// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 11.0 linux32 Build 157 04/28/2011
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gT8V+RHSdzoa1vERBsZ06ML0/vKl/hnpdeNiBkcc7Co4P5WEnUExGxLxHMC99LPV
iHh+w7NHvInE5nqZB7YHTyylbtBcs7aVLgRaV+QfyqV4ggDbkf44asaoxp1sYuQa
Ey54QUWpjJf6ttGGgPO/EUGx+Y5ica7OiCNStGiPZnI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 219648)
1ljpjUGoO8nVncJlPYinAoFmnHofUuajfzn0ktcbu7KSKobu/WOhNuD9ILf0LW1Z
KwW/W4G1NY4xjjscF+ie38zU1yYS4hC+hcZRl3PROf9Gn3A1Xciydc7thuz7SdAk
CFBMp8B+wwnAsf5geHVVfevZMCOEGUrjHmnsK5r3fMl63JKQLOEVl++La4M78mkd
Bm4Y4+HDFfQ9c2pay5MuqcZO1sehlxf4sq29/VLeT8AJJrABt/eA038shxYqLOIG
JXdy6iECPWlOt7KVsxZtBiBuSlR5yJQSkbCr34tMmEcyiWQ9xJU/IywaSb3vy56u
O8G689dGGc4Ffcohu6VcXTp5fo/cx179O2vZzfWrDSUvlBriVOHNxL4zU1cuTFxX
sln4jw+o46t0ApnIqQ1vr/6BimrROolarEg8qh09xIRpVks13VPcEGteyzcwb2ke
Q+BQrmFlpzpTNmE1K82V87hupRZyxX2tO18QJIYXsCKGVCEyrbxGNihzftdot2na
3fcwH/CYsrrhjczBvlekkO4ppG7VCOJx1yHYYIAXPpJTiVQrihHc/qYgx/9I3c4b
/IAADX4aD0uS0yZD/9ZnoPHtkbOzsVfcl9avZHCRHvn4qo+kahXAU/j047nmM2q4
4iTnbvGSIJ7i36/YErQnDd2Sl5gf+QE/VHLCvoPtlcCBT6VC25L1nu0eoRj3hAQj
Lw0qPnQfm5ZefB+hRNBV3kC0bLIpQ4HbP3ZgiWC8oqolfplpK07r9QCYetPZvatQ
MRQd5L2O0gmEUcpgnYdor2H4LOURBWO6Cg6D9EswwSsRfBmTGbx7VSWmYWovekff
HPVFwBKf4DmWLqLlHX/qk9RaUpE1oTvzE5ZyJaXkhFGlKH5KRiyunjJ4pzbtu43V
2n3bU8OHbQaatqEuLw3BaDxDQMwzB1xE+YzF6a9OmZvmP4vERB/87+2yGs7tMahf
h1tUi9aCP0m7E24Cm/GAC04TdJzKIzSNQmBI/bjXqupTko6oTHDr7LLTeFNPlfNl
KrUx7HG/kEV/f98RhjVE/m1jj2f34fJWUEPghSPnku/PWz9Gfm21nhqlg8e3PWDD
YiuYMfK2O5j6WzBMcZ0/7jdSUT2I2htAPv1YVFgqXWCYU3YG+a7LlwdiQ49Ft8Wi
2sofGLk1N1Qb+HPBQ/fRpzxiH15jHHW605Z1FI8ETO5EY/iWHPDuuw9+SzY6eG1J
bxU/hKg+MMyKP0vdYQeyMztHoTdg0OOxy1uaVbariAZCG3dxua4+VwSdHjMYdLNM
7tn1RmZCsR76weQqdbaHOi1sx8A6GVQytG216j25CgBwLrrRSFCdZDKUudE/sdtC
MFFLBz5XOnsSEPV8GS/WjRozqjSPP5Qck8md5bhS8VDRV5waMyAxsOJ8t5YcMoxs
LD42LDru4mGRlKQ1TqY4h/OlQGWJRiOLe7ueHmOS6m8saSSfwql5yIsfje8dTu0+
AjxP1kSCmblABdO3+l0ESp35mCLv329829w0uO43nzp6EOqnIoi8m411HRfZ+C9M
DltNCQZQpGOMSukeF1ZDv/ZMDy7m6vq4luPqMx5InRz44VoIw0guksv+RDz/dAZc
JgzPDJ7wWswfyol06bRCdh66vEwcpkY2BU3qqulRYI1n8v4HPmQh2ZqI6eOye9Bh
n4QZWg22usj+iVYbfpcq/sYSYBr4joHxQzGKSTB0m19gDCQzqbtBxcE0m1oiOQRM
WdMchm+tsdfMnRi3tGHSkpTC5UmspulSb3bLk09Js+0uBMxkLaUi5RpIJ3aFZZNI
3xIQaIyeZmtScTiNKPxDGFLFHHDKXY+oL8IfpB5g97qEu39t2xQT0l4QdCMN8y+r
BTc6+W8xwPQ97+fe2eJZKF6vm4m/K+tzmnYQ1HlmZ3K2sgv1mpPymmdL3KIOr+Ku
5eojNDhrW6vQDYHK7L6lNm/8QNdm8bMZ9026m1yHnOZsfEZxfUCU1c/EePamB/US
+sNMNZFkN5YXd4q27AmdC/bnh0/QcL7Kv43O8jVjPsRplj90ymTI4F3B9jcRgNP1
A3+TXc6geHMelgfq6ZaPf0AfxIN7CBPghO7LMUaDzjbg+YxXvLOUgJrS1f0+lsOu
MicUkV2nJO8TqRwMXXdNa2aWXNZRd3cgPWAoEl2eON2HlDkeS23eN2sjAJnsJktC
xq+J/yEWuI+0O6A/K9lJPwE52KRCDevskbTgpbofIEYsHYKpaAU9o+oy4AZR4wgV
OSvuPMOkT68M8kFxHPnOANvQqm7s/8Qn6f0iTrqoR7jcqAIblUXGpZfN1uBjlIKz
sYG3iQijO4t7reUifWwB9tRn9bPkqafTji2xYiGPTKd/hRR6EjBLjXDOFBcGyj9C
kKfKv6TjrmdccYgg1loqOT4smIacdOd5n+IdwK6ynfK0M9pDYcEuIDUTANIAcany
Jyr4NyCtfmLtoglZTe2Brjctg7l8xsuF+D52XQKJNScd85z/obvHVstiUBvvXBmj
DFv80NF5Oo8fr7Sc+3ci9Oh7COKdeHQkbInOhwVYCbyL1nM2RtoMocTDT4SiikXA
HmgMtM0hSJWXD2XXffu7Dc5esIrDE4zJ26kaAdqhVcEqZPN9kZ0Dz3X0bmc1aYio
RkMgMAf+8inh+K6zYvUNCoE/oyn4UTxiKi2FemTMie0waVQbeWl0Rcf0WIq77ypE
Ud+3q+b13vYCyuwbM73AYrSx/75r7Q5gUlTEiF3Eg0JXPjUcNj9yKnNUldBdnRxl
mAJkzsdYEB8JwdvKg5RZKFJT9DtQT2NMc0T6D/durnl5f1XMtoZuP+ouZyvMhQbK
3OObYl4OPsZhd9W0CxCObinUd2VflWOVus7NR6wLhsR5NycaLk/xrpj0pUg+YciA
OvHew360YoaqrOH5oq0c/wDTdOJYZTesYxIoZFCIqy9tPzGvxBq/W2tl0f91JhXh
kAQ8SwruxydmFilYoB2swpYq0fyM2GaOFkwOpTa7ELeKwIUH05Jx9cCzEUdOLha3
NcRKpxyd3X4eL7ZiJkpH7rYlrTGvNIY99A02I8AX/Afb/ZRJgDQ5j0cPL8alMuRp
HZeeHBpQJkVxZbMSrmztyof7rxX3qCqyKRHDdgQCFr0e4GRl+2rTJbQDarLGF/ba
ovVh8PxKeAKlR8dfNo/ovzVefeCuYdZQXCbu3PtbU4ztanEWzwkvZtaIzZ2AOIz1
Cij/KpFr7ZmsZc6FAXGB4SCAJsGMnZ+crXeXXsGnrJDX4wDplyCuASRtEnd4O3UB
jP3Kc31U6tzF1QigJl3vDRCLHSNEymfGjE6OWRj2XWRTuWveoaWAPP3KSbglAtgv
1HlKtrH7+spUmaA1uQTGiRKMsAj3xpcOpSh3OiEp8Sld3MDl4Ar1Mqv5LaI8zrFE
JLmQUhIu9/zvsi9aTZN5fn4gMBbr67HuTNOLeAtfLdAnmiyHVmuyrh6lucZggNsu
bZ4oavG0mGkrT0KnKqZ+RapBPqZaFz6zOQOM8gvz2f5XgmOyHeBIMzb11MLw6xa+
T9D+wepz5+L7oqUb0s3edPXyOUK7VITfK2PJtmls4p8xFKexQEPg2sUGX2V02+42
wbcd8ynQqCZTxOJigQ4+nOJRoTPifG89RXV/HfSCtZvcv1/h+P6e+h73JWYwSQWN
/EqEjH3yqOT0KJB5bzmKyM7DJ0b7eOyLphyxtfY5XbX8SVVC/oks3B3h8FZIiOOO
B9ECwW1irCy/lpsksQQCXpgH3IrW/W8GdfIBPvvbTI2THYFuIO/RRTxc/E3Spa9o
PKYkzWu748WyRbPbvSeml6Dhuhi7Mdgy1b1f8fNIn1GIc1fpmHDJBPj5uV6eO3tS
jVsWE8ZPnDvPegw5gmflaEmrqMFMKTK49Tq+ro3su/EeQ2/qmZgH/HFGTfB+EzqU
YeYQP7Yk564iUh3x/Z+BZFxXZaM9a7kruAb/aGHxRcV09BEpnipLrAOdVMz3G2QU
HV88vKmAqJgmHD9HZru7tQ/UK4O8b4ofgRPP98D44eAWY6r6xTqsetwTR4HQm09M
g29D9zkfGUrLkM/sSxfPijHEMqcArWXN4LoR0AFk/wmf5EhGcpOKNuMbD1bj4DGG
CzNK1AdWgKIR146memVkRhkOtPYBOXCWnRLNOP8i6j2c1TX0Y1MQfPIjjkjGWe+l
kwAd3aQ0cFoJ7rmWD4bgeLMOEjm2g+mRGfyS9H6nKwyTfFqDkVXk+VFKUufB672z
CSbqAGj57ylOyX0sBAsSsG3xGH+dnc5O4KJBDQyMouPy81dLvL0/2A8/t81X1Acg
TbOeeyHpU0DLZmsM6U0+hfYFX4w51Agmufr1cm2Msw3hGWsL3srvntfutLckaMjm
bWl/Ou7fC6EQuxetRWH5JJcJrwY8M0hyEm0h7qXRj1V8GLcRzFJqaIgSrzZ1DZH0
gimz/mhrpbvJIjg0dRGFJ9+AmRu3dXRPFBLgXePrSmbJzb5kGE+y0sKHUpAxTn50
GzJCVqAP9RUJYSFgKH1QQFplCinP3OtAp4TBK4MAcN0XWWZ34vmiFrEZjN3Q288P
MH3YWTZNbFdjWYUf+rxzfYSO7RvSR+DKukJvSN9DMXj5cfviuU/0JReSeCYJIxoU
gEZp8MwCkJs37OZ7niThQ3vBZWQ26qdYgexAkJVpKp9p6DiMxd+zFVXayuNij4ch
cMrL1dPRqutASnXgc/NcUtkZMFTvcqpQJ4xFFlhfM55iaYv4EcHCUlDxfYOiVtEZ
SfT5HwJzNql9peFQ0t6hcxjpVSvfQqxg/E+4McWAcgQSyfh4gHIy0HjheqQZw6Qh
d18pblD+3MQMpTqJT6GUAhcGDDjMwFrB4OPuKplSSUymU2jurfroOjLi3sp615M1
EbzJNmI7RgKHkdezPgRDXF/YrehB2KTmMe1lYAezIGlyliOhxa+8ceZd8xmIAxfs
MtJ1JxfQ5OrMzV1MN0js0xjMQeR6NzcALm4zCtf4CRke/NXZ4gsW/W1DgZ/ZoIPL
Na8hfRuclKQH/0P5GrEVWEi///6Xoc3qo2/fm/AhRoN6f/VUZPOM7NuJ+FFzHZSo
i5hlWiCSnKD5hsA2oW5Lbh9Mkv9HHIdHotG25zDj9V3oQcTaa+T+pf0tODUXL4Df
ANEMTNb4lXVEihWTLP7xtcf3bjyGQAFhKBhBpV7wRWuNzMXsJoHyS5xY8aM/Giyc
8bp9TYvSMd9rralIZM7SyZBegNVqXAW8CAZn4uoxQtJ/VTT9V9EzE4DY2+ybuVaB
4F6DJOZpLuGMEgireKATpucncQ9dkGByc/hXmJqAL8etdAUCzLAxUssisN4N+f0O
/NrFHOricchI8gOmLeF1+wLy1UFUv9V2vI5w1DZcTMJetweeQJUPFRhUXyUT/zx5
DA81BAiGKmFvdzYnv1MR44mvjgc3UZLubceKT3ForpreXWdrHIrDNGVHguQcKHqv
efTmD2d1qlCyU/++mp7zwx01ErJJUuytLLWKc8WJQaWZvPIiMuycU8gigctN0Sbi
4SlOeo0CmaggF5cbhpKgWmjvvOLBcLl1kVKG0ZH8V0cMVEwz5Bycd9wcLvDBPVvM
2EnJYXCkgP++LP0MjBVNncLRhFHj6rH4G6amZwGaQL5DhGzQ5u+nh9Tn/tmZ18vb
GEjXyeujbQsT+xVdeUzHSX6JyweQYcJTQPyczkbMSImyXMpUPeavwv9YOHNz3Teq
QZWwDb/aFQsCKvGYf2Aq1F3h3IY5U5LxP0LRgHQyXKljAtZMuB3PGfcbzKSndWfJ
QJkUuojs6SARD0WaW4z+DLINT++WK9k9oDJdM7dQ0hFQI/atRfEN/LfvA20e4k40
yg3OsNbK9q2cWhkM5vIAKzPU4RXPtWC6JlAUZHWRmGtl1TLq9HVB1IVygTaWgor3
uM9+xfvZhIcehc4QSQfoqZyZESInx/viMGz6NgJbYvypp2jL5q03L8cSyQp4G55D
USNQGmvWsXl1bigA0Qn7pT7lUFVE+14ZFxYxGEBc+b5/6ongBFQ0Xyx5IkLrIfWR
mgEBYmnOA9MtiqJ7Sh6C/8430uulGGvGEcZAxzR5OfHua6DvVrllblX+68kfhIJP
A9CIKYj9tWo4LDnEUuxxC5SaPfN0YpFCWSMMpFImE0WMNNGBzeEmCOzFu653uFJ5
o1YdXY4sPMXJGT4I8Cq0ejnU3V5QNmlwQYrGDSxCZfvBHCDhKqXdd7Nx5BnAMBkw
xWQtVGahapIeLZoGRLBpXpp9APxG8hpg8bd2/pEDBahQdzivsknnCudfitydtXg6
iiUQbYHjyPXPgAeglbAGhR0+OEvWlvTG6eBxjqFwYNTL98w8sEWW36j/JF7YfONf
UGjMBBYtljMU9bljwOwr4j70JDQIf0awMhAQS/orLQ+FNJuOmalAGO6Q4RKjc162
K5TAaTYqkq5FPYtgBwYI3HSa77DlTHr4dPq1FWqkL4APXa9XA4TTti7kbtySxxrp
Y68qizz42nz2hwpgtsszaxMIoRRqOdJ5c0VB0DTuV5zcyVMuPI9EdPgGf4/7EgGj
9VK2mk2l6bU9fC+PYqPi3MCRBSw84zzvhRO2xdllt+KfagQQuMNNZc3haq1OB7fN
D03DPGEXua2hMu6aV0MKp4p5zBMSqPpsQh60WZ7WGnO2ghNTRnaf+Rt1b53Qx4B+
Q6OSjNpdYWDsAyq5WnaL7l3kkGSoA8FRe6RF6KjTbDa9HhMKowlsyFO2xnnd5Mqm
7wtmqYXoXW8arVE597LGk+83bNsC2+AGodKxXEIPHLwDWdTHCGfo4tXBCPKYgwXh
akbaFAoHWgYB65bwtT8dlLvilvRhzQmtoESiO1LcHY1bkINDD0ER1wDgL9Qs3vUV
DPLRIro2mYYaq9NYHMeJn6R63trHYI/IdDJVLD2FLzfIcVCytb5U3HKO/xyScaxx
vJzKvGrev8E6zaqW1WqnMC8UDu9rAU6LGuESC1hf6j5PpfP/DGIl5/KRP1MBjpxY
O4S2X9HabA07EPV9UIjFLeo61AsuxaIT+W1pYpr0m/SbVgCXbQnv2DRtPf/PbrCZ
qZoFlBCZCO6Ho4+00khH5I8CcbSGMR3hOcaagLiQS4HdrVPTcLlWzoVeabjEH3HF
HLqa4hmI+gGCoMzFUsdpD9f6aBqHRJN/ilR11CP3xqZBSvPfDFamBuupDoW/NFz1
mWeAkAWtvcZtBO4FTDy0A1c4K/WR3F8HwwuYoWpGkxPAfEjjJ4o3/y62gEH6zJKw
ePsf5vzUrvXZ/tF1Aw3ifu8g4j6faSI5PCldUdlJxN/5ksAChvbtGj13UAvS5uEx
OaVcNwiZxByWHz7IVdacJKNalWU0RNk5lCRzuLrw/RUxNn7Q1RmgLjmwgBAvEUfE
hCpE/rsuYiJ6h+Xcnk66rPWBrp/uP8TKljnRkoDIgKpJK8IbX6R8v1OXBcSnCDDA
p7j5cEBTbZ5u2qQqNCEljJ0ELFTitNkU1VKByHrSHj6/UI203PzGSWYtRerFA7PS
alkZfRccj1sbgwm3NsVJByL1KBPUnFswNbNziNx7/AK3oLhW47FwMzvtncrOnjJc
EhIkjqj57B9d1xM7JHpg079Ir2Ye8xLNIzHh476gQUGHzOUcVX2A/jQxrPG31GtC
ldUCB9+MIOvXwaQKnUwS7t2SnD3rKjlgkOQX6qrLDYzTiEEVb9pC1ahER+OnImQn
cKR/Nfl8r1xTBN5FMoKVCxsMOdjZp4TEDtTFCCoQCsP9y5uji2f8KVNnKwK2ioU1
Mt96NWbNlHrlfZwkizma/6e7noV60puZjuR7iNbfYqPZMtVYpQVca20q9Bkep1Eh
4jSWh6OSrbU2XOPIjwheparJGl9Z7Ytqn7/cGg8QI06lRQTUeAEoF4crLeQBwhZq
ysiACSfMGzoGuSVgDkB+2oZaUy00S01DYdJlVvf4pSYNJyC9rtTpRLJx2t5ltSLC
3KSAybwjaIAo3PNIF+pgwVslm98gDTiKCuS8avCI71CjeXI+o9TzCsGm6nDjQjHv
eBNdJ/UVap01pchro4tCTgj64Dl/wpq6CDxQPVkmGYbOvpOTHka8JZY/rQ9Eq2oj
gpz5DP7X4Ag78E8cBAX6T3G8s32oJBsnny3bO7X+8M4PtEauTZD4gGTSYi1ViHhx
iAxA8s0Vk930ucesPM5JLzC5KSVTk4BbWbf3PWTQoQa1zHi7m8wsRuoTTHuJy4An
FgpMJqv2nPWFhIBx1YUmknbnG5z/5wTR1hCMNNXjSRJGpj8/W85Jjz6aRjJMe40R
AR09FAy6bosQJBY7po2+hx6lTMSc2E2+X+Apy5NAaOpWSB1iKdNGZEoX+dQaX0Uq
d+mlL0DQoi2mjOQFLIr8uuG8JSJ36jw9uai9KXsOybAtX8NPiXFGAzICIA6d9fOJ
Iedd13U5hGo6jcREHSBoNJ9RujNyJJ2KKC2MCvT4bKI2V9TQ06l4Pr+0EE+dj/cz
koRCx0hs3xMFpOd1SKA5VkwZJj4x/QIrnZhnUAFNhZt1YZtNCltQoDapYq9b7H3+
pPx7rXPA/eN2axQvNTx5rJ5/LyNSJHLiO4I43dR7Z8YDH+Dv8sRi3RQD8C5BxmtV
uOyKvNsJ8xHzKLOFHghtBHklYWJ7MxzTxIDJ4AYMwNBe5kkGlSY/xClaZOsivbUk
r6hUHhx/vzWp8TmJgZcl/aDieXGY4plOKrYKgSW/UcmrIb9nAFjYsPGH/jmqigpF
umi3sqHrqcnsV63MSTHT0ryxaXDrssi/qS2g+DDFRCz4XkbTif7YdkaKowqGZ1mN
EtCIAI6KpCk3AqH17HuOH3o3H7o0MKxhUgHtmITmnBJ2mDiXkDHkWtHRjze6b6z1
Tc0jExv8uSAUoIjGQRxfaVM33E92TzYDX5iEv0NEs0Mj/E8PZSbxQqyACxdrsM7S
inSercnPImxYxMFzLnQESHb8NZDwwUBal61mRD62pHVJcngBlADci35+//SAmIiv
+tcN7WZNFbuwr2+NpKQ/JOR+6FIGIXwH35WKMS9OvqaZHxBiGIEVj1Bi5UC0ahXq
DvlXBdwvBEwiDMZpS7B/RPq0KPBZCWOOFg62gzQI6MAGr+4VQtgNHf74m2+wXl2L
/poBE+Y7qol5UrmrnYHUIFNhoN7J43nbWMcx3ShpUsA69btFYDbrnLMlf6WGPz2k
Q3jamtbJ4gwck2eEokwT+oifLua3Rv+juipWysby3oupKro9YcMVLqsn8nfgiIaF
GwTvivPzhe1AooVh2sIu5sdHHPtKtSNc+THiie41SlLFxGBBOZp7UpKf1abbvSQh
NHuMZCVYDG/uIBMw0n5mBMGeLfsyfRdtuDgjI+z4nCIHC1CFaBfW3Ie2l09MvrTW
vY6B85oHxyU46K6almbtu3mIxe7rVu/MXRW7Xum9fBYHSIQoB1pdGX+IdsL7Uv4v
rvdHpOFr5Mb4qGBn1EEaq/EJwo1UahBcD4Mz2jqGO7ySZcs5S6nVqR4JXKOSBPzo
P5OlQisPHTEIKp3gxlMJO9v6rxFzUGXcO/UW/tIM899HydSPAj/25zGfHVsQAmNW
LJmq+yl+tcEakl32QQ+eXRz+lJFq2ZubkVgnQijvuHUZTBmIgbfzSJ23L2RmHwWv
22UhiU8YsVKwRh2dHJwAEMpt9DmCaUmBEA8Rtdr7VPWB5bAuufVEUYMKSEjgmk/d
/EfWXic6ZtgkRvievny/myBPQxYSp4OdQipGmXqcV1HOsAC/iU5tutB0EhbrJ/Fe
sF6Nep9Tk3RUPV9AVnk2OZJxSMN5dO+Z1MGDJHljzJT37j1zpMz7Wo5lDlz6+aL/
3Tod74fUxHnZdF45vawBjOOyng0aA/XgM5G2yULnlRlFlay41RjxXULcvxwWfhHy
Tt+NRm/7TKnNLcRtiWScuaTVcxayQsM7AY16Z81/S3kKiMxVR+lmAhOuSreJ50jA
uPQzIItlk3t8yEclZDIe5VkjLGxgxC2rwdltXjzVZvV27KSrbppBTU69JSIFU98O
AeEa1eCXZTvqq5gUkBNidQ57YgiTnBbVrSPTVlGsvjv/gDmQgzZB5XwuyVPzNHt2
0acozo9NHwly3wn69xR3JB/1R33BmhZ/bH60ztF5/Vxa2B+lL4xZSs/aEbnovyaf
K8Crve40DBi5Mo32ZXq8PTWCMnPVyYp2n8rkvP+zPyVADVpWJ+Xuq39t9m1HrbdK
a6FswzZrkjauoklCNV8MQTeJOTV9HOrbO8zz5hWmL4VmC98tsNeIu7KHPAp3I/uC
e7o16OV9fHpxMBKEwE+8fUhEaZPF5r58DdXblo2+dwDKThtGMQcw0OhaFjbusdog
qLdCkkrNeU3WxvAH7xp4LYqA03izvMlO5Ky058if6lAOhRJ6NcCmxlJjLsc0jjyO
oBuzrnraZ+r6/xdeqDRWMKS7gVp/JCuhnV8kfZBNTvaptgtkBbKWop7t5odlS/D0
9Lr4VOiAPXPE3Mvv5mf9gVurS4QFmVw1CFnnccYHdhpnmUabpAMjXRsYwJQ99+sB
3h0534Bh0sxZPSB8ZdmeBVYn6Vft3oluNCLBwX0Oo4UvO6s5qmtKkVsaKfOmMBTG
MhosvkhNLdDhSfWwNvbWP8TUnaifNaf41coisWvsLLC63Qppmuvw2KNrgzgLoSMT
wOP8Do7O9h2MVCWCDGC8mjrvACvKgtcYEplYoiXE0swXM8mUF6tlj7JGqeNpEy3g
0mB/Av2CvpgIvKlAZijCQz5k/zui5mq2sM3OjDJJKqa4ZVUMhN0ijhXLW8XqSFQw
9FwAQ8EyvQYhoUZ2EOQO7P1rAnvMhWqW51AhKNt/GThKNnqfG6AqTDQAx52cllu1
D0i+QqQbDdaHA9TYCYAwrPT1ax6FdIOHGqCQK2Mhs8GstBDJt1L0m0rIUI2AY5Cb
U/Coo7dwLNJ0bcZ+OatDPXSIDtUAXLLmBRhfcaXLzVEJmnrfUtAlUwaK1+9aYSLo
iqen3gDX3TAb69xQdwYsIAWbSrwjDkWC7ygWqcl9A026XL9J+xu9+FZgiGY5mm4i
XmbvxXVbG+Iy8la/XyBRLFhIY4djnROfiBk/5UkiTOtI38PEt4hYcd02q+uhMk4n
3uGR6ZLikINyAjY6PXYlg1ja6PqEQP8kZEQM8Ip60qT2+kSmIwF7CGkP6Sc+k+y2
okuRxFeE+qf/P/EvbkR5SQkkcAUQybWQKoGcVu0kQyBeXAswtyMtC/my5r2IWtxg
wzBMzQrD4Bircq29W2o7oY/NfivZJADHkR/PTJe7pmYfM7a/TXeiwj7vUcDudz7q
1k9cLiGiiEQymRUu8QbkGDwZez84Y1YHrOFdiCyB+wY8vydUOgLq3VcUqGccjdWh
ZqSA/eMcC6JL88Lz4cZ7CKBv8tWita+MRqPXUNGa7VPpz53IeDSrPRhmIuTzbN5n
575Z71bUm4hh2ci+n7uOgLIN5BrjWVWtqGYWJVyCt1jdv2/DvHtdTRHsHAmUD5FT
9SzzAiB7vhg7hSwCWkdgl5fGQvy7G0ryTAUeojm3GU0qyh23S2kxL9wbHTmsEOZy
NyT+K5i9Qru6WhPpgf/ztDJsaJTTO+4DxAHjTQPhYF8F13ISdyIJG/0iGrGRN6bx
/pNsoiPnG0k8Vd8IrU/DtQVTtVgAQiLQaW6iP2GN9CTPLOatfokjqmiFW1ELfMy/
sW911lsWl4E6OVSiFM6MewvGG7wd0+O8H+f8dmaFZ5IAYh5lztBmAEGj0nbvTueM
D8xn/mVCGe7vHo2Y1UnXjpE/ba/C+MnXq9rwtXveehxS5iBuo6iZhx5ui//uv3rf
YK1YksEZ9IgB+rFtJV323phjuK2wsmzrge8sEzFe293Eo6WcCqoeGntELQXMJ0n/
o4ie4xmXnIQKA3r+w87qnEhktSRuvi5od6trQU2M7G4ul/FbeFnN5kCJTxlTOWTB
kY1zDjdqKsYC0Wzaf2tp+l5AXrOEPbl2T22CvJlljchYs82onVWBnxBYHKCvc1i6
pAiDl7gjR7q7sIYSjxQ5BUe7IizUAphgkS+8g+R4mLQCz7sqZK1O21LaX0PkudLf
LjwYccPbIUmJCMDAPhW865n0P0TfNY65Hl+7eUt2tKXM15cWTI4Z+jO9osbKdKRP
DJalRoR6wJP7dQke1ASD5QAPIJpbTpDQWjM5HEyfmQS7MWOboNA8Pl/vccjlHTPQ
I8FbdY1f9u2BZN4vxmNApUrDC8FGd8dgYzEehTwiXup2pABe7DUTtjD7yuUmRwMZ
yjw8O1oCGIsKcGaI8OQ/6z2zcsJF1CVtfJjPtyodktkyshh7XswP+F+oAsZGkJrh
3AdmbAkUN9v5NgdoKYhlSazT+IjW5gef/5smOgMtPyHeTm0Uuofpc7aF2FIAlqAb
tsbXFnIIVOzDvCBSvRoJZHKIp9Zyjxf+SrKDFoUqtF1fSPcANWZ5nHys7Z+cDYPD
LIvIz3cwAtWfIwOf2NChJQbmVHqqmry+N8jmXwUXzD5J88VmInhnlWeO4jG7y23S
bUJodXfKZgMHuqL5oPzF0artOtZOlb8Lg5puS1DQu22lJTqaMglXS4PihO48t5CV
BJbUJxgH8M8F4Y7Oli6A+Y2q8gJbPl3p4ki6C1u26HJ10fjCzd68QuClDlNZgMWh
DnmWKLjf3DzDCMvwvMPaYaw1bQj0dGUzWDMffiHqVp3LwZ3llUYV8SmmG9zg/gHq
eC1lLQTG44HKKPYF8BoU6RA0YEXJMZdGLpBi4SGGzckwRfxUhYsfhlkMuS5LK/rE
rhSWnwGW10y9OnuWOIKVDCRZYFlwrNpLSmIGZidvZnpKje1GFjP9Uni4y/8wqtN5
qw2tNDgvZA1hPlzMFNODtIL9rsI6zsw2G1DIp8ExXlIwTz7kImX1yHFhuJd48D1S
TqBxWOVaNWvXjLzLRTMHQxUo+DgpjVuDt4zn/nyN/DRpEyu5jfDG0+ol74mrVb1+
mc7WZF/KaadQZIpmSMBif+/ZXcmNAMBhUfnUaYNJMzPQsgiJBAnZs+vdPPOT7HNM
/u6ihXprKo+gmTqb3Yn0evl41uy1DtowX6kfORJwc5qpL+Y1o/ZaK9uj4t0hRRnQ
LgpzFDgldaRM+IZj/QVPCVYPtMQ8pwHDywc+gtLaNenTjK/VgDmLl1Lq2WcOkBW2
reeUToU266dPl0THH7MQXEV+wrYMRYUr1E8P+ecFy/60FNv27EiYTRqI5quIIevK
qtm/WIzB/oxdt2dmvIVpodeVHVigMvAXPZTI0EloYMWn7D59ayMYT86SGJQFlZk6
SPKT/aj2rmH18w5tGRFhUndROOh9UUA7wR1VLUPLIW3gGjmJU6k3oNgOyBF7WRY3
JogY/RKf9jLKB9hzF7j36VnaVWTUyCq1u5BR/T4dgfFsxxWSmTZjBefR6cEuwQrK
c01qPedbompIQ6DIQxUdJmn9clFGmSw1kh02avgkMAnwQMa0WvxXj5lOnvLKGiRD
VerA6h7i6nLN2CyO47NApusPnRhnyD25GckVQ/VMaTHnXdKXp1FI5mpf9GF7rJg1
EPyCAzU0KawM5FbPAcoUYs0iUpPAFbwY2+ZHuk9IYjFLi/65VH1puc0MakR1pret
CslpcjcXdv/FdR0YD1pMzBIIJ2+Kqxr7vP3QFdqWIDYVb+AgKo5vCC7+mzdyPW0y
WGfx0TbIeDAT20kHVwaEWs3utdob2pfTya9uycKoKu5Kj9oRfobIJCzkeTVmANbo
gjZZaCe3VIaHU1SPZ2MRB81pmLQGl3fkqQTPdInzMi/bLbivrIZNfFQ3rO+/0e6w
6k2f/tRv0IaqpUm89hf8sXF/7RW3r5Ctff+ZYe1sDb+Yz/iig/KlX4XyUumFSC9D
tYjwpF2AkS4a6hHZH5heVNBHhRxpd9oPIbiGAzkNSHWARk3S4RqdkZGnYu41rjot
dPto3YK7Xbpys6ozvmhskdSTW5vUUN3L70Br4m6/a3GlIK5yKCycYNL3FmE5+hvS
7w9bByqZqMfuASxDqfHEHjXLZXTaYki9stCfKQMRFqMypibmp0ybaDCZ1alcuVFE
zJj+GKUqW0gtcyw1TSe1gyKT5U5eneDVWOAs2JsBgz68Ype7KEl7TijHdsOd8oUY
k5hdAGxdk35HCz5l9C8rDoN2LFVl30S0cq7eDvrAoA/8NObWaYA6cwk8ZdmQ3ivE
0XBxHpb0s/icYXv+4sKHa24W4BqeEAb3NP9wD+V2lRqBnsQAFjP+68iNLbWHUkIh
W9ssJ2AzOs1yQn13EzrHEiMm+3+DwEwSTDNE3ijHIeZ9QFnrf6u9A7Zw+/y34ZgZ
rsrQj4pK1EPnwdmQsWibdRIwcwL9YKGgfsFrGrG3nDObcAvpBiLS94WZLQyWILLV
FEWoap+585X9FUkQbj+uPp1GS5O0McKQ0kAhBl7o5hDQWoLDwaXbYp25TZl0HHB9
q5CmwYAHx+/dlhYayv84BfOJ79NmLRd5mibHfVIjOGIQCVPD0Wr3XPqFZHLHPoiN
l0AS75n1zSpC7BYaGpIwLkHODZxru84goXoRidVsywV1KqSyLdlV1np2tEWE31F2
Ajyi9RAovpiaEgOeH+QhycCdBgWvZO/ehlxqOPZ9uyyIxKotxJtMggdiTooJtp9n
7M0Pcxfkd0QJEO8XlM8H/J+obeVrx9fFvOQy2eE04UXIBIIiey4XLxwqKyynXEo/
Fu+MIVzS9G+/EpHOO1aSjTuLt5d4MPgiacVu26Me35hrji/91zHLonRynWfvafLn
pqfFCc0m/34n0toS15cHHFnEb+v3Oyk6JZjlwyi+2KP/s6AhNHaEovrGVpAsRmnk
kZXVUIOqV6vYGP92bQ2pSvfhUtVqFbWgX2J9WyfGxeMIT5DbhlFeOqhQznAAXvj5
p9J1+MruANwX1L8nDH4FRi7xki6pb47eLfC+864c2RKz87XHfdzJTAS/C8nanpud
vNl70CwKcojj0IymizHWGOv6Zac1f3d4Sbgid0XTfLOP1HLwnRo89XWIBleRYdp+
4uZs9Z7Rn7hU7Uh7nu0jTpzF8PhRlidPl2Atert0r/fxuMUBcUyw/0aoj2Dzq3dG
f0zoYlYhaBhpaw9vN0mq1aaN+ckCZeG+8ZEosWGc7GXLnQ6H3exSLp9iJUQCr7M1
ea4XOBNs1IwJ8rEWHPa+uZcJV9KsfbpzIH1IyObZrWcGsapigxZ8tRlLA9mZzSdf
WfCf5UgiKuZWLhfyKVZkitDnl+ZxJRi3bW8n0QURYbRyY2A5Cw4pGjh0xX5yPLbe
U0krPU/QE919xHfqdCu/toQP1NeVORTaO07S5VFvpWZvOIChhTPq/sJrlzwXPUGD
osWqI5OvaiSAvkQ/XgzeNwhe78t8w0IVc0sfEP/F3h1GMt/BSAAgoYeNYusxmCQk
3HQ0bRdEBJ2Ea2qIW6ZyixKmjQG89Hva4vUT+fnGES9P2rmcd+djtQX46kj6aPfs
HUWSi5N1HSG41Sqx3XiAPyEaecvGEytmvF8qh/hmXOXJzi8tXXNVsFJf8EXN/MRk
71/7KS22nNWb2qbqLv+T26LbSYoWVhUViyzorNJ6wCofo1QEIYzm7yXI64DTfFPg
mrAMJv1+xOwdjyxe6GonWZI+OkGXz12jtfo92KGQUjlCoPKyKnG3t2XC6+j9Cvgk
4hlj/NH4yeWrbojoiZ1HhuYrXx2xuGmOv90uEDxRLNe8mJrzKnnTNjmh2F3Ra6UG
zvyJc9SfLjsKzjxfpWM7dLrMB2UPJa19APqgN/Mp6x2LKyH9yDsYs00p8gSwjKeB
aUF9oUSYO1L2cX3jJLzIPT2zYPn0DyTyRuO4Rx4a0NLo7lCfGh1GH0vO5AzSi6I+
JE+FOIoFMuOSBUusRHx78hJNnZLXMBEWnJxc8l4VPULV0Wm/0wwU3Tey14jKfmBR
QnVlE3lIRxkPqaclWdDX4C2gjpEDGw8VORIaE07tvUzshME6CK3Sh4YW9T5yY45F
avfGoOxiHEcMStBMqMl2mdYsyhQR0CG/38tgFPmrfDlOroN8Bhyc2xr6dpQM01AI
yJligFYgRxHmMVc/EeBE3Pu+Fm2YcmyHBvYNUxeaEaB7Mh7/3/ciUuZr/iW3ASVD
Td/hFnxXQxT1uNkMovqjsHljoxhsG4Jk4QvK2GJWT2C/5XcrDCWU3bHTQOmX/24A
ClaAWRvcxNlGxVHKcZvOzPigPNAZHMPEbpen5zijSygwCO0wgLBbphuKjd3QGQs8
KcBDHI78ZPYE+IOhrbsbmTMF5no/tvSg30PjwjsL+CfRtZ0BnhmoPOaMPfS6x/ZB
EDIGpUsCHde6rvZpkc2orwOcjBKNAqGv1kxuknZdDLZJiruOfrfKA+JZtAz8IaVo
Vn0G1NoLK26VIC4z/2b7vIVxU+tnffoLfGSHgsucoy2JoecEKdJhKLcs77HIn69N
6cF3mKw0DQZ44v/U98PoiUYEIDH4mel5LxzIz0Zf+ixmPkOPa4eNr+MSBXFSMoK+
L/q3wfOxkMky/vvwk+i+CxTrsGfzb61aEA9DBQqMG1pDPY6xw+7DK5YBJQDySDbQ
jAH7Xk3r1HT+YRezk6e+Zf+nCF3dM6Y1LNohx78qZM+65sJVApN+ne+/72YlyLM3
Cftv99NpDM2i5EnRk+2qUOcIp0uWcq5obRQgtoJNEhisAGOUHIWUQqiEIxFB28f7
3ZcZXb3mvP54RxgSrPrBQPXzVXf2wgv2KEx3ORrUDun5S6TlJDFvqlUb6uCl2tIm
lPr1EJ27WFSngA0yccXf3jGo9RTL92+A08u3e538BCJNYmHZgCvFDPrgf3NvtCo7
jbu+Chl2do7tmiR4GCS0JrpCmkBI5PVWLPxF8QiZ9fK+uMTxDfADUqkfsklWarIS
ocxhLAtddAKuAWsIV0qEuaDn6GG0Zap7ieCap2rDmJh835fpLqHF0FKVqsBpFDW6
KAmMaKMiWvDM6YzFtbx2piHVho28LBSM1nz2AD1ATCINPrgxIa5gFsOwyoORTZcS
0ezRpOISESllsAB10asVtRiYxdR1URa/D33HVGshboSjibAmwPdvpRvJ9Rg0RWjB
FWALcAlU3Z11GRG4rdINdWpozmLyo6dveU9rADqXfLKJAEnnTOdywwnVoIdG91np
+JSQSiFjXIS2OpUBK7d/UB8FGhIYD0zNKs9cOm6pmS0PPd2iePZrCmjehXjCwY/V
rcmKy2BvrWcfyM6IzDlektjOGE06cuqWQ4TMc5WRrYV3t0S3hmgIJATX6VuohYqu
wzyTGELWcn/KLlMhDVEVwJcpK9HgRL7pJGafvGY2Bx4lu2isujyybigfcdmuqt9M
F38gVxT7CTmQV+j3snOgDe/AXLFfvMzjXIc3+pTx0p146JlSSLec6OKthjRLEam6
QkuUy4SpgJ+p3cJvBH6Jt36n1kE451EbMD18IJunqRDw4cuUXd4GCWRUIFaWI7oY
ouEJ2LwQXEHLVwPC/z0R3XdQkdn73glVXXfqK2/yRvoWGUh2wLl0j2OfD+tRL9qw
w/ou+bXv/ZiEGRo9Ghycrfipl6yEsVPu6FEBKH5ldrcl7kHjw2ujTl8T1qIBES0w
nJUgYiyFLqiTLyFSJc8xucLMalPKaec0opG091FHeONVzNPrEy5EEkADk9Khb9Fx
tNh7D9IR6OxLpRgphd20uSJx7jmnG/TTzPOdbcfx0dpZ0NH5CZUnNErP5Flt0UOW
3yzJ8weLfGw5iOfV+mMRCIAAwJr3QjpLnjZQmvd8YBMqjL3PuyakQ2uB19Aqp0EO
HuFiaSXEgXp2fAofxwokGw0Dt8xSmbqNPnnvbfgdOhA3bXeGslRRiKubWbXlgNqu
96uhmZEALDSMBzaxFZW62dxBjOYcm8s+9WzDmJQicfQOXq9umvpgEC7sqEqLhVc+
292TqgJPa0M9G/B6pJeT1y3/Lxu5c1xWXypRFrqWq4My4L5W0vtELDkhM8yalmzb
VK2voTVTArKPr73QK3Kq0ddhPg76uTVv1BIeOjYypz5Tc+KxR10pf+vkupxuGOjA
07tWf8sWNOtvyv9l0B+zWdtmiXUK/SCYlaHhertw1tRJG7n9k14g7hYqBv1fsAVS
ktWq6m971ZIWSsqrWk6hjTZplNdt5YwTqE2mRu3VfvyfNCgrn+BC9SEg/gv4R96x
ka8jfVGNRN2U0dNJeOqU/Hurkcj6oj0O+USKYXYAOHVvqtMIkwFqwHcYVmooLxNS
WlzsGhui/3SJodysg6QAIZZuFvA0t45ktJP6UQ9gmgkkid3Ys4xwLbKSkBGRlToi
ERcHEM+nyf2Zv+nTqizQdsa4ljmj2/vaPn99NOUnXNK/koM9RZmxLZiY40evzYmi
E3qJG+AhoI2sG2rDN7DYj/r3s96ETWGofv+zJAX6ubpGnnVVQ9KyV2gOUaOxnUJW
/qnqB0cN66jvQGg2LyhklZFkWw48yPZZMXBqyXqcM67CCD+U3jszRGLHw/kKHl1c
SUVHhkZCqAJYPM/jVds1oXcBTy8EBch5VJXGqfDYGgWkk6lobNINHUmKovgH2QdW
SwJxGd7L0OusWSq5975rC9DAaTBgtRCzLmbYO9IY3frmMB+gaJCBXbbPRojbG9/d
s8q+0l/RmjRyYxjQs7PXcmmbHQk4V/Msm6rYqio9/nWaXB42RvkpqmA+/E/jAPRi
KVW6PIoHJ/SQgKw5AwPbjFLfpmvcLX0wagnNqEH7wcUgEQyCvY767KBxhwG6ROwo
KH12C+e8whlJjZz3rkChP6s26V0JbE3Hzr+tBqqgMna8gzV3Wm5Q2R+NFckgDW9w
ugsY8oNSNcj5KpYOA7BVE6C8fG2UkelZ3fJoL5yZaMyJyAwV3l+LzlWIcN7gEfrT
Z0D640bXkKnTQfN+X74NtK2SeD7eicvLILGNlkHOAGVnySccR3SvYXJRDv9i7Q6s
dEy7GwtM/LkKvf47E5itmmwQ+RBAtL9kHa9GN6BnyGSuUGtPXI9ccsbu3QW8zNp4
SnLZa2YbuPYfTAc8BmQySxP7oNvPQKlomjrCdgN0gaDYHkmWkK/dq2+Cf8LslkER
GND1EBKviVjZFXYpUMh/3Aia6CKsLYMjm+fC7zYYNqje/yq6ubC4WhIDyTimajnq
SzvRpjgX4vDtGLoNsx8c2CRlnbSQiHiJs7TW29YGDA8ztXCV9XeFk9jYswOAbDz8
xiIqoV6p3fniYaZLxtcUTKIIGhj6kv0eY1AKe4tDY7I+8DPTj/4/hRpZjRnjDTgD
giSzu76LQx62IjKZHHufTQVQBpEffFGMu9Dfb9liGKhcYcXvnFzT6hQJ7iK+Ez47
amDlFvbHLIONJMoKih6eqNLoPl10HQ6Rkppkv7z3VjHI41HWKSQJnZDEK3yCUg4E
TmQUBrgduK9CbCEsV6ZaDYuXxGb0nKaN5ujmqLQnY0hccVbBbyDBpKbMw1DPt4S2
amnx7pXcJUNbRzxL7gwLwP71KcL+wMkK7+RtLSNskkSNkZymhReE8tYzQGF0EEYs
z4ec5RZ0kWhs1xks+lFR0zEwx9ptVNt7p3jiKiBvetZzypOJOYYNq1oVH81P5syc
LwUDXlFsSUEtYYPbG0anR/WqMJh5Hg9likeYp9uiGAOVBdY8Ahy17YguvrGyrY+E
YkNzVtYucjUhR1bk1aF5nNDS7vPu0usutORvILCzP8iixSYzRD88+Rbz89LG6w6e
X+tQEFOqqzAaU9wazChUbXDkcd8qdHXs9oDAdIP8tobj4aE5xPEublVM9uZPpNH3
QcB2k03Gtx32Dr/2J/RoXy7ZtjwsL6afZ5zwN1LymPvurZ08I/pIV/ZhvZ2YJ6kZ
y7RLV3HMJ3SIza+T0vH47qeiPOkTORtP9k6N9AEtr60Ocw9lKfYLMK0n4z37N98f
Au8cAS3vt6hL4MqNaRFcv6iwEoukOe+OKBXhY5yTCUi/pG2KUKACYhTVCRkI/r+e
DbotaKkCql5As/L2mbGT6cDEwTe4KlyUccqyakaENJCBbZLzhrfMxfDQXtgpRF+A
jp6BJkQ+whMe1Ync03PDvEu+Nc3kdBdriPcExWF7BBsOGrVnUp+6PhXwFHVBZAbE
u/YV7QkhdEjFRIOSmMOqCzjXasgGe8jq4Ss+CiKYwwvNFJOwsHUhZOS/DgCyhCcH
zyhPpG0fH3JFZ5Tn0NUpjUnpJvvVs3UNaawCdDF7wNLzsBNuByLHeitcwWbQPhiZ
wC/vQ6of9rfS7yNr1ta4t6q7lOBnBZCCGJp9s0c501Or7RaLGM2wKJbszJmhG3/0
Sh25BFircov7RhLIdE0djJP+Q8JKAeE19KbLLCE3v4VrINQarMX97eETqus7h14P
gVbMKtrYvEvd01qRZlUdqRosYtweK7kLzPUmxGsaOz67d7EFeVryMEH7/NZwBIuZ
74vUiEspMnAtTXeJHLUw63A2UkzYtOOP1Hr8OwP0IiZXGTB+z2ycSxGDF05TTvEN
zlUWmwvA+b7gg+qBd+OfxxGSznQA5vUcKIQYzUqBYRTqic9HZiZ7YIU5qO2LYnP3
7Dbt/thRUfXSOWEpcHiDNQAsDHXfv9AMhZQeE9TWrRw11o7Tb+4fEQYXqPRdZ44Z
zrOEebtfIGcB13aTLt8SMfvedgvTfL6l0P0ZOhXdV+0qMLXtJM+NZzWE4pmbbGN4
pjYi2SIcaPf20IvXa09yQmLWBpHw3uINlFBHFC95bshDS0UI9uiBJcDaaoh+ntVA
eYgp1tCZ0aA99fDZFr3jD757zw57+LMxw7HG0QVb7560Ku2L697t3IhPjmuB6DKe
wq8GcvUIQzYXdwhQ40s+KjomVpBOcRBpVobDPh/vro/Z0e86b4ZX76AZGOtvICUx
+bXYROS/noPY3Y+G9VZtqGFmt4BGZPJZ3gd9MBpXaOizeVRI7qMSEB71fuQlYjV+
8JrGW6nTvkLRuiXu6lWb1JfGiZQJpdvKfvZOiGR9uMYf7LRHgk43QZxnzm96qF9F
7vRaNeHmTqWkcTzSe8ZEfYBCJsw8y1LK9J+r9KUoR3iMzVcmMr0/bI1CRAVpZuXt
ifMzv3u61iyeyU0KBzNHLvQFnRWGx9fwakVeHfH0L9JRsIEzguJUdVR6PvuHZSrP
7mAwylYjO3iz626sOfmqjZJJB7NPv5JwY+4T/cE9Nh4jl5emSgZr5TcrqtGDlcL/
MN0GmkSEWjfQA4RZB6A0kayF+2K0S3yEbqJup8DUv5elk7IlUYSRu7zdF4CRNLYg
qZ6j5x/kHKqIoCwFSmKfi4cWFUjBzZY2T6lJwQhEKVkb7RvB5TeeJbLM7/TjtutC
gVPM8Mi++jU6eJxEh9+r4yNILPrBEshKXasRmXUKidSrJO+mJ7cuofilqKwZCnep
9yfTSKLfPAkUDijtHyf+U5SKSPeC2Y3tLaZ9bpIhpdNvVPohOvKYDgeKu7A4F1tE
X2FhUDHJG7wgyklys6MxdnYn6OHHHHkWE58PmL8v0VqTKyZebSWKVHFwJhK7xuxP
FUYizlxge2/Gk7S0thiDe6Afz/ZDBfHX3+5ZYa5q3Y2LFS4FIWSMU8uxYSwnRycv
kok4rzeSlsX8+701RwCGU+NRhRK08qUd6nwNukd8hyZ9jGWeerNdlncYpPs6OWwq
vui3vOXv8RRShzNSwDP/bbsf/Ur+YJRbvZ34I2ZdpyeJKpqhIJh1GM4rGk0lCidv
U95u0r59HQvjiT8rp/XvwcFyzox3wfF2hAAJ29GjJ/hChQhRKGMVnXJ3L0SfQYHb
OtHsy6Vyn/y/cQZuop7C4zNfdtRGTb3MF7g6Uvozmqt3cGnIz8Le082BkRQB2oig
b+0+eRKFISSQUqUnBLByWDSPtCYEpKXNnEQnoClN2YiEAlw7ScaOtuFVMaeNavb+
yiPJSf7r+WBm3uJH/R4g03SITwtgCXeHFOB149Ic0UV2pnC90sdt+AL90KrbPnEO
7ZTSClT+T7K8TwGC0GPbLly1gsCRGX7deWTv0ikBOVATXpp0pSCK+kV1hzfMDVwZ
xLdCODPg7incLeEExQe9zh+nRuvLjS0rYOpvXx0gUs3h6zGxszlmnpeVdSyRJaXZ
ap/yjBlJjq6VdOH08TinGvpehcVyzLlh8yiVuUpxQpX7bDnARPVnJ68pha9bHc27
aroLHmfcxwYGwdjMUWTzUQjWc6UW2SEEgf2YTsB0yUptM2LB7aDIHia4B1Rl3s5a
qXLkAWDy0tkynMixvRQxzTpclOHuCDfaXTU4SSMmCZ0XUJYoQ3nCvxrcvp6YvOtK
76GOs1RdVbRYguHpzsxiXh3qQFdzyvaDtd1Yf6RylhkeIzhO6Do4LY2oqIl+KIm5
E9b/964zrh+TxBsVOtkK0Qz80yR9cRACUGLsodqFz0WzgXO88yjOKejWFwyfywcw
zZJTweIT6vjRjC4WeiobLnAuJ3pQ5L3R4L8mCy3L+cUjWcR9MwBqHTsIvONg28TO
AE0+pQ9VXwUEBXIuFDV86urTL2I+FYTBM7gWEbSMKH/9SKUSAq5phU4f8DACHGpY
OFlTSYBVD2ZkNxkN8Z4IOlb7JTXRwMpPxjtgY9ZEYsxiGiwbe5Ju6UU/VPBbWIk6
CC1/09h2dyxCthoTWHZywJP0xXsjCzZLemKiwv8JfTKLHRRkeebqzlzn+A9Ry2Fv
h1D1q+0eWgLtZBVHaYcIbLCB06XC+C5hZY592O2KpDlYpgaUMCy+YspQ21gKybMs
QZWU68X8PxNfqiAlOn4NaDfo4EpBgIOu6vgvrVdVsZmgzhAcwkfYeO9b48nIbz+T
SjVHvlinTbdm8+Z2gGCgR2qW2n4D2H4CHsfpcBX2XBHGQ2BkkV7ks5dN4Y0kRxp+
rsLvpPs8AS3pd/BvlkwZ0M38n046xC1ZI+f6GRzgA550OEpo/xv9g+sRwI3r8ZIJ
5I1rYPKzb8likE+8DLMd9gWmdXxLX7CIkKW5tgbpYGveWkrZSbcWfdi/yRm6rGsH
qTNmnDOGRyVDZx+mHa/7x3cOv6VK/HjDAT29m97BsaYD62a+S7b0fNjoCAL8HY71
FRdTIpjjw0BRTDuGYrkfW32qFFvfN6H7UfcOVjYvuofSs9x059cIFuQm4v22fwBL
JoBRqOjvqoWUIzj4v3raMWBkt/p608kK3LXDAtWZDC+wMEXnsLov5DkgggOJoJy1
lh06c4SQlO15jI0NKE2oLjkeP1qV20ScslLJgsIW9bv7McHOZvNltiqAjR8l35UX
Eosm6HIciP3u0+3lZaxzOxf+8REamCgHDnmQNIYELb8a3L/r4VhoYfHas3I9qQ14
NLPL4hnsHOSJg+EYhvy6TztQt919RFI27eDvu4iJlwpD3Y5r45Fypo+7jRvzvZIt
7DkwiOfBNeUq0jv0BLgquGOZbJ4Yp6SgTpVh01knTT6iODURfE4M/QHc8e1/gLyZ
TOZoKQcz0aGZrJlcpsfs4rrO9LTH26jKZpJ6lqCDKGr3G5XwEXoPVq71UO8VXNUn
+SY6cmPHnpqX9Slq2vJel/RIZAEcquVXZfBZOMoIVNusawVbznbOrAj5PKB6KHOU
gEob8SfzcB2/HpZhRGLRzeXLGF2qOHU69j0f+5MPxfmWriMBgXSnof4hL4Q1GW3z
YjWtz6HbUOirzdGc7RHmffvzDa+Bt0tUh+8crRBQjLu21ogiccxOXNbpZRrtCnyZ
0VVhtSzyWG3Yuzchb5Y+40Z/SRw39TeDaMxVghMTcHM5jZrm8s0XRsKfPAmSo1eJ
x+arHKZqAO2a3BWDANNvSie6LGBL9gkiU364c+l6YweZ52DUzzcgG1QMOlANk4bW
2CD/5p2LUXXI6VntDMAj71KuxhemgMzmeb58Vct8asWzqjSNEj8SVicPBglZ8X9t
p4CXdlyyaaSOeOX1iAsERAZm6kNJ3HbA7jlUo6oa0LzfW1lhKkXc5VQYicA81L55
6wZoof7dAhF0cTjDrWGeaBmmtgVvTGSbVoFPJvCFTOpApu+RTzvDqk6WcRTx24oe
N7eaJrwuQUTLsJiP6bY5htunX28jQs/r47Ew4ul8NwBwxz2uMBty1lTbzXZBlx4y
iIaFeX+qyJqwutBRWdzwsGTopFKZpL7Qv5Mo5/i8JkGSDrXIRFBD1OM1mDaHhTNJ
RNT96cxtrvphV4ag+tEvRxviNAHl+Cl/oRNno1iDjfQn0E5GHMmPS635Av5pl5cj
O7CWc3TK4XxCP+3S0aK4dxtEsKChpkS/T5tLXJY/hx1p9FMaSjqfzxlOtBhoHhl3
9n/I7GKNe8jrCKkyLWf4ZFXUP61N96qaBpB8qfuFVN+SQdNTyLa6s8acR8zG2nfs
AAuqcuEuNY4TK4eGZwuGYGFnxE23zMIxiHJzkqOwKQUZGi/B2ILNDxFaGan8ZCdG
tmqRmb8rfTdxkEH1gvO5hOczPqtJHVY9fIy5D/vU6rW8EQ2uOOu7m0mxUsgz9LFE
QwOlKEaAh6om6PMCHRzhrrxe2RyEKCABIo5QWaItUYCELsklRtVvBppu6cOD/ugm
jOzKkZrtmlN+gmSxx9FUOgMv/pBzRl6OU4yjdc1WXGAO6AYnMAp30Lxde/Otnm54
nRVMdnL7IqFuuMu/yjOsvls+MoMu/okODTdTllOYTY4LNkpYwIhq9mWNwyB97ruX
qKIemjwX+xOHx0j8KbbDFLl4+9qiB3oH3qkxvVwox9kEOTYKYvgUbPzoavc1bomq
LrFlKBLQqgJ1P096EtA2SMY/+UXT749K2P5Je9ouR5L7U08ZhHlzymPS12wQgd3p
h8RpkOHiHv6HPfBAAaqn/7JXd/oX19G2GvlbBTAINuEw4EVJE0Oinp3mAYtytwz7
ruRLQR1lOR9lr1cNWm9v4P9tyu8Jyg4xbM4O53RaKp3Ac21QU+UjMiokWQtHSmp9
h4dMEYi8iw66L3POngV3T/X9VcZOh3WYvgTs4TlI1gScpxvMvS1pM8+DFwJAZQ42
eGCBGlGoElN7qxv2RATJKQF40JUZkXYXgNi1BfBAmWZaFfXCwQevJLsrz2zaAd4d
5XcxSlddUyBPIQ3+8c6uSBBN1OGP+knIvmNR2HYj56YeFVDVK2bpBP0Ngk3Bey4N
+vt1WFwd96YBw7ZK1w5SVMhRSvMaa4C4J5FZzYKj8+CgEY3AZ2XodLelzuvBivp5
h9JCEofYW3aMqdAdmhduKO1b9UR7saAjcgtQRIS7GVv006yAoDE9YkFOO/W8AAhl
ysqN2FexIbQ0s8Xx5ngVt/Dhk5TD5Ju0iTmgrpH1Hi9ZFpfVGVaHKGTbUqsfDdg4
RyR/RfamwRVz6X2b1EdahIa+SmOZJwLidXbqTv3bwWo7MpkQwSOhV3g2P/+tg1Ne
aAvumoGVJC22MG7m7eZEDvm+eIGiPVv1cipa7Z+Ix9/HRfSKJHwnNto2UnENLm8p
lKXER/yhYzBKMOQjGZKiRgg7TE5RdX9f8TJNn7tqAYLH7eaHjiDQpunIpt8H3VnA
rGIq77uXTQ+Rz5e77gVgtio4EYPXMtjI8JEd0DC7Z6T6suFB7uz51ehA7+5zrRF0
VDGTIPGntrahFb8M6Ihi2MA5R2UFOKead/phye0f8TMZNig7Emr3Bs9AaBgUWprj
buaQICoK0tgMd+biVpe/xbrYwrj+uLLEphir/SPCUMyLxXaXRhtIiU8g9nlhorDX
ifA13n585NNZ6R9RZTUa6swfRZu7lSdUyXNZcWwnkYVKQV1VEPXDMeOajEfQbrgw
6qJOSldM6QSnrY2ynKxwJNnsiKfKsaFrVWZwzRLEMXUoenT5lDd2riBPRfGYcIOp
7qlQBuTBXc9JtQXO7Ih+n1AMuvYgx/+FTVRxfmXgdOLwgU5xgisY/rQHDAnYpKlt
fjG6RRf6InEa7k9/lYWUQsMyTUtbibyeEcHQBhOov4OWwoVRkYB74eomcaF5PlEF
EKXEFD0YATSp20Ut65l/+pGRTafTbUnOrg7yja97fghDacxFOPQ7Mj4l/9sJWtuN
kvXxDrl+mR+pqIWMPytdGThQewcKwByv5Z8dR9uKVWmVji9K6aqHhNRqjse4GP69
UkKmDpABwyq0E74z7KrEP4Nz+p1K+oQqF9c+8CoTZ4bCYi7KKiEDDACgCRqOzSi4
16pkg7lFtbTaQmvMp3oVaG/Jg8TVWuxat3meF6rX/3wvA1mnGUk9tvDQPepqsw1/
uEbSBtaHM7aIvnZxRZs+3ze7+nFK36Q4w/3ilZREDmYgMt+mBnNigDIMZ9JBWzZF
UWwzCWNtIScmy5SvqYcETssLPivRMZf8x3aUH9CNNJr0BbPiWO08wxvohbQO4v1I
5e7YQcKRfMuealYx3jOdBtx4NT3ZGN7JS+/wPPOp1mUVVujVC43ZB6CSn7An5T5p
Fpq/f8aECV/oE5Fe5KNkRnvlt5bM5AoQ/YvRDeyvo2Pc3c22+72u5CaNO4gQvNib
E06kczZ++JSICwtvInIYRGZHSpNP716VdJ+r7bc5AA8/uT4yDueEFasTXIZWKRLp
IhYmuxMi9lUA15TljwbKjrZ6HlJ/6FDROL+u13X7H8JtMAplFHCEtrameoLRvYKk
tufytQlAG+KzOsX6lz9gI30kv5PkOufrg7JwbcdW6SXluAYDZ+CpL9PToQ33aNEG
hLoFWQLkHQJYHmWy19nR1j1OSl27nuDoS1ZKC8Lg1/oq2pz9eK+mMlUrmC5n2paV
tQ8RVhVshjEGYERzAeBkG7Z3oCdBqgeb5GqQdeUwzwmY6qTIboCW2Sj87tQKX3nn
XsdhwylaPfVW/NenV+Vc8ub0L/rB994cMhqE2UrpT0EYvolEG8Ph+lrgML1nV+Ah
4vSKt7ZVSKhv3SGNN40rf1QshKic+bwOA8ceKobJ1ba+E20SHRxEaS0NBjbW38Zu
H+LIKLBm69SDUDzK6xwJnK39GsBG9DiAg3EPGuK3Qkzb6EUdACSKWBAfolBi6LWq
F1uyWDsMqh7kKL/RFJosoJkaeeZtypiH1Mki8mK3qc10SaNNHL0uAyR+JKIdM2SE
4rzPrIAi+pS9QdU118ZTQmBfG6tj0Ybtv+4TzJZhm2B00YEpD7tQTd3W2IvVAWG7
PNHVFZhrgp2+PZGHgo2vBr5Th3h88YmzdZscXsnIB5mXjZmMWBSkW4QTJeUjPS0d
CBezZGiWi7uP+eBlTBNEV0RgvVIvz58vd8aSj/JzYLb28INfYotm1d67cPEXWuoh
uTiDnRgXBCvUwnDy3Rvf3JR7GLoD+aRdfp2BpOEdpe3WsoHMnHeQ6jlR16pVQKKe
FaE3zGauW5W2UR29OiOrkhsVuy47w/MThetCSf/Nynf61u48gjpX1bSfs60g0ni1
EE2Q6wZvgJRSvdKBlCis4Plt6nJXCrsKXXAJB6Gpfg0zsoGHLJFYXpdTDvzGDgbl
Mfa6SLjfxlyz/OArZV+sivfba+pjnbZVu6EQvq6Jiap/C7iqNsguqd1ZntAeVswR
8xhGZVyUZ6H8hQD++D/Ho0z4DhM2K7cjmMjGnDbNuSUH6rf7ow07XQJgnV/adZtj
ANh4g3NCYq0QAJtEy2k/Wnje3jwhZHlX577Tq2f9Uti3/ihJHhkXqwP6mw9M2S8n
yW7s3DkGU1U7Q5xo0i3KhyKeeQtBo7QIKJ3DaXbzpAjdA2kbYxBEJfM4VHIU+qXv
mzAS64CL7yEQTLl3KCBzx41Sq18ah+p8BOSXT3Cd3mKHvQMGA6S8wP8c2S/PoJ7w
/g3B2lE1nOZApAuDz4OGIYvB7c8lNfmecAdVTis092gwnqbmMSOjMFEk4xlLWS9C
HuYvBWd6wsw+iq7ldA+LuZP7irPcq6OOl7+8neFFps6k+TILTNGrBfrCceN8Mb7u
3N2Hsgq45CJg1UoNtDRfcoc1VksDW9YXGzBv60GiUEYPelboG7uWvpUXMfjg89Vv
CkAV9S1DqIV8mcukH+do4gfy0FXAsqgKWK8/2ko/4GvSjob8DuQ81tG2naCdNB1O
WumTONrAUihkCr4LxsoJc58mHA3IrR+9PhIh0Ue7TndcSdqTh8lrLkMfSzYDCeEz
iX4eJxYxtEoASE5Ayd6092x/lzBF1Mm/PZ0RX7eQ6w4Memebb53JuZHojxWvtj3A
bsxgaduMPbFcvnlNvPEiky1K5+K8eSAKHAgCTZMX3ggL+QgeHplnEyH28GuytOJZ
yQIPXS9nf7fJBFz3BgEfKc4fSK7DJDuNBGd4j5834vIBokS93t6emoLI3FxjJPDY
NJVInmd9nmNEhXVJROcFUJ18hSg4BArFJnPc8vM7PhW3Sh0eJzpLfUTnzvnGchGI
I2xt5Zg+c9qt39p49ZW5YuI+gV+VIwfmWWZxj4CmoiqUM0YN2lbYDLCl82/S3Pnn
DPxGz2/sas0duVlm8n5/L92NVhw9xERoyPszb94QzOmynIBI5ye2SGJd/IgvwuD2
CdJlnNpja/GBFHXGN4XYdm7KY5MCIy+oyNpP5SCtyJXrPBIHMxKY/xlRhs6aa0Rz
njw/Cdxssy5ffcpiyxRcrWqa+LhjS0Ud88hAoKO7xhIDiQin2cudaw/BAJY91kJm
GZxkR5XvtlBkyGIkrpH/dTG3c0vVHpeGFyXab8DFmta1DStBZ7cYTFUSs9j36/pk
nVL1Dh0PwdnA7takxu3igVZnInPKRqAVVqoP1KeUDP1mQFupXjZ44sV8lPu8jV0e
6Z46QZCoNv3seA77k/IHCQY+c0qQKR60y8mav3rsCoGi5JM833heSyM0JYXktkFR
1ZltPOdndhVDDq7naMtsetF+0DIC91PUdzj1urIAW5MHgNMY1RNa30OjCyzGbtd6
VJYwZc+ZW4N4wW94VS/Ih3fxG4odBeeReV3d3km9EWFyLgbQBySh8pFvpK4Y6Z+8
UNVO+mzys3NGxYN582F6BBiSOGUmlrUJDT7uExARBVfH5Xze6/EqyEb/CDnkclyE
JQRcvhT4eI5QQx9otr9TN6qUF3TBogJrHylG/07cNm3Dl/YizQok1s3ZgTpDcAFS
l4uEv3gRxP7uACroAzqmJLHDjkSJRkv02Ivay7Xx1pO59BKtfQchF64oAiq3uZP6
pf5jruCw2QT4+zKye1gbczFQ2mnioCaRIvvHpb9o5k2k+hfcUZj5ENbrR2jMNG+P
gVFUZG4c7HnerPPg1qVg+C/zZneBPdOqfCeKiyvm6t7crkR0ouEX36I2I/hoPLN6
eqaOzp5tMjngzQu/H/HHIB+jUjyBtWYjItYAIuw8mcUoR4mUH5/CKv07dg7OMuJO
5gyMyiW1G8ARHvindP2E6TJA2Ao5zC6luMDdjYgAwPI7T0QHIRoudf4P1GRTilsW
6BQWu5Oo5sjzJYzNB/s2vxWS2fgiYeIk+mfKtIGl9jXsq3NGxYUZVMwqmrjsB+Kc
ByGXHcRrZJViJ94NPi4w+e2SeY6sYc+q31uLr/m9cpvvAZs/ovZKKfoLf841cfhi
2asy4tkI1PmMVsPqgsYDs/DQQuGg/wU+o4r3YRmcgcVz0/8WAOg+Xo4pcLErrsbF
i/l6i9iCK1pPUskc5H1LfR3IOJsxfPSOXKJhXu1Kb1+ilufCExg5eGpZkLEfJvH8
93CPgXQMzvWQSXYjZpXG3S9JUp/cFyQjn23kPwurvaVCcPSozXZvXagRVwtqjKxH
K89GEAhOPabhOQCXMb/NwDs3QUYdrMizKtVIsl0rCJvmmSj1nkTqoM5k3sLFCsuy
f8Kyb5A6Ld7VBqrwyh6n07rIvTCPY2huRaaOHTb2fSJc57DK4DjrFxtl8KWa5kfT
y4t2tiNHF5eJmc88dia3mMq3gYlTzthqrJrAsarMwGdro3HGfraBCfG3dGaVLH+Y
ORPcFFBEI9AfbR1KZ45LJEt47iVxAVE+8WjChX/oN5VDugwOLWpJq8XYu3TSmL1F
ZsD8jaie3POJRlQzTw0XI3cK0Rz/UiAW2yEUms736DhIesze2Bw1ONx88P1MJ917
Cr5gWzGjI/mfKSsbP66ePPurUWJ1tPn4x7p0WOdtT3Ce0CHanLyEJhoxhqTAbOsH
TwuMVyWZn2j4LSsPuZaQAXKQSGg1xZBxSFwDQC3UEZspGygz/c4s9vyFYisSGmkF
sCTlxnvuJhcTW2hoWHFXW8ogYvCeSOcdLzwVa3uGuCSJsKuJXrEr+UhsVXm9Tf9b
xZRKpFPjK384HSi/s8tVUkZ/i20vVIbLAIkt2V8aRsaQeHy69jZj0jwtJHF9f27B
KgcbYC69zVQkYYBi9cOUQ++xIVX1rzxy7wam8mmVw6Hqts01KrsiUVeOdNEtjLO/
EsjNz0e8enVjTGKB69c/Un+kWzrAV6mXAoGvQhV7k2F9fCLT+ZlxZV9eP1gHEzCA
0TeA9qOuoTE5TXE45U6focZwwzj3EQkIll3I8WKXz2LLNOkw76kyTat+iL1Kjncp
rFbUvLBu/2sD9F3iSwjMDFcuJjdpluAgBJPlIc9LbIht/rqX5T4nTxhQkJ4q8qTr
5ByFLrKEHe3enFtdI2sESO5oa/GPN0ujasgYXm6nn2FcLzZqi5BctjfVTj8p08il
RtC5JYRNpTEIhLw4+B78KR9ShbJMYOqdYwoFshhvvtcaIe0wtxg4ezapj3nBJnEH
ihqgW72XvU6FRKg1+/luLdZ36aQqkjdubOLxtr7nUIRzOk+SY3ONPskBQ1rXcOiQ
vRIKnVmXrdbek+J8x97J49t77tR7Q1Jm9xaXVJz3xysJRS5aXuPRXswhXPVRXVmw
tqULhUWcsbGdHywlpBx+ktNkCN1h2y/XdNVPjpWtBY+QsIUkWB9uocqQARDNMHh4
EzpmlVISWEbOpaufC8fbSExJP5uPQ22Xw1+NubYf/BsTHCdDxkeSf276z1SVDhYU
VIvGK6Xy5/MHm4eySucOFw6ZWXr4EIxmgHmCO7iLi0BQJtwBoxnTS6IkHyE+ecdP
taI7HYwsFO2+6PJ8xZYakwCZQ2yaxErsCeQ+SH4mkFSC/9sVb8ifE2cSeyxNsofk
DD6imtIMqagqv60n/gZq7g1CtbHd8HwozlalqkemLV4lSIGz8nr9bKrJB/sUi9/E
UqDD1YajvNBZvo0AAcaZPv7hfK5FT4WezDGzg5i6Qudvv5oijOqcUq6c8OYs4VTE
PprZn46GMlT9/WJDT5owN/fdqhcAlMwm6ljhjRoP25naoDlFltDtSmGI+Pdvqa95
VPnoCWIblQhrInU+rn3RO/anGVL+9GWz5imJpJQ+zxfbs6a7OpIpe6OIekvgVp60
JhENyrsb7m8vkg8Wh4/H9v0riRihB9WiYM9IUxVS2ez/ZCsD89XT9q74YDwYtKhH
Iceclqlu8tFQuw5NdwlI09dHtJN7YIhpR7azvbCNd2lHwmUmcy9HkoKqkgFjhrkm
lBkG3yWNwDf+31UovaS98sINi0jA9YEJsPQUYRdtbQD83MG3UT+amiVH+VUsTm+8
RRvpoGXTRgpLkyFj3q7eWc8WTzhDWgZ3F50b7xR/eu8qfHUR6TA8Ga7Ji2aIP4bl
HXstS5nxkgAxWawf9Bbu9fJKQ3NKLzNazZeeXQ6xaspZDQmEodZILrvNdmbn0k72
xyWJmg2M0uIqObN969PcYbFz7tz30193mz5MUX+S0uzLidXpMtmNgr/gb230gmlo
x4lHCAs+e9r4iHy1zXGqI2d3hSNBBFGHIlfKNNDA0RHD9xrUh0Bmh11+x7TNHeau
KBopYMjt2FmyJzcizDnmHN5xVe2jcm3drqAQmWQZLDFSHTQPa/DWizP3avt08chR
W1KlgthNZGn2svhKSumD3ssG00tPh1FgUTFhtIbjsRA/dOEYf/IdHNNUCCFBaRP3
FhXQsZF182hLdAs/7uTZw5nvXW1jCDU/pfh24EXlaLFXNN0YsXfzdfGbQtXar3mF
l8Y+w6wW6EXJ9n4ScutiXQFTzlpwrjhJTaONk2ZX5/0KPHwX+YOhRKDzrCJVAsU0
o+mjg1kaCk+2NMtEEJuQL6dj0v4tJ8QSkqHQKpzlNjAfrmBocI97LWPljxChIvK/
Z6Fml/n9L7WHqFH/C7z2xNUw3GwcPi4GXf8pEW2/jfnEf230nM7SqEalPD+lsVqR
Q+xw1Aj21IbwkWJkB5bS7DzlZNNEt+UbZ/rY/oyyPtERmE/wfhZCN6W8y02GxoOI
YA3eZy2xKp7ww/fkVisrSBv41tWHNh9Jhr3bhk4cUNZJW6ICg5L7e8nPbpvA9k9A
sLu0CdCx/pcnG1dphSHH+RJdWC2WnhYfERnWX8C5lxhHKLnOt4/1b9Bk3s/PPNCJ
8KXiTc8UyzT+c0aI0T7d71cUEG6qqcQtkXCHOz54aLVdz4k46wfSep50H4oPkVbW
S3zZfamfQVGzcbFV4u0oODX4xJGpEx+o7SEI7yC2eeIgbT6nEiiyRJaVF63KJA2N
Vs8nXSd8rLdTpsEhfMoXJ7BYIpCF5xP71N2EaNXVxdNPdJK35B+1uY34E6/9ffwP
QW1nnXBSokzW7Ce96mR1vHzH2+nPDQGkQyufbf5ZD5BtWyDDbZAgMxixiKMUy/7I
pbjOPPl9vb7K31gQAY5cQYQIOzIj1g7v90u9d8Jpe3OdJ4KvI7XjsYyhKeRkpZCk
C5d+IIfDbh0nhBVsMgC+385LJ3+5DflcLVgQ1kMtJ7OtJtjLMrhg08Jsqwu73vOq
exFta9TjhDx7NrV/+aM9Qua+ikvHen6iMkzHLwWzFQLOL89VkDXmuwaaVvNzErsy
EwgR/uAQvJhK3yx9/BwQRJ0sSn208dHdBMqFbfvAqLFkz6rv0LNnb6gI5gLP4LGk
vW69wMV1IMkZ5mSvLZVOWQ7lw4XKHWN6YG9LX0dBL4LSXP0dnGF8ZLfSuvnoQVvc
gafUhGFdqPI3XnZtncBcpKTkBw/4kbeTHXU/5RNLtKDfwZHyiarXw9RglQ3lGbMC
E7jnmDbE2cJTNLrpteaE2DBsnwe1dSk0kBO0GIr6UMa55PkEk4hat9Nci7f6aea8
NvHpe2xixgCwplnsYdiWQyhoBtEEiAQseCG4/Cs9ULxv2OLW7bQb6GaGKOaFTeWx
79WoUIjNFS/LQP1iMSLTf2J4IIyeJxPdM4ysxPfti0zG8NiKxFzOfu+1MUm9UERu
wdmPzzMMS/ZJUtKO6d08JJUhumR5eFcOjjlNS3RHKaCBw1Xu55MDAnmkv1XHgpdD
qsGly7u501MmzLJnBn0KWecOdN8/YJUsTcObDxRNWyu2VwmWGN42JtYOGOIGSYvU
7Ylb+vJCqKAhn+vTzPwjjuPkwZkBOdOLJVVhwxb1bqSIYLJO+9NItpkKLcUsCV65
tI/vpm9uxvPY+e5Lf0Wl0xulThXD9URiMdML8BfgXjEIgDW7vVQCG+1c2IJvv4sK
zWtPocDweEOJspurQVHSBka8CrBqxekWtCLA6/Qi9wyy1tTemnIk2scBrrc9YwLx
AsRBHm3qefYk0Pw9b7pKMumwuskO6TGkbJ/yG92P2LZ2SNenk33Ql74nuEwN6KRa
M15/7CJV6dZowR6I7Y3EOUfN0vJ2kJbwLEnhDIWonmfZiO3+uyWv6B0uZ6YUEQFo
ano8X3XZUkDQx57k5fkRv5uIJ8q6X1+V47E1LUNqDcLlUfV6r2zUmisOwBJYmJv9
KY49+2/55SgoIaoi+xm9WZe8dzYql/KL4S+t8dj7FUVdW/h9QdOlyRGadW4u/a63
yeXq6EVcX81A6hfiZ9eC/k8OkhvzBuT7XjDaraBLRscfaPnC7Y0QMMy5zuiVE+ex
LQ1bRpcQmiWYu/SWpwTnVmMXXKDpPZOlkSLVQqGuKaxrz2CjxvzWjthIAJJ2CjQT
Qf/oiAPUvcR+pN6lVtKh0kRClhpOv2aU9NsFTZDkfYYJF12I+Ll2+hrjL2+J6drT
37RKsBq4jcdAejy+lHG+w32lpKNvBNsPXaU6w8WvuxRkTPNO2IjpGxrJpE3wK5MU
VDu0Zoef+pXmRvkWUJcoETi5D6gxgUSIRAVLrLbzv9xsAPXXSBL3ZzUEi8gxsEQs
kHfoHs1ZT9pF7IGYYtVHwcBtLn84tYG6u0FcVivhALrjAldH5Z4h7g9M6CtS+tc4
PQowWniac1tRgZ9riWlKnyaRZYOgYACKK/dRAT3CR46KG8n39gTnLaSYGE2QpI2w
KHyLfC2c2cmRj1KUpwktvgnOBUn+orWOX/J1DR0XiX6UHDf4Q5u1YmnZS7/2ORc6
d0aiKoVtCE1MvPcuHIs5mq7DYldIkrKk2aBaNwh48Q3yvtXawf/YY15r3oJJgYSl
zUtyiQRrkWQAUlD3GswMRhntFxFdHqe1wuHhNgll2K0k5a96ScqjTeAATizBzEFL
YPygTgQ0RfVrJ0n2Om3rzQRGHQWqBz8q/dc8pOkiMtTIdBejT3taO6SSMZKJAq0t
emt0xY9FJUi9lLkZJ+3fJtdmF9GsqW6qqi138c4OCis2g+3sS37HK3Mr2m51A/9q
L+Q4UveR9MK1miKnljWjNaOSem4NY7Fyt6QgdmeFT5Gs+nCWjsvNGTH4zpxonhxJ
Ye0LNe8IaVyU5CQgJuWSCYXBLz7YnX+pijaC+c6ynsQiFGBZehTZAw/79E0wMBkT
KjupF8e7G7RX4LQqTbYiHIDlD/zbsgC6qtQ89bRYzOsiJ+jsjteF2MnAZs6Sm1YN
GeCY0QHf1Cg4/gJOjI97qX/tLwOpBfiI4DXhZWVbJjzQWsP/XIinVMZaKFL/pEem
DyRm2pDE7dlesC31qbQnesUDlAAMZ7Q/863NFHzPAcE2rMSt5i0OIW1vPqpjMk5p
K5SaDpOpSfYz/xjj8tfDkA/9jTGnM1duJaUmq5z2ECauqtFt1T1T7ZHYIfU/YaGV
8i/IYQyZ+JdSfs2uj8v82jU1OQA0K1NJ6gvHZ4jOHlcA0gApffYtOLea0TIpkahL
0JXpjQknKq6238hyRAn9mmoy/YLSwAJQKbnO23atLe8b/uyGrFK7SX3Lh3n/MW2k
dgGTIogbb39M9PzoQ40qyZAWATNInmHLLr2HTfzoEcWueYuaKH2u3ru2NyGOL9Os
l6qPMDYIl7OqLwjrxaml9OWp/FNak2i4cU6cQ7EIlA3jmPfJVioZlhIvXcEpo7ns
UwoJXmuPamqFTv90C19wQ0RtNJVs22Qc0UviqRtVxb/+uLXDBqZBUUiurqA8OWyV
bF3TZ2/Cz/wRWfipX5S+b5C734UPZvME6lYIuWABDY00/xsiPjESXsJ5VNR8UYix
SkdLJS5VEP/1ejvR+7NUjHnY7CGrp9B6Y8kJaX8OrFMeGIiI0PNZzLnz7A9og7mi
YXp6H2THo8GhvWuMCTSI1zR+c9UHgBd+srONHP+Cj4ag12UMl+oQWIV8RnxdsTkL
KnoOyAea9YPW+asOroEn0XFhDPnapHJ6keh+520EJgGLKpV94SMAJh3H/oWYJYv+
cFPRRUcQxdo2waMdNxc2qBTn9tlIPg8E4t72iiYaHDg/MLX+GqgKQotAwyOL/mlb
Slqjyg1uM7vIPJkjR6UPFPMpCsI6X7+OEUilY7DJ963+90HUPSInEW9Vzj4vADn1
ckO4i2ahqBAiyoPpOamHq/AR8E4HaupUTk/xsKGfTOKOWOttar+xpZ7HTt6tebgg
kJJL6sehPthbXbgT0bndvl3qwZocjLW1AU1Rd2DwtRCOgQr4zdNZaawKgRQvkm+6
GKm04vgRQLfKGz6QRc8joDUhkgDKpjuhH1JO9eIGL5ExMKGkAF7dMbM6fe6D3zyS
FhkpV0PznLltiAgYyzJkvwyrz773X9IJJ/H9nT/QFNPouUdXPGOQFMbz0QL0P81R
ttTrPam/CDiUnhsgOIX3/vqvriVEeaESu6dsbTUO6/zf6/K7OATxMUDaA5mAfKRb
kdZtsIHHTy+GkB6yOHKcdm5aCQ/6uR1AygChPcVwuf2izbTU8WqqGKau0rEpXf5K
Nih/r31+Oy1XmhStGDlVNFgn/cipFVx73HafiTZo+kGjIXCNvF77O3i/Xh79bN+o
FDTbXxvPeoa4sGajYx9WO9LIsbCN9nHIgnxhue65gEvQ5f437hSz8Ln5EGmAkB7a
RqLZVIEPPI1YGYmGPzbn9bcw/0q9JIihmjseB2gYzkX/ISBuqWh0eenFXy+mwctQ
yh6h9gmqQ8vLgbJySwRcxUL3c/FoQ4zSiOsWDvkIegZqQQfovohPvXsnYlSCuYyW
koWhFA6O6nsr0NAkqxUN1UGyfJPx46O2l+RNkcDMfGlL/ys82AtXT3A6U6s/fQdj
hJfFezVYoCrk2l97TWCmnyvAWwoj/UmNcnJ9wOvEhjBqXdkCDlCUImtTjM6sg6hI
ZiuVxWdh6YTfqLgnGZBDqHTnJE4nPPJfu9bw+ndicaed7zY7MFJI1o8TYAMtOyiQ
CUbDXButh36Og/R/Kj+MheOYnAYzSggI+GVVitZ5n12IQkIDcpD6HM7+36+zdgKf
GT86UXjzRSTVxrVzFXjICPtE7WlFk0S0jfNTXbYiFIaZ9FJquXIect0Da4Ge8mEw
Zm7oPtS/r+fdNtdbAqtcnLSF/+wuiDBtI1VjxuilFUPaS7Ww8pRpSsWB9e/PeUNk
zI27NWjY4Frq2HL9xu5O7cOh22rE4ZdqVD2m42/D+pFvlQne+1jMp/AKTjIA2IeP
ij0/VifebsMg3Z1e7hcwuJ6SITWV7mHz4xgYQzWNfjq75MquXvSSKWcl8yLCy/qU
5bEBemTv3IbNd19DezM9jaHqFWA/XNDTmO4SX4brIfpkeN1Y0zyfPYDCcYRxKC3K
1HtLcKIWVHxo3r334fR2dG0nIjvTLkqTQP5US8UDW5vcsAC2ZENEvniQvCHO6300
vq4CFvFVekUDDcXn7AU1jw4HKROKYnywHB4ffz53aSmHx/WtzSX9wyK1Mw7p7Ims
PidNLLfxig7DfLk/8I6D9UcZOISwhc0z56jd0vBX6CC7+NUBResDM6TtnLFJXA3S
haoEORFD1wFEJzsDfTAt5HDVpiYlGa+tcjnwuHu5ODe08cu0XJsa6DEdOJu0erJ1
lK4XDqLn4iEfqtkWAJDDlphC9A5ivA4BI62AeD5ZWfWD2kH5uxmr2VcMW8UhJN0R
iFcKigVaQqe4LoC+Z1p76cUWoa5AhEgaNqcIPAS7/cvUvc7a+rEDRdD8FdcTSH5U
Z4c/YBf+V0OGNRoiImJ1S7SYKmk4Z0it62UG0Ww5uDQVDxXWDvEn5AZgtj/ciVtp
L9/wM7eoY4qd9cmW2XVbejlM6a9XPcxnVCDENgdaTCKqf8KbuHJVGyKSRgPEI1Th
1SzCvDdUbfBLOLMP3kvgjMTuu3X31lZ1DkqyOFtfCALg3ENbV0Y4L1ky1lD+FQf7
rgGAPcJCOBB56CcBrJQstsmB9STQYADHx4v1WvvvTYTUmUT7XLg9SHnHRKY97osZ
+IBBtFCLay5nyvlBORKGyhmTmXBpSDrKc8ML4wrY59ALkgug5Ofwzy//rbIIqu4X
bGTUkcBngXGlvrY1YAcUOJ80IHPL/zx0UFTCjAO65MmUmchiwQuI7C7yXnaa+sry
0LQ8TDqkNv8fkyFTWZL0ujgr7XGnM/7c/R1yx50NSCLt7Gfe5eYSANVk5Rn4Kt1v
85fikTNTrPsVXJt46T9avzy2A1BAM7Pb1QlcV9qs9B/nc8kByRpWP9pOQuxgOtau
bDXTjcTQp8Me9C1KGmcFUs1RmO7BixSPwXYNd6D/yP0cfmf0agWKuWo1Edw9VaZp
H4RRcZ+WcixodQAwQarbbPpKCt1S5TULUgbb2eAm2CFc+rvhwf1DL9X1Iu6Kk9Gi
j0aH2Jp8q1AwZiBL0N9YmrpJrW/4zpbYAFHwCRk8pU1dbivV0Zfya5NBu/OMGxdP
dz8kKCF11wKRynlo2zExZvk2k8lxfTCbCY7QF+DmPJXJ1alnyTbVxdpWe9ZZdlk6
5ksm9HeqsJxBO9kP2peWtnNcO6BHZV/vYWfF2+HEwRXEeLu7lOalv7uBdmk2Wa+6
zqVrVsNeD1yDuwp/1PkeSEJ5PaLfq7pvBMZYK+fUr1VCm29GOC37RMTbRhdPN9d3
eqFuZ125OoVywBknsidbK32u0YQQnPyc8c68l9P3K0vDS8amMpvFr036zThrD/sQ
iDTlQ96Zym21ADw0IRK3qhFOwe1ede/jc9EiKBr4CjckkkNKnClda0Ho7G+L3f2A
nuaJ9GGxxryPklKCeuZmIpXh0QEasALZVKN6cIXYCU+4gqRTdvLbLMLHyZf2x4OM
ryWVVpOI5qJeZBdbFR2vwCwmmnij0zX9WaV9fJSCPaLecrZQIga1Xz6T4jReUiq0
D8leFhTE3LtS8rI93uDCp41Ko/kdd9EpyVQK3GXGfVmNB/UIex+ki7GhkkSCWTT9
diLChY1uPVwvwOLetw/xrmfsSzzzZ8aLTVv9xbMRuBEhvkGflQOlPywl6eHs2xWv
6YWC9lINw6Av8US4wi3z9nVkGk2HhhDHVEhj7mlokzZ4hlF2AcLzap2jJjzS9/Ao
fJKUBbk9UCQsaztZLVgDcBxUbV6cpLYdQmXlGednGy2UiIdxHXozJcLE9EhdcPxK
MR1MoQBC3CUGDglANj+Qq8Wm++byjXDD/oHojX0Q4+JSQC33aSdSf884DG+3/WsZ
TugV2xUCJPy7r1TqxIUK9ym7r+bLFaqW3NJeppIFpTjOSBrrLNHoZByNzDIG5WCV
Nq7X8/V2RXTcWAQ40Nb5KCvLDpLwxN1RnmEcT+Cz2ZujS8/8YYptUbF1YQghmTAJ
LpB/R42i9NrzXvDl7iApY+UpSyUIUP37IFg7FTiFlUfSl3JN+BP+8Fama5XQ/0Nd
P2F8vhQju989nYNlZjJYny7SP4C+7oukacklZYHfipLIEFRP/ddpDdSGW0JL0Dsh
q1cWseYif0yToY3Kg1Wuj3kyIhXACCSDQ4WT8jYPfG9urKx55XJlQH67zxR+oQUl
yBvvUV+sKifOaE/h3dNsF04bQwLR0yJbrriI7irmarHf/30VBwaSHxhrC7L7VBFe
iiuMxfGvGBvXXUIbLYmtSSnUnkXDpbsSlBcupul2Hl5UM0LQD0yOd5k0XAC6HZQK
1b43RbduhC0KQaLwcGX9PIpplDAtQMmqlSkBKfM3UA5lFtpITKU1FLPBIZ7ydfEY
yro/XhEIefU9CflR8uEU2MZlMjIK8FFc7iXPs2MhJbWa17dDTb+PcxmJYDqC5y0L
8N+s8uLzUWX+Iyqgbqk0xkDX1m6okGase3RjcmXoFvTP4ay/WGyrC/Ynrr4Fj/jR
0X04UJzqN6Xa/7XqyEoD/jSpbbQBiv5vjtood0/M90AiydjHC1MwJaSo3wmFOiBX
Q2AaN/FMkwCZKOJ3si5mwreUGWnLyJwFFx3iRKG3wop6vhm3d41pO9z0LoZwJlro
rZ0oqeARMLUrC/7yfiY5h+ZIZIAvVBgGgPNlDRr3KNKsAdk6pFKl+WwHIKVuMxR7
nvm6UuIg8EgxbFYFzv1i/chn2QAwpNelFwUJ+Syq7pQwjqc3ab2DHLHhF/j8mOrA
jf0U8BUVeOIieauw8/ouatLKNKtIQSV5x/lNt+P2qu5+Vkt9/9xZWypDVn6pBnpn
rrVkSWEjiQBNPm9zsufRzbER4cKO0Zcc8f8mweZ99hix3PhKStVUYcsDfWYQvMyW
qVudMAZYZL5DSRHVxOFqKCZQMMLMSw7PpomTI8AUHj0IOOGYpe2DoqfAQ7mxY3lD
HgkyGk2j3YgZDkF+32ZGdhkC7xZeNyOUmkd49oA5kpoWw7OdYVCGnqS7tq2bvqn7
QXa0qrfRus4Noaya3jPDhjysOKJfzjJXsn7x6OBcpoj3KdxR27vuG9r5R4nFSVPY
ibc8UMjCAEQ7jsQ3hFO33yXRkH8WPgghD/Z1Rbst/922qO3FNxWFK5iUDA4zaBL8
PHsvB/ccqZDHJoqRocSGKvjuFgluIeKEjTFyqnVCQZIaessELoavebsLEh0JWxPK
7hJgEX1UKc8eWMkkfAfd5gF1Wm2rkFAzt/Ziqx6t+jznx02kN2JCvFU4a75zLhff
8WT0xgPSWa9gpcxrBwQ5HAZC5P9RK5CUgoNc+sFDNFN8E1xrXoArVfTzXgOtF2wx
azUEBh8EuoNUdiSokC3LRAXRocpYg9KQJJ8nLgiqRrawjx205hmvlSgBRnCLjjBY
Ga8th/Vm+yO2qwbNQo17OIYQ3ti3J1/7yIBOc8bomfgl1m8MO8BryEYoKvmPwMj3
Yd2u8Hbrn3P6cyZ8IjMJmRfSboY/TZ3NmyftgaYGQjpejYwY9gK3ZZS7NlpAEP28
a3GIstMhQHExFDKVmVBSTvbS9Zg9lfT8pycSWIYDAFeujyxJBMNfdOH2FSlwkutS
DkE1jN4zSOumc1IIjDScfeFHWQewWjk3RI+c1i/vZMqZ3SrJ5Ap6LQj/2SG65zfz
7awYPuCa9N7av0SyFvSTzRa2k6b3B1yOpk3FRWnmShghJoHLKhhWrRizsaBhwu6S
M0Yc0zgztwG3jCSDhvqS3mONdVBO+/XKY/6A1t8pH5Klnc+JIyF98TVRV2aa20xl
Adkc3x8J1OooeppQWcT4ZgsJ4YySuxH0iYS4sy2XGH+/PsQqDh3rekbY6ZQEaIbT
7TZa/vo6SidXaFeKy0ZdvbMV9nWReMTW30aTcRvA5zWNgLNfO0N6jDQmQZgCpzXh
tHH8M8Us+lX2nfSdNbLrtveUr4TAqGaQcHRafFxD/Oc1l1Z18RbUi3QQRTYKHd1N
HXvZadYQ2Ykx+YT+vDIVmH6jDGtNtdNwiVfdZun7ckg/HabsYs/S09XBvr0g5tPe
+R8KT9rlVhjH14J85kPcqPfBZLzoYtaUdhMMh+eyXp1kX8CJZ49bnycMHR/UANoC
5589oGfseOPh3c37jAHi36mR/jdWWnnGett4Pt+vSw9RELx8O8QLYZ2d2HdqT2aL
jW67TDH1KGzTnEERkleOMMP9eiOvCHLM2ZN4/iCN763kY8HQy9eOaoqffKbUp3sG
kLiSk+2uCCVVFg8br6K/usTusFIAJI8Pk4GkAog9fdf1VJDArSbpJ6D83E7BSM9O
Qr9TuEgM5nnTSzN3JKm5v3GUgGurqjORU4U4N9Bwmt2wrC6QyruZcTlQjEhFiYsX
hwS7sdL2YIAv/SMP3oZ3KMxBhri95zsXa2N+OX8ybxW24AQM+EHomQ3rJ2w/n2YC
/q7GAE1LmpYU6kKRvRRPjpXrRcySOsfAhn1fBswPhDlLsvg9VbLEVD7bzZva9+G7
ABT8tu3Pp8BmHlNJug+Pq+PFao9itmlz9luYLnQrnv/ror+v5wjWfImsakkZepem
fzh/RftxqfAhK7sGCWQK6UpbV6X4JrAHgEHK09tCTsLdc2tDK012WKL1Q+shOlf7
fM/zxW9FxMQjBGDWF2LqLG22b7YhTuTn3CfpUaOyxCv3jN/cP+pp4vS2oh9oNCL/
1bSD3VVZFXut15mZABpc7YIDETr2hMA88jvinTAjiBuTeX8qNGSdoyw7MBbeIoxR
vFBInbUQnDCquhu0aC15+j7sAfJkFGPpf8m8GbsfhHlG1IdrIKGHyQpvIQHTaZy/
LxLNjeszVoG1hf7AYf/wxQM19w4DBJG2ZlTzGXrE3eOq04dOFWc7pfvfYczPrUq+
TcZeGCojcphu6MheJcvWRoB/4zx91I3K0XMrr69pQRiLmgrlVO4F2R1Rx1/M9/UT
3TdcZ4DQOSnDhWiNREMBgubovNz/qNvNeyOsl41LuTcDVri4GvWdaOvD9M1O4tX4
qeGW2NDGlbkBrZMt8VbvuPCXnAXrbLv/rh2dh2fQ8LXkbqkLZHj8e+MpSZl7FXGr
IeRLRBcP5mwMwu3ze5fqqxJ17eYVRBLARJO+bKsnB8h5SgljHaQtd8WkjTv5YAt2
Z0+NG42T2wIso7N0CDqC90a484zHPAlbGRQsnwwQMsbTh5ahrU+HX8Qb34wWahGz
fplY/YDj3sj2rcSFpNpg3nlwlrGoG4Mla0XCReS6KVpVEL5dDxOjYXvtAbbFyUAF
gSSid7QUqwLiHzXStTR3mCg0YoWiuWD7MPhTooMrgr1HT+gdUu2HP3zRuqU6K/pA
yUodKUPEsRjIV3a/NqCgx6x7VlZZW4YAKJ4f7lbzWyZXa/UwLxIuH96rwrxv06/k
qN+uHJOUITIDRm7W+g+8/Ipxyp8MXgySu+26w18VA6TvlhrYYNY/o8DOhyDTth+F
k7O7InZ6W9MjrbotpZBu5ZrEEXFTnLQzjzBB5Bh7dcEp+zK2xrX98J0N+s24Vs/W
zd0M4GQIz3/XXrIYMkNxw7rgVhU/hgQhiL0QsXEZjuybYAZWPGRe9+vO1e/YX+iS
alL0FGOaaxKYjDU1dKl3MATJFznlu3kTW7TcdBzwgHyRbkEmyfa+xWFdCyFb1xF7
ZfPbASNhSueq8BjT72MSWt21Be2pze6nqZFhrRbD0VSqpfxV/H5EUzPIMc7dEFQr
U0iFb1e8wRjhhCVSBU6i/qS7NU2XqXRcnIyWzyIneSFZeEqSKt6lixInkUQNRh54
SkaOSjUnoln7sDlJhlR4Pww5DiP+WImnENVEAiILI67GXeEcakuyA5Ezxz1yn/73
iypcTXnXUrlkaBMz/xy3THfS31/FICsIvRX20x0hwcgTGdYD0akzWBTPOYqmsutb
mcNSVgI3mZkFcgVQRTETMXoPs+ElG7quVEk8WzOdCobptG0FvgJdy6hyi58D1wrI
CXBO0Zus/8Sv7/HF1MPPiy3AXdziW4iISxXgqA+Zus03HLsLs1I/ygo5aU60Cu/G
R7R58YvsA3PesrpP8AYmVem1ceTQuH7qFRYaZo8zQgsgB4mdMg++2j3sp4x86yDm
YgbQ9g0UUvVmJYVPiQinopBLjXVRFtJILS40tF3I0Rn49uCO8aLbUxfx2xtgY5ho
mlYvaY1tHde7tzq48CGxnCgaZzWLje1SV5ceMQEdVBHBXcAUIjdtTOResGV4dh6r
Jz/3Glmo04tHKezlxE8dvoYwhtO/XbkemybSlcD/1wCLitb02it3HN5XHSkxxiAM
WPVqnJi8iNQWoclzoU1RMlF20RKTu7RgBG9ZPUbXFKBuBOm7QTSP21hZZPUYhSnF
FOgF1bQRqbUkZ1mjWrbgnJroPAdY+cocdZC1DOA1QQffBt5bYFOh0tFnLGc6SQQq
t56pPZq4Ex2hKzUrq5tOEgQ7ZeOXTUsi2CCIGPzTVTSGeRztYPCrZ15fQqP1GJ98
hNIC4FXmkFwly9bF5gZO6IRIXMG31TtsA497ecs4ayBL4plF35hm2vJJlvJF1tB4
bcz7hwgwwtz6l+Rc85vXhMZPupoRRE11mkuoRtuPtBTzA7tlDgwmlnPKFAOFkbcl
T/WM6Fv6ojFFzM6LE6g8sZD7tw5Oqx0evJQc9wano6rL9V+aYpfY4hlRqAxmcZPN
JK8Uvwmm8w1h/Ggc3n4cSpKHYHi2+xidjypRVAofvwQcW9Sr1/2VY7m9+oRfw6RH
oLQDyMLsRo/IFdfnUVybAEdQ3UtB7CXB2dfYEWj1fq6NTlkRl5CAOavLMBNcKc9v
XwnNxjPbf/vwEBE/Ox8CtrEMRhoMKNl/kOUr0JVEV0pzsmeA/qJ7XqunKlFhmsyn
0MJLmuceg1HioYF77XM4dg3KJOfHGNJwOEVFXslTFUYHoD3zE2MUD13mNLsk3Uh2
b0jwW7II2J6NPY0qdvdNXQiY3hq4v/9zThy2BtlmkzEsyujQr4MHasNKOg6zrDAo
i1jedRuuQxn/I7bQLw5/8yJLdtv9+cH55TWDXG1VzpjltgtK0dXpeye+p9hn+BDq
uydlkPZsT6f+9Q2jS6U6DHcJ/AB/ODyw3+I+/hX4CzviN8UodppGATfdVpbcfOOM
7WS5ov9iNwQvpD64v9L7V11NF12XlnF8s6tAMDZcwv4+dxbTR6kM8jpHqVOkc6XS
v9Re8nXA16nOlXrBi4vzVmeo1gdReR69JRGSbg3x+d2AS/5TI+3UuhyLvXDTO+pB
+B0WH36mAz7RXYcb0Qi37agb5S+LdQBHxbkTKWtquyZT9ADdkFr5we4ARQBx7YSt
BCTSa7B1OviWqgamE4J43ISiKJYSDBGuOEZR0eUi/6Osd795KAeQQXMzY9Zdp3q7
OjrFwNEWRCiVTy48t3S4Keq4tf/Mr87J1n7vhZZcAYFi8Xye4e9IsweTRjnx2/fa
T7VRj17t+m7xxCHgLVfoaOACt0opHdiih6957YsheMmHHlID47doiU4Cgvf/+u2y
xst6DSD8Rilv2Y6GrTB0zOFvQ/+jUFJJ/KeUB0fRhhZb+DeObp18hE3Dz/HGl8j7
/ceeqlMJ/lVXuo/kmme0gBmLzuQAqpHTzyrNU91oictMka6uroMJ5E1FYK9nGvmy
9UmtKBKdkPgrtKtv+OeOmCvB2jE3xy5P4e3fdnZHVRa7OuPZaow5J6OeyVnJv4Wo
fB+TmoKj4dXLnV91UyCCRl5rlhB/v+q79IP/7IfanIpODu9gJciKRksS3Flt+D4U
BcygkHS/k3LvYHJHaCsWdmazB7zMpcQuLn9PqOBNP+OGWNUAqJdkoa7ebHtBfQnM
iqqcMzfxnOnDvkrMVyj1vALhQKcOVz67Z1xYNlD5bTAQlahE5LmhbQ4rEiLyrfVx
XkxwSxfBg1ELzZ8VQ2dTNLd1QmxOAvL0CtHqR8nP34e/HwX/jhM5mcnmPb4+8Btc
74foApqtCx/VbBNiW1s/n9Tskz0/hiXOsSSb8Wyp/EuOS5c0RZ6gFHKTzfROiOGl
0tVdTooOJGvRExQmNE29PcxGwWIURIZFCbYVzmFSrf4B8mpJJdN+nQZ6Rfih7O9k
fhKwJ07idCLPDi7k1S8KkWV9r0QX7DiAckojlXOCFeA/KfAfP4pqxGXZCTmsFHxd
eFC8S4dI4ylPJp3PVp1KwAB7IMhu8ztwBS7HQ2gUb+kOKkeqZdr6CSIlrtiWHGGA
udeybe6UK0++MJItGFFSX2UlewFDc48Q/QadRU59lAHFmN+49J9CiZZIWOBiKvJl
Lj9mriEBKuXtIabsHaUZ1cnHMjfUwpGx3RLxdH5+/mjMaTgYF02ptD0Vrcmbgpwr
rluyuBCySdNb6sHJiBug8qwFzP/ZBMB5w8S2ppdG6WObsqtL5cAQsRj8BAp/uj+r
fSkQjLRf9ir6WycplYtmeLIhXEekOxBJRLrIWgLjEAoLK+4m3nGtpQs6zHltdeO9
l83tvXG+4ZPZVm4K0n6UytP4x7JJg1L5vrK/Mm29uKTPQsJOEip/feLsTEGXWwAA
QXFmRPdVR02sFV9dyGuAU28fcgdNfNg4cG/ZQ8lRnqteRKF++9eRUFUCLFspZQWp
ZqHn+k5ST1twbqFbQLG+1oj+aTtP5cf3ySGsSDA1Mdk5kAPyOk5DJRq97wYIAADx
VTev85rzoxKlKe1UiKni8FM/mwVEsoC5e0CR6BUhPjVAlBV5vAuwgRz8/1wHHTbq
m/LgerXtQCMBqYT0bRNj7aG7hKn0nbQMYAuPEX7zkdCDvLoMYe+JSUhfAe5HBy0H
qrZhusBnnC2jsYQ0kreI3MHKBC8OwI+TUiKuHMv70zr6QS1+H6P/rnHI92rrrIBE
sl4j0fnf+MxMdk671uPfyCN835QjTKFlb5r+P1lbgbGVBAFjjUmNTj3m9LxXK2lu
D0s9TiGbvj9dtUTZ9wTo8sGcJPUifHL/8+Nhqqce4YOwYhQwSQ5/T/ZZDDD8KREV
JUtpKsFCVxQV1mhi0g8UpTCuWOnlXGy7xhmMo1pmX0mAzJNsRWejaAIfFmo+58Wk
UusCC4w0Q4mNySPXOP/7DsmcgpqXMr2AD0/N/aBco+L0pFTMcGjUXLzEirfIbnZF
pd5c7EuoN/1ISBYpyoMMI7LBN2Z1oM5QF5/NGPBOKmnQdeLfnrKwR7qo/U1PsXYB
liIlS3grpZ7xOyKIdyU9xsucqnW7kM7OfLDygQCKyc24dYUtRwJW2w2jAOk+1S0i
BMtLws3gC2YZ/gP996mSsj/xvx6+FBvPW3POyT2k6RhnyyrHpgqMEVRB6cOS4fMI
LPNvIu+cTD6mWLI2lTsYcEed560H5R3mycJF4kyuVt+N+UQhNtp+txmNZWwVuGGP
VP0JuFD5AHArsxqbEJrh9bwYEOP6EWROA9oXPYlWnT/p0AKipwIofNnLMj+RGlyo
Sa11bczKGKX+k+8nOZ4EC1D1iVoyCcBOQh0cgkA9yQu7wvH55Z+QXlbJz800zRhU
ZxpYveWZEAWm12KUr5pvzHGRXcExAtNE3Mxf1ER5TmsFxrt4KXvA+aeuExBmdi0m
JG9tK9PF01U3hvIIC/r9ZTv9+SYNLWRZczKAZKPjr+mv0BrixjHzfMvZZyLOygfd
0fvR7bKDW4WHWIaWfxJmhsbP2OkZecrS/ly9BEksFD80t+rZSiKzdK1FQzt9f8fU
EtSxHi8ldlSmYKUdJM6GwJ+h5u6XmaWswINAUSEmA6qIH0ghCr9Eagz2AUCOvRZ3
uZTUaqK1p7XuTWNjr6Dpm4kra4kUWNw/Vs4eamXB9pdpdA/zublSFzMml9J07HJa
JPw7+gN5qHyc7GFDBFHw6yqmUQ9Alb+QEMiLYvYkyYXg5kcEV1Y6q0/K6wHkJIWI
pjPSSOTeiNfa1idpg2qLVr0gsdYjWBDDLe+ZjKAUaFC5KzrbKyfNw2ff6L1kQ4Fq
+sFUbSuLbWghXjGMvmAhaGUpKdfd3wd5HZn4lZsqATZc+gG57195e5yZ/b/3u5Oe
ZOwtqbHy2VxE6Wdey1Z1s0hXX+37gAj3TGGevULnOsNNy08qv0NRIIC2x+vfaRzP
Cf1rNafQt0j3wCZ3y8wuRGRtmBal6GoEVE3Sbp0uMtWqehNUoCMfOuxN0J5avAAX
iMqqBmWBMKu6B3K1UXYU2xqUaU8UCqHO68HWdL5o6uQ106HFLUa6725bdeMLVBW+
KadQHC8sV0+7oxhAk0w/EGXr/TaB0KkQvvUmklCkwaMc05I8hibAMtPAj0YOatL0
V4RGIiLz4HqPDkigAGSlMbuneaORmfVxuribtuNqhUfNzLibullvHXeFP+TBXw6f
ly9Y6T+mWhyWeI/u8tl1tqooJSeO3LZW5bKrIDwCikzJBA0Xt/Rwi/V4nY5hI9YH
DwstKEhUUkPTqTwmbtMZTqwEx9FtKWYVMpmmrlOYK6ZrZiUbLLur2jgsX5B7u+cx
vy6v5LMlw5pguEULK2UgQBnTQI/ypNT9Y93M4WQZVRYepU9scT/ILgzXbI1v4qos
eR910aYFOyAwhk4Ys/raHtGtljTUhOdy5L79KyR10R5PLZG6/dYRPjSL506AvkAj
iuzu6wG4TIp7rJEbTCXS/6Ir+AWfiVgM9OYo8WbuVA87SH0qwApaIt/yD7XKA01r
SQqHkcKVx5X9QZGj8OpvfYDWOk/rB4hpmMdarEbhyBjB3jiYOpyZua+tRL64CQCi
pHkzffwK+xvZfn4tQCK9o5Qc9EQGBIQCb3u2DDoVMtdXcG3HNyKbzhDCxQzssBC3
3co3KMTaWX+YN1jMrXyMzM+BbCTpCsXvkgR1FP/6NurgSTpcamnc3Y/wyVDfPgq7
Hnazb8e1TzQ78eV2JCAJ6c/Z/eVtuNV3Ne7OPqYy8KJHT8TfvAo+ZMr8Rg0XcyKH
/jaX/jczgYQB8EcxLiPL01oVmXzAn8MHj4gB+TUNs8dz2yojGjgsFrZR/cP/ZD3u
+4vDjtknzAEfnGXiiVDG4GXPKxNCnO6HCl5RQIDM6pNN7XPXR9+mmub9L/XWKNFY
xXOp32xRPyJDjA5GaD1UmZFqsHAa4CSj+byapho2Tsb4CEHz2Fj/0eshWUBdwOuB
e8zxLinT8lm0KXKv8FCACQcj1IHKpbCRl8F3j7Axw4cmwqMjOCYAJrOmwcT/EPnM
BKcLglxtfaABVlr7+UV1DNcQBdHcE7DGeDEKag8XUL+v5Umc93XZhD4y1OV4hFB5
OdGAPTVEIvkd4IOJlTrykntz71kE0w3fUr7XzcW6Ws+8/ABMSrzL9OzUIfGTFLNP
cefro24kS6JkbNX278/ojXRFJYRSximRkgPyAwXTTFQ+HSyQdsCjaAl34xTMDLte
KiXTnJxiHHwEJaQbKTFB/macDr6lhwgMnr8y5yyIHNjk3KWzFI31syDrvYtk/REe
ih6L6VZY/E9qS9wwsmCiDhSfObYg7ey0BeNeqCyc7LvKZSUlMufh/IL7j6prCpsy
MBA6D5N3omMF0NeGhJ6tG+RaGfHkmYA4gKG7xj8H2dypTRvTjJmfsNpKC1ugSgZa
GoTbsOpOQUFt5i8v0YpQ8qEFnSskmWTq1hCh0lmgn3hmTChxMxUMTA2pQu1ubvF9
GWEFL8zNfVwkFSyGquervxkpzIRv6b6LtxrokOqzSf38USZLLJyqdg5suaw4LSu5
ivfP0I2Ebk7VTzpsS7vYqhuX2SN4UzRDZR9K2qhqE5g5FVYoWwti8BJ1agdslRho
tPdXTwmC7KRJq9EOQOoVEsEqUgGwJDb7TCxBqmb0PhJW4h2xvuLp8vRo77F4TE5T
8x27h6S3KdcYZPvtlUmZEH+fvZg6AlfGalsL+6sNtfoT1w6ifn+OIhpK92tOOn2F
5xJcg3a1Ul/H1ONz9quliJttSpcOtV1EQYkSyrBMFec81Sdvf4+UyIvruFA8+Gv6
uQUYPxFixrG5E+bdIFSiL5kJ/SJrc2B3b4ak5JRBZjuwcRFE22nTfUnOJ1xXwNt6
UN3V6X+90NqdsZ1ewwZZOZayUgw6DspXVa066yCZSeIghmNyhojAvY6v47ldn8yA
39zX09HbFhke7jiwP2uX4s/WuMLurKiSH/ji/bBnlFEwyuDdlOC1ucO+lmDKF6ZU
o164OFoBOJqNQVqurBncblyywOgjDD72Q49HNzWJI12Ge1/Zv35dPey7Rsy7lkuP
WD/CVOx80Lhobtcx+AHzbeLANR/r+DmjxPC3ZN1/LpuDpcg+DIV8JJa0uUVDtToC
DZ/dUDriGPAniCNanZacBboTYhwKRk3kouy0GvpY9R7s6ipVHoSIMD4A51agawwU
yNHmyxs7O2IyoRjY3sz1fz59A+lTvUKYySLlNfUUv/mm+x4pvszLfjgvXQzbklg7
kUf+LtnzIX0tkH+Su3rayC8VEQiM/9oyiWitVgpBFJxPd6mcS1AcwfDpUE3DHt4u
roBq2cmslwNhLRhPGyfsn4OlAzturU+z5U9ku42f2wnaz0AtuQKLo70Apr9AADqo
fuaoUnoP9fPCxxwQO/Cux8Qqs56AV4Gw3ju7/h0ReP5kID9vswPyYRZJUja+pDu5
HUmDtjGakjN3nlIE+wzIq4nFR470oMiCQMda0vwGgRtCpsj3RqHt6H5MNIOUgfow
mohjjnfwEKp5MzMKS2lN3JkguppfvY91GwpuTxH9ADsKF3nB+PsR5bGTkjyExzt9
+UfNTyJj5pzvUacQgUvvFmIgQMnTmL97kQDRaTAKTRiar3TPGi7j375d9R9MHeSB
LJRjJHtD4Us8RXfLeE/yV5HEOELlOkScR1tqi4Dn9lU60f+MubA8eKW5LhAOvS0c
ctJAr2VA3T4N+YN1qizJlwIuxLBV9V3nKOiaMe/LMlnWhN+N/qryAUIwNB8IyP8Y
gc4FoTAHKMSHiPpNgIeW0hpZ0LuN188ONpd8U/Ud7/IbDOsqbDMMDzkF7SuP7mCr
aAAeVNT90aY8M76Pr+OjtcPgOVUgkrDem0e4SqH6our159ScLNmY797qW6CeuYO5
cfMWaZx0yfUEADvylISKzaK903ycavax3rbu2MLS0LIQk5fodH/EbokeltFEG0zM
zWd3RdteWCAQZp6jM0G8fLAZL1vi8tvmO42HXRz2+4CkmOI/OP9jpvKfRJrGgcJv
S7ikmb5rtK5fWF6T+8+T0CwRiLg5r1Flk5g8uWxhX4jNG/NZxQ8Wufi5qJhkIItu
q2Bx7DIG6pdM5nTzPfNgUe2dT2CL9AsUboAFesInFaXkLIuDSVLVWdKQyuwPsYa3
Wq/lRZ77FFhznQlIXMlmGV6v5SmKO9FChrsf309Ll/z1Lpxj+YhZq65rEcLZM5n+
EcdgqT1vFtdoLrPmPcny2Xfmdw65EuRtzIHWnXL+u0mBs7vwGyqJ6ZCaqpFK24pv
B2qzuyteR5DHgj3vohae8MKGmf2Y/aN++bqVkH4h4j4os3+6aEbvsyTSyBE1Dx73
GTP9P5YY3Y2muwKNzI1GlTwMpdvdXvjzFeIxOKSUvsCQgRzQnDxKqIC4knbbRCau
CxhpEXspOPEuXF1oaovkbRmcToWMSRCr/9cmlfrYA54T25N/4NL8fahT9Zg+udwT
VOoT4Be1M23EWRy1weeBpOVZf0jtwe96d/5ZNt7zok5k7HSjH8YCw/6rdLpj638d
NnGXPv1Ei3E4jYHwz79HBqxrqmgvEmFtXBQSKkwKsSggP2GI0Vx5Tg76SgPBu5rl
kh9dsVG/sHPasKu3xfTpMdnWYYI2iQyQbrkvHoNtlNKd64ln10XpypXKtkxUbxve
tZpOfD7iCZwU0YMccZP9Yj3vgOsOl4tZ1lIavpF+8L/gsXOaqetPb1ND93yGamXJ
a5Lfm9XhMftcNkHTJt4kqcu1n9GXkBgm/gZ1/GSqb/Oq4I3Or+yE9gcbnReYeBV9
7kT2y6lRMo7Jp5w9ZDcASRigEg75W87Sz15hBSOaZ4ufaNTmK1zPyhUHTlR/g0j8
oz3qdho+v4d2Deu3ZwAdIcwNS6F8fNyxVyvkKh8Ut5LdUuM2wDGxS5v1BUa5adjK
Uh3bxyvOiZ09lqycNCIHxnxXbYIXupCKjt4mRNklEBqg0UI7FR1X4LSSLl9x5B7v
CCHFoxrafTGLNXl+WGWnNShAPSHAkJQpxLNZYZgCWqkHRysTeudu3+SkxgAP8r8p
IfnHtoqvCWZzuRVo56vW2Cp2WBL542119LFSuXMoKaTNrV2RHov2fFXJ0nN9JV0J
ReaYIMBkTn+ZoWfxlJup0GXtcrfpq2aGIJ+z8bkFDdeysTAbA+O7gBjQyTlhKlrt
LrusZLYScFaKq/D8j524hc0HMmHjoDY2RxDuYnY7O5KGNPlcvxB9NDR0QlJZxSao
/soiWraDZ7C5m/A6Y3gzPO3kJmazJMFKrn2gN+wpowholo3cQR+tS3BpfHy0BFIN
OXFTSyJpDbr9XkjnfzbK7N9t6YVpK9ZWs4Olo0Og7/pnvsQt1cccxC6MWgQgz/ba
oxY3NB+gr/LQUaNwicOyZPw1r10K9s2XY5OxRUITWWY3waCq+q7xwZXkJIUVN0vL
BV6W8d5l0U0iEJxFPNw0DI4PMn5OvIIRxm0pt8PUogAQV6C3C4ExzaB3F4pqw806
SxgVB/FuxcXulM5ilFcHSuewh7hb6zrIC8EbRLrFp3ZoEc0j1eNhg7eOYi5AVPif
WTBOhsPuPqqx6vrP5naqvdLX/zsOKVhYfSGJfVamXvLQ83sNyRBe93ndqZmf2rAz
9t5CvI5zzxw+HAWhbjTCziJzfOvHzk85IGqUhwAd44vF8I+MsCSeDaoCYTd4WqW2
EUfWcITDLLc0EVvnjad7xwtGtH0vu/T9z0kjLt6Lu2p0v7eO++qnu5InogHmeeb+
bM1bVQEizLBn655KZDLvH9jcyYrqgaQsGv1kIj+CDi+bNv50t0tQwfS6lwk0ULMC
gRci/C+8Cxxp17FxE/imFtVjlDHBOBW9GNh9YRHkLteqXc7IhGmPztzp+TMCdk85
F3LZZfm0XMUqGZ85EdyvYm6CQhzzA3NorIWa82faPEb98Fvl1vJAwQ3QfnAXBfBR
eC7lfLosiMhNxttf0HbW/JCQKgBFwPxupRyt56iFl3C2QiAfn32OyXggefqOhN2W
RmP7aersTgV+mLcfUTN/y0BNucNqyLUaG4K84prN4bOu/B7uRQmmkT2le8byFlOE
H3KoplnLPEswKGB8Ly7IbhURSOEVq2aBaah7NiF6N+OYIrMZfEL6M9d+vazHqv8T
nuk2SNtNCUoOabN3eRNZimRLPJMcB3JSlA42psR0L+tq3CVseY1onO3TXTWIOZtK
NT3rsPokWBKT0vWPBsCcbQ2miyGJBeRIpMxdQf4dxIBkaCuHzquSI0Vf++3QcgnF
uha2f49YnvTZ4S3OdKmXTVxQfoYvmt/iU+Jl4YBFCt9/IclI3Juh1EKmDuCCP2JA
gtBGcSYp7NbjoDpYeWrVw3KkQXka/B/SY8TwAb6LBfHjlNYwiP71G6JW0nWma3/9
bGJd5cDVknDUUESkUROI7aYB28Cu8f5sISenKnmzB+0agl0ll3PxV7qbSnbY5Hch
9kDkULFOwQfRHhBZzEogjt+wUVpiGJQ3ENREMhBqe8l3sQYa8z4eGXay5H+eIMyk
54HfU0/OIss7MTO0QQuq/mPBT0+ssrZpQHdLNrovLrVr9rmdZNqwjVGiEWrZf4uP
UX4ah0s3QWpka4c8cqI6zgonN6oBGe13/MkJxLEj84qMIWqnMrSCv1RQdbpcysCc
CQBi+Gnp74xx1Hj98IfATXhS+WmFZPoG3eI4aWJq1dDN+wvRbo05x9ldnCiveGj2
n8L8W4WUB6ISsC9vRrmomlFzWecnAlSohhLqyTs8Zwv4lfR6qxaq+t+KUzVQ7ocg
hpKGar4zPpHFSLsLI4/seDzKpBDNLXhU8f54OHjfH9GDhndKcCi41JZifz3lEe9k
20KomRLgIvAcxJXsapAtRrSy93LYqL0kE3gS0wSeV189W6qfV/k9qoicxKCqymXI
r55etbj0eAk/O3EfLy8yGxhkedvzQQ4xs7TUlzQDBOf4KxXzr750goSm0R+o98ST
8UqohKYxEJego/JCgs82f73376UAr4tnMKgQlG5XCnBiFevLSqamhb9O04ZBz0v/
6B+ZJ6gzm/MdMARAMoiKABja5tLLg1f6TnGFGftJoroacJh8pzQOkGU2HwUPycIk
RBCjaaaY0acO3k84X3JsTqvfM9UtOteIy4ccOFbblIrHSCHtQ9/GYx+sFz2uQg32
Hj4gUxhoFvinKaGA5Q3RZl1Twxmhq7sxo2VnX+kO3YF8y1xNRXS2yF3Eff8AK7s3
aBsfL9P9UVOGhiEsA8y48AMyD/HwTI1vrR7OZxm5R9cpRRXsDm7VifdyDKNyIuDD
ED4JryhHFnHKe/KTxUP00HMzM72dKcxtsZge75H4BZWSa7AnNTr9wAerQZ89Gyfy
tBM0H9+/rHu3rIA1zVhJ3tN7JsaeOwswbazYOyVns3Q6nLVr40H8RiayJGpt7K5j
9CYp8IJuJA44I8X6k9ciwRk1wRBEK51ob0tEGLnnlQ1qPkEJQfz/Rl6WhE85LnC4
j3x95NzuiB5ySydkIxZO7kyQpH0RRQ8vr7fSti/8LiMTJO3nU7ZVtKcbEzU2noi4
DX2CvsItFFK55znBgYF7/bbY8yomiW/R92wJ9xyDRBKQ5rSSQwWOWKHUX+iAg98v
bpNNMMEh030SygO7AXXKqUe9z5m5ryKg4ehnqCIKvcHMGeDtZ6CcRFRgLeIPUWua
MOmyp2JIghpIdH72EIpe0G9SK7zm17vYodnQMzXDSDQuLxS8nbuww6G2z7CtBzTE
kJKwctx2SpdOwONFlsoJx7AyZs5dMkZbC0ZAPinQ3IRESziyswzeaUyeEOjTBZZy
wXa6OYdq2kZ5pYTcFfencY1ASVNP8+zSKxZz5drGHhi3RzvdPLzXFg+IrV7O4RqP
v75ayqjfgHqjkQvXQ055M3sXJegKHgwHShaXCQCBa3qCa9zQjRDwDdVVQIHMgtm3
BLp9AO7SpgfmhR488oAjDAub+5EfedjsBRLmrySSOWi8ebf/Y5riVEuVI3rGTq59
IH7kYPgmvzGkUoxwMJJ0C0jixiBzqvRldfpfLcjvqbiAEAp1/4Itp4PM1MGz//8D
xMO56c1sh4OJ+7vtnQiwHFttgNxAIkFcaRe40O/yH1PfmE1Fti0yJTZeWT0BeBzt
hq7yxmF7HyqAnx6vgAir7gLhYg/VGjH8twtUMeaTrCtHc1oWCbzMKyDf+Fqg4egm
9ty4X5ZicZCwYgv5Gsdj+hKNAq/UCIlhxM/C7IK5UUuRxkgTk0q/THfC75Q+HXnZ
+j5k0iBBHdwiMxN1Y/9lc7+EqiDMUuXSElYV8ctu5lvyFRw2wKDBtYzbuBkdlGzD
eDATY1jbTaj6hn8aoMtPDy3WtWPdsk6D42Lrg5ORDBNC4hY1Uqg6SwHgaJL6GDAq
dQ0/Q6G5HdD0wGtJ+cSlSReWDp7L/M53a0zqpgDacsIznKSglv5ML6Cl3w7sFkkw
iIuMrcmlJBDhXKTok+KdaJYyO2esxOMdeHUw7CT2tUVsdlmZeaJugn+EYo45H3Pp
Se0ErxcrMn/7FWvKiP+LvsJ2wlLB2WJEfJO8C1tQoEctceAcvDc84EywN1AtmEAZ
2B0n1XkbOxQRtxJCciU+Xcf/Yw3b9WztI6eUS21uFTzYRzzHIG5xo0523uX8B44y
pbLqkEaM8c2CWXlDRC10obZYbw2HkyDwfOC5JCiSsbf/LMtu8SOi3/64bw50IaPY
S9/PQo85YxN3xOhNhD6xkTNvYqV8YeWt2txlRKSm8z9XE+rYoV3GEBShdEbPER+c
QHxvXOeVrO+vNsWOd5XAhlz2JuC3bRFmaMZTiKLUAQ0YB36+YRN7MgFpobGDCUk9
79i+4JeuIVj1Z7epocw4niwj/8JIkT+xgATTASsO76v5QSyYeeTESDEjG4OfUi1U
S8FRdrP2LbEPhj1oi3QcgPue8DZYrHhvDz0dxHNWfHLYegEiMQyfyzVqdhVeYyKP
liT2sD+2j9RzXkqOQ7w+Gvv6nptSGPahGawj1xBkewiRfQBV3G78fW9plYL/otki
OicGBBAxmobhvfrSQXA6vrLiqFOcClssJfp7eogMwNlYKzwc9qOXUeJHpFGKEJJU
DFWqGsozzNs8UULF0pOZaB1ERc8iC6a8cYrrZv2eZtw0W5WBlDIfQ5u2W4NV7ybQ
QLSzvlPqHY/8EJY/6YnSDf242NAho78v7rBwMvLqcXWwhPoDSs1G3jBVedYOgL0m
ZmzmtSo1azDdiuz3hQDwNqyORvsiVqsMFeuF5J6+NASCnBv3fW4CYpOMEylyg8Wl
+w+AIrMJARdN5ydvQPaVLOd0HxcnvOukcnXw05aP+Fr7SSZRzlE5ywoAMGKL9OLs
qFYFpVKLOPutsPH4OpH0Z5M5DRqkmcp79YYL5OaYm4ffwlnueAmM5lOMx401Rq7s
P+0oSbScGRtxAsKoeFRX1Cbd9OKXXv3lMRs+VoI5i0z/PxRYqcIrpYXpoc/xr44U
DArUyPzP86sjYOro6RolSF73M2vqLd6RvfYbljn/RUiiA3Xu0/CX6rSmNsM68oPR
LSbnVn/y1/7x7Gc3wiHeakInQgj3t9E3yVnygNdcn7juTNXrOm1tV5ycWPiz64sM
F9oZ2CRH9o13GqspXdeItlOB/FD6m+jZi084CRB+8obPqhzkhhxkAo6mLXysbJBL
/Ufb4BbUFlbSpjOR6yjb+sulN4zzUsv55J6KBy37R8mrAICGqD6kcmhFtzS3zAUe
4kV+r+itergjDBFHNz9sia9e/74u2FTza98NWrI1BBcMXOE5MRKNdVMc5bMDkraP
LoMZQiIs4nTUOLNFUxpcXvVDrAtvpoXSG60To8SKZONbv71RJGGcVnqkwRmKw65f
6rir/DP0CYl8phqcK4/ODTmkBscHQz9JQw3H4Gu+DD1sAWD1ipU92g+zn+SaTB5e
8ZlHhAZkh6DzvZu0TM/BwU7EWSYscWKBxuT+Fbd/Mi+6uP2U6JAPmqup4NZIdxjv
fS/dPS8qc1FYF4I5QuvRntI361VLont4oHluAC1AnGq6FKWUk0z51MJrqRlOQ2iE
JV6htWeGp8Y5D0BSFuVN6yTFi0TKd6b2XXllEOaTdX7A1k4FlBGtdFiQllDwcjRl
sf/HbplXW5DKX2aCG6mERrF+FQyfkOWFccOzb+gsmXHc+1QZxdZGbRzOLzCS6pZT
hTTA3HtpMt4dAPcdwXjpysJv1S/IlsIAiYSJoPif/rBZ4RiQmMQn7rlv6SK/9WXq
n1IIFjSoATVBVpIGFGTSbJ3kIshnkoKYmpCB3/fF1fmryUwyfZlzqy0rIH+Up8dR
XbWnpVaydSY2n8hPH8WzIWPOZ3Z4dgkrGDxaRYGx85aNgyCQ8XiDyCbrBoe3E5RT
SdA13Q5afYc7r27ml63e6dz2V63oovzsmi9ahkMQaRhLrze6pVoaGM4jagXQhvpE
kftpnog9IOG2YOE9XK1XoDSvjAnpAAgcFBnfReLWJAaUm8v80MwL57jaYt848tK9
KFxXljNo2z/olnaP54zl4M56md/0mo2vu8XvS78xlne+63+x1N0V0u51g4XRsvNB
cDtotFX4GNSXzfpCvwIgGkqM3A5kjZmjnAmTCTY+In7iSvyuryL9Ubafv2wVxqqG
LI+5u6KIGoGIgfgeGmJcMJeBWqBuYmRFvOUpwhwgvceYG2DfEsmTNP+aUGZO0T2G
BmPwAO7tSoEwTkjUdVzg1UFLtA2atO/x3MuD1HCDx834S5FPm00aqTKmz1HU/eoD
b5pIQcOZab1QapCQM56GG2dA8jXUrojV1e2uvs2BjJVpbjjVVbvwFEx8p7q0w4Z0
Kl5Ki3jTfaD4wImVr2WEo1LTaF12A7xL9ZpIVUKQm1IZ5xhsZ3J4nD3Wziblozs5
9gUNarQqskEJ1HWibK68l+nPb2p0LQjElpVVZXov0e0MU6UjeegId1qQoLxyadZU
dv2nmmN2P6s7q0S0Zo4VEX35ZgMr/JQ7KxS+Ch/EXyVEepqOkY3kCZKr6tcifcer
n0C2DRso3s2tVxCEAuc/hk4413/U4vsZqxLDPkXAoLQjPVduBw67uEroG0tX8CrI
TELqTNwu03cLU2VAa+mcs7I0M1s1KAHoOopZrEmjTuHHbmlPs3jdVOJbz0E1OLoM
5nQ84yrZeIYvJuAspUnlWhllQb9CLBAIGIwmtXVL2IQGoRunYqF33MboO81K5HU9
uJazm6CLcXbq128w6ot7OASDWGk5d4TYuCPO+p7JBjfuVufa8kHDucaRdhLdoCVp
mZum4//rElvTuXNglhrLoLv95pP8U3meDohrq59A+bw9eoznl29I8w1bJUv45jgU
5kiowg93V9r/TZLYjIJ2cs8KMpp/ayDrVA38A4RGttA14BYjLVE01Ny/AaQx45+u
TM0ypJOIVh+cDNMlsEcnvC2wZcCuWX6bi7c5JZ4pT9rKCdDKpV4x0RqTBbwOB1ej
3XZ+XZrRMJ9gP2rgnIWmF8YUP2XHczDOr2jFmltthYM8sZ3S+grEaDBp9QYatdkQ
jPXcrXgOoIcoI/DYGINHq1ehgr8r6VRawkKSxu1PNso0bdjNLk3T+qcPERdRdNYp
4SjgOdQBUnN9aeg0Kk6L+qdNf5PU2CpXNv0Ae8fSEqHWq7uV72qJ4n7VFp+C01+m
gjozFPGWM1W94/+lZnVVPxqS6w9U0focW/Q0Yd2AewgWypPUeyqPxd37OEMCJop0
lbaOWKEF6RxABgG57jeufzFzOuCGtZr2TcW9E0Ercu578FUO+0nvDq4l/X4jtZWB
Or/zR8ifENXKjR6VqghrIJzBuYeDXmN92x3aRcnd7tFrCPSdfMdVBkIEI8QmtcL/
Lf5dsBmjyJIAnIW8LCJoJv0UisX3ZjJD4JJjTRUNgzmUAykf6j/76cXJBlgY/csh
ZZHci+zfMVCy+7kEKJMuNPFFVPRW0Hxz1oysZ+veOAnsDybdB7BGJlEIrrFP/6NL
su3KBnrqg31d+23yTca/rLmQ3TrVBn/BLNnTmQ0qInKZeNMRBmxbOkLjt+JKj2AA
TRF1wHtapT11+nsCcx7wxtCwQMMqWvDfl6MdkS9QJN5PGFFM6ZjZbLK9heZx82Ac
QOqSbvy2K75MrzFEtBG+Ex9hMxI4wvhmD25Ny6Ji/kjJ9dn96oWxbDNhapPiJmiE
aZw1f9qpNqwubmqtDf6rKcD8g4W4q1KgLyctVH4eKAWDY4LrQKk3iaIYsZqxUSj5
AxlFroN+6Lc0QiSMf0gebngv0YNnwD+yKK3bVZwBF171ZX58hqcyxUYwRGgZ+wyE
L0D5E9Jq+7axjz1bqEnzL5WI8ANQ+kb1PUqFQO3om/7NmLbWZn/EqY1umAdhIt8Y
fqb0pCb0ZjSC37klSmjgQgizpcKQyGhj7DT9KAyxPDGXBnug+piiToGqrD/ia9X3
FDxGcH2SVsnZHswabcqodwU6Wwkc6xaUR2nTdd1kSiKFAE/qTtES5Wx8HdYzr5ho
0VcJfCsbXus5E2xASc7ZROhyPf7VyB5cUvsp7w+a8SbQjoL7cZu+e3UCmMAApjkC
EiDZVSPmMsNGFz7qwS4fpMLt7xSTJV6iCnPDKdGFoFHGugshm75AvzgWojs7I3ob
2jik8AVpIC6KCN2BkZdvE18pd64d8k7vaNUqwf0ftTy1H8RDjz7h3HzzGaWmy9Gs
mPr1WZXKeGBdFTpHff0ROMchjkXSX0/hPAGDf74I9J00yEHTIm0A4PwYVmIsb+Sw
bjpPkWuWJ9+asxg06P1GdL7BZanPDLq+R2O21gZnaWLwedme4rV6R9tHCjxw/7p/
hVyRAV3nyDEL+ljHjC7bzWo7qlyZw433C7UWz6O/eNJBBPYM/1b0jJBVd1UtGXlr
J9dlVEvn6PReUghiqoQVEfN9NEyzzmhCSkfPamFXO0AWju5rRNZxGCkhwQV2OueN
Q5Q+755HuyrDHTgHdWuFg8TBxK90Ke7LykKdgfKGgNFuG7OtQMdJaQXruLKQ0jUA
0oggOkNTv2dnSoNjF0R1JXBhV4oL+eKMWgnNB/eep7SEVV4MlW2+xsqstb0xVXll
rkP/Ul3ZxbxhrIfNBZvlQgo0CAS1Ta1q1YYKEFFpCGN40ujdyNiUKb7BVuguAEk+
IvnTxwp3VkKNAoBVHqZgaDC243CaUO5a+NsPqww0b+rVtZztcr+8ACI425Prh3c8
v7YV+/8UuzohFN+Etc+LT4ytKk0t8H5g7GMtWlHLy89GTOoqhCH7i/l4rVNvOlQE
ga7MkcJT+PoBvEYnjHX7hU2Ehdsy5oPkGMuuOrAcFvd/lZuG0Gx+lzO7iYhiX/2o
7/I8qDw5U9tm6Iapu5yfIw0zMNRIYKSIW1+dhTlP7mDz8M1pYkMtXHfcRyNKPs6S
5dsQA8GPlRgJsc+BoYJReAcT0bzlXOnbRT8HqwD3C36N/N3FXHcoDAvv8rw6IGvr
nB+V+LqhYHOL9clkfmHGy23MuRZBR4/wTfvcRfbnjpDps3dTOIKBaO3HLSiZyxSf
L324PYNwdFCUwse4Xv9emry0aUMaRRhdS0IGf7tzIz2uVHLgqz4PdundxQq5j4Ol
yXrZ8a+CiJlQWTov6GnLoa6hO8Ns0krj1Zl3PBI2QzRyHS0BprX65h5heR25O0rK
D7aKShNq86IjjA2lruPCs3+MO24fQTKI6XtfMMd5agBXNVgUeBWw7SLhgzgNI9RO
0TPw6eigwg1YNMAj9Q1fyW6DRNpdc5g+YOijVEHX29ITZ2GIE9NJhoupfeTL1D1D
14n5eAqC58Z8SzB9wKX0qKASHwbO2UGbXkKeD5lYHuXOJX7s8+wWCy7lru7/uVMr
uslemjS67JB9bdKDIdHp0hBb2vUesdMbVATYJXVE79mL0k6jCMQMHj6hSBPqudU5
VOcJfycyvr/TU0ff9z7YMiwB+NThn4V9tpP501PlS7EgouDdPn+Xk0rrbLu5Y52r
gwzPIIwa0AaoNzTesN7q4CUHriZWsnKIUHpexkOQ1Z1LBM0FilV+Cz48RtyvAa+M
tMAKQpDYlmRDNv0qCHCiwOJTSpAoCSBmc+LpsVkd+mpJIPxmldjLxACOR1PAUGKC
4WRdwar77KO7ROwJTHtpgDSy4DfqPmaAkqJYpXTXyXnOEqIHi1xAP5c0wIp6ITst
QCqWoPnGOCvGHHUqAhQk/P1CdfH5eUy+VPrQ2JAc+BBW6hjVADVEbK8pAUozt+oH
E07p9SCPofKp48gmivY9dvgEUW9hg1KStUAbbTyJ1twB+FMk0aYCInrTztogEnR6
AKzs2fX7B5bwzdLT8bEZhbkKLw6mV4iJn+lsb9bfZ2ibTVii73vDcM/0CrKkdV6h
WLixhMFsqObPnpPDZC5ZKQpRyTlVCRSeY9xtPdaqfD8a8S8nBBsXsBYysP+3rGut
18cGTj+oFxzOgLBbNdnIIbljbouMRfzfpjHd36j5NvaZELBA63TQvcSCMbtFVfHr
bFNGfbi/bqfu9Vo6g1h+hXkh+eaMZDeKknQV0AQcMuS7gi+JttdmOQMhBKvyUir2
l18FdE9gHMMAFYfNIEPtQyjgjbix81AsDP1hTNIO8q8KW2fKhQt0m8Sda4D5qE+5
eqc1K60KssTc7klerbfSvAUptNswNSpLwS/k9bTgUYSeFufALcmM7xIZlQX82zDp
TIgRQuHPYu9TJYCAX9wL65vlaJCPwQns+mNawrnKLaDp/ovEHwzfkPoKarpQkPBE
qRs3fZaQ8mgMwGFp9evOb++jzdzU/LuMCO1qGPFGS/vUyrA1Sl1+ehy7MaAG9h1j
vDOUEuGSaf/cM8XRfEdiJr0uVmskBIC8oJDLFozaWI6JavVHi6ui5dbziCcYRVUl
wSBQVW+3eFr+VdXS5N4q7w5Zcda3+CWKhROU3oCatKlLzMjNNoOzYS8ZHr1Rbjxr
hBETDHUZ3PGPoIiqU2trrFI0D08kZwJ4m7eJm7N7nvTBMHj1lG6wb/Xap33G3sDU
aYRyJwjAuRRipBWsQ2qp1WAZ6Uk8moCxmNpV/PwL+ZfWXIwzGjRDGwwXukbXfGQ+
04PKKi1jdReY0sRj2F046kY5/iuqX37WjFhTBCWAW3tyz5+esLQhtEWJxvd5idz3
L/gwwwe8GyXWbvt8IxcBmSVRwR3OyXColpyzndidRpi99bjGuIKm83+5XeaCtHUu
3Jq77S9gwoH96sEpFSvVf4cbY2yJ4BPmBNBqG1lseAXFQ0lHGlkyvcJQAd7jTWEY
Lyp1WUCn/EPAb1Civ136sNSC7GLnzPlDwvb3/DEQI8q6pVIHXa82LIoViiNZSfMX
0qkPT0ZwBXUSCVv5/r4LgXZmuZi8cx7pa46GAY5EvLJRezEDBKKTQ32BEe8ugiam
SrFaAT6TH1jhvmNjuBt8/CN73P1Ktt4PIijrK9GP9cJvXO3G1u2bswj+CmtH8+zx
wDi8voNBfnQ0AjAL6HXHRgLgXIGO8lWHKN4U35TuaFcKBRi5h2I9ZxfdvepHBEVW
SFR1yToFln3VVe27jDSvVeIFgTdrXlpN6Wtyrh2ogR3ayqzo+0w4/E7gObCc/0HZ
AUVNSslZD2ZJwXyZaZe5bXm/Yo4UhM66a/uOXXNU2VnFMTjHi16LCawemfEL8mgY
hUS+RtJmbpZq3ArmDy+lypGQLL4ysrPdKFDcs/2PiPyvkWs5sgeMkEA/rjc+cc6c
+Szuj1sYrvdisPDTF3rcg8SHLyVXxJri2pbhzM77MsiUvkSDYqFiqO+qpk/i+3wm
evzE+mm/Cz14gt06IEVRLhWPfnoHaQrXHdndW5CNIm8xMizOpLSKXu8UP5GNZZIW
PpMsLEJ2q5gpeCT4WbjwF8DVtogjUprsKZ0jMSqbGc8GWZtabnIO+7aC1L3xkM2z
5vALLjzORBnUB/6P4WTfYmQer5qkc+ZWZYdXOe1m6DjETZNnhkpM4aU88bF2yBzG
3INLjGTWzTCt4ryWmkvPSZiWop/CKcnskTf0UbrM4muHpbvrCbmDqaDD5nXEipWJ
l3qsIjKpgBczsKA6hI2VHy5lzbdGqXOhTfSQ7h8f0MLPiNFr5DAaEKDf5CMe/XKL
DhqZn682G+E5u4r8lo2esuzwZCIfXTHZ+/YV4D66xmmcrRMTa/pFY6ZHwf6kk89F
cULBEPCvTlsysYsikF+o1Pn79u23Rz6EGSgbw1lyU4AFV3t9Uhgkv6VaJ0IoV3WI
vbMTJzxtlGAM7sqBjausnv4wzm/Qeuxu/maE47JpFXP9LDZ+eE5ERU5HPNY0vyGY
lVnQCUUBaBzpHE749Rf9MIaZjjg7wiYb13I/lO8T82oNl2XzItVPSIMZyTwK3Y3f
1YI3sudEuzi/8S3mGFocpeEvCwB6c0odHwhalaG/P9XU6nm/PST23gO0feUIJ3kk
vkSTJLTQJ/nxuzegG/iFYZV22sPxwT2Y9IoggPJ0C5bjdpPQXkLwC8uojh5bIuUb
4HNmeDCZp1XfM3LrnhLn0T527+mVarZ3KM7ukGJLlMLYI0dbLzVRLBL9spd0lqH2
6M97vYldNHCoxeurOvJ2nHag9R1HuAO4edMeHSghQCqaA5Je2yE9MPHEzYpbvSG/
xhYeHlDJTIWy2+xElSorQ9v6jxEvdPPuIhPGekhmfX8uY7qH9//a51hVUMgl14cS
rqKIM3LbSuNNi2sXSafiUiwxFx8qNAWXL93Cxb2nIiU6G7AoIe7EN2k/sZRGbln5
4tMlSDNIt2R7QxVBY3CIdZIsU0+TVFqb4ufkcslDTHMfQ31a5NTHp1lVRi5ILSQQ
Ff1CH69w1/ao+Ia/rmPo5vKe5lcLLuL51jeIhdmhsCyDVMUcKdlraPjqzh8a9Gq7
OzWs5+O0vn1ZATiVIWgBPURAfXNgP88LfkfbbqS6Z7Extvuc8X8ntbF4s+PobxLi
IdXTRsWEEFh745b2/seVwsu6VYQ1igkvnpZblexK0Q1o9qCVnE/2zCgdB5MVwrpE
VU37eK6pM539b1x0UuWRJlR4Wg50sm3QYWzQQzCh4udqYarFJE+ritZnboI8N4WM
gTmNF2KOblvU+oMRlhBwOIABY/94q4FbWBGj5f6tFFceZ2AgrhFWl6xj2gOvJ2IW
/1SiEuJDvcJT0EwpVXrJTEfN0OBmIoIxDarjdK2jDnkg7Y2qcWkxXCSjejlR4gt1
jgfePBR0LlX2PhkNxd1XfnN77XKOQtUuaAcxjc57fzzgeywTsszyrGfk6pbIgWJi
hi3Bo88SjHy8fCM2Y6LdJbrpjjaTaQB00s/bdr4IT50M5aG6/jVkTMLxUw9z1vTk
oiDCbKNxlt054MrzxcjPq5pGML75irRZieQLu5aveW+lEfdlLiDg/7+SHw1pU9T+
IDro0sNX9jxnRDIToOue6aLNp2WR4Q0r0jwAHzuFlukygI6JvuJD/8qbl2FetjNz
XnSAW8y/OnIkgx9zYC7ayAPIv8jMlSSVGzplQCq2LYt6EHW0SPdaPa3v3CVpfVmL
gmR9nEfYUv1rU2ebPT2du8SU8zTNImK6TcuXRU9jQKYP15CCYSEtIXZUoZDl9KAC
xN564XRYjuhRJivyM8DEZRX0e1ykefexkLvoP0KcfFbiv8FdOabUvLRd5fKNosTz
ut9+bXKMOU9k3epf8jHcrDAcBNp1WEEuVUm5hhnOjYAC5TNOxO72/LSUJ9RS21F+
mw2MFUB0B2MFeaIsumS2P6HMhG7YSLjRVcLWVKyu8mDkfGBfVdbNL1DYaafWcDdn
fcQc7fkJniEmARRWLFEzRgbBLQkfwYxdeMIyLxnoQoFilFA+HeTl6LT4uytBXFr2
PJyqofPOnblIxGwNGnrE9dolNqmTwtkJfpklqPcZqiJ14ep7t3MVhru7Pr7m+YF9
d/2thfxufRqp1GJ1c8I/5nBCXmaMUAHVRUfRTXYiwe8/i2Bo5xzji5x26jMCrN0h
AKBt+K2I4ZtjWJS6UTCnorMvKfUddNjiwnim/NVAr7l9R43oqPhhYe2MlrXfgPTy
Lq/QCqz1bV8O2pmnUqcgxq2jZhKw80cOc9NqjibDqFdhAnZSnue2VRLe3Mho5rxs
3UpHs0D1LqJsPUTziIMbRpNufTPNZ5NTyS5kyoUEcuXt1+IarLJB5On5hH7YlHlg
fC0IT4pnCQ5AJGtowTwlNd8Zso9JSh+j8ux774tpKGFEfAfIUiO1MJMOjOthUdgp
sezLd+lXbVaTi6i3yg10E/WlsFc/FCFp5bnd6Scni0/ezYPNwpRLwAyhzuSa7LvJ
1n/fcg6hSrFc9AcTjw/CiT3X5dDWiX4YuM2MwIFWeK+L1e85esgOmhFclEwkobcU
aWpjHT+r73Si+hVSO1cSF2zIkhWqA7tv67MG6fA6dC8T3Jd48TiGF7NvMrGdbg8f
x7fb2EjHSF8SNE/tM1GXty7uDZWDaLMIueK7JiLxN8smxksLnhi0Baaaz0X+aPbU
3nZoWrdPLW9/c7jyCeVJjuM4kU3OP+YdsjNLGZSNlgUlj8Dr3SCnI0IytZiWGdp3
XhhNp3UomtYBmzwV0xLOhIp7Z9ZBmKx1UJVw+36cf9jsW4Rqxsf1sPzKfdJgn3LB
n2mQmVCMOpGzEdAKo3QNr7zbBvTr0hAkxAm9YMsXbJVLCKUK+c7CEc5AiX4M3R5U
hEKkUa8bi5540B2xqoEK8eTKbMU2s3g45w1kYCNMQ1yFu8tFjVl3rG7njo50VCzA
Co02T2UcVGKaYF8DI1vZo1Roiq1QDv4qBj4z42XLQGWD6eLYgJbPLv4CE/gxjIrC
/hPLnQ6hxDm0C3mnCwR5IeTdkM9Dm3ARgukHetkXXrNpR9vFCNpyteJF0msn5y0k
5dGUsAgSJD6UQRFVFgDewsXBeIfjkAo4cCHmwJwwED1SrYX/TkTYqCSKq33WNu+g
x0ECvmn2XzMxKp9To7gpHKtvy2cv6P9NPrzmq0g/CFxaO820lLY9izwTqLzxoEPz
M7OqUlNCCQ8z7Ia3jN15PlmxT8qEUt5PebbVO6demv6JIUGlIw9TTcQHbmmwcyer
qzzEpOrSMMyrYpIU/QTUQobXyCocB8k8O7pwNt7TygCu8nUYIu7H+kJVDieFOfiO
kMkaDIp1VfGeud5mVuq3xG7AGuO9BltZ1+vxg0Y8SZANf/I/mWPeWWE9pUtheLZM
P6gD7RMRTqIh6lnhh6Rkc1k88vNakjA1llMLmsCt06ahv8EBszunajgPG4WLLBx/
6uhA36X2Dx0tnPZwbGEliGPARCY4IBuhwLD+iVBmpkMzwBvBE5XOW95/HbZJ03dg
sBNU68sYh66JGimmPT0FYoRo3ElLqX2IzuuBE4fw3q/8qEJnchIjnZczNGMct4BH
7SvlyCU5lXXAWDggaJScj3nxcIXOsCesvDHH+TJobEXzVykK43j4LUPjcuU3Qx5d
XINMnLxlTxTGYh3Lo0zd3c+pOKoWbq7K4Vt5AIE2SkyKN0oTwTBaw8HlGnqnwM9F
B5311d8EGSWYHs7I9yJ9d05bpbKDg0Vb+j6gA+O5RaAqCvSG8RZMBm3LKV0jZPQc
WLg9Vl20KF9ipC1pFJOvaI5l/n4dlLuLy2ruRz0JasbMpwCUQPcN52qki0b5T3cW
4/Rg7gF86C9yZeB333QuLs4VYvVmuMdmfpkXrGQneSa33bXk+r4nP7dRgT9q3Nvf
mHNkO3//GHwApeovqNrNv+SI2ip5uwcolzFobEXovC9vNn+IINbNOlMLPry4FDpU
d9so49MtPB8izo3oHyrV28ZMkysf7q4ayHs5mxPnoKIO3vFpFcCHalLe03mNxXZj
utO9QWDIUlyYBBvZ9Sktrjm2g4jN5XZ7LBqocYaG5SsEVPrz5S6tCtdCWZQdBjzh
/+P8tkW5717tcO2BAvjeYJyV74tcm0o2P/eRiE6Fg75//eK680GJduAuumVk9Hkb
Q1qDSojSQ+OvvQlO9N4elCuTpg+/6FGSTuhMRTYgJFDGW9hfe0XRMF7I5hUabisg
P4aNBPVZ74w87daAebke0fRXf+U1uL1+D5eWg8tQANVlTTt1t+NQxU14UuZIt4wG
2DTB19wQcHsEHgtvkORVNcaIZXDKwNSDKNze6qfkEBedIXB0SZE4UmwjVkz0riZD
43UlQGgwCijI0vYjdh8Nd8FFIBaLq7yoz2Z+nZ2EArcPaG3xtutoLuOZpWI0C38e
wsnwiyMNg6YnlBgaVsx3rZi8rAqjyZVkcDDbkRdjF3cC6Z00DSv+UFr1xK1G2sn/
/7NN6WhQqDj8TPJkJHsbH9SvUd1oD8ym2nxNDA5UvDaJlhsEA3il/JaUu8MfEtV4
bQnc439YoTVzuYNE/heaYmSC9/GRd7+ETFZqt1VLIk0YTcT2skUxb0rOqyd0IpBC
9vn1c+m6WFIZMKclTBZe+whlLe3nm9QMDeog9R14VFMrYJZqqlZoh65pneO89/ST
fOcLu9Vd/uFXF9ITQUSx2uK8NqPBZQcDYvIOAH71iKdv2r2y7erjJ63zGboQJvM2
iwC96GblWeZrY4SknbSsIWyLdnRAkdiERS9ibU7lKCCdoGd6j8HL2HKfGN5EL+WP
gexrtH6U5yamKwNRf07ctJcAZKjNjjd49kgXCLQjMGhZPOOQYBIZuDgxNInO081k
dp52F+6ISPB2EimuvPkZsz13pY08TYo0Z5KY9GXQVTfZNFW2mgCb9HiZE7XuKqy0
Mb2UNG4uOhhKQ1mHgPpZqkDH/Co7K62yXsyNJa0jRLudHVWjsk9qW2Na0bitur7u
+Jp8//sd9K/ghMjqIJTES7+nO6FDuyobWh95+L8OV6R3hMLG7yQMYMPd4hLVGs++
OzmPZ7MR0TYQyN+OmqhWPSJfhj9ssSJMoRYkFLVqUZiFvZUTC0AUwojW0DL4lg4Y
94d6o9essVbNo6393oCMT9r3Rzy81CxKc+jdOJrtqPsvyEQwB+OVg8LCD3Z+JnDD
wdAL6K5h2PtzdjNV9F3rN1BPME1ye0qeR/Wh13qfntIYT1UB0/8MvUQrVbE6BOBW
1W1U0X1IX5xjenssMTMTQqQPOfH0ahDWLL388bHpUCXkW3t8Hg5RI93jvRuzqNKl
v6WBAGtBLahNu2m+HPQogHk1Rnoea9iANN+ZPgJhJeGCtL+vjvzSr3vk+F67ON01
arJzFalKLhazhcTKCgQr+AXhaHC5LXJuBGVQZ1VwSSeIgW+63/6G13lVIPFXvqEa
HG/K4Huj1N87lXCDmEQMk9fWf9PwojrsWCBS+vgDb3/sE3WvE3Kd3fAWOuMY/xe1
vdwvUV5uzGb+Uh+gVRllQQFkS7pUD70g3MAFdLiW81ewmR4C1c9KADn6UiQLRLZB
30HtT7UnuKC4s8EJlO15Ai1PppBq30IqtDeMhjDefZ3HuWHLezG2/ogd6yKzxXpb
1dckzVobcsVF+SzBY6A8xdGCKDkBGQC+O8VDV5017fEh6bOnzrjwUSgMhn357OKv
4Etk9K9I5+/A9l+yxXmayE6+/D4eu1cQre6Fm6Y8+dPm8XZGyxukIsykED/DxGO8
SA2Fxitc8v5IwhJK6uPfU/C1Fhv+7NqYME3vueoiu3LFjWSac/MmtDj4N0+uWPBy
qWlTRaIh6I+Y3WRfLdm/Wd2d3vMICLfxv1iqV5PlIbLUIi+V4Wu4loMgOtv76RkB
EXcy9tjjCywhgUoklFxAAke8IJvm4LsYzWOtUkSyhX4R/KrIOgBlerrGvOHLVFQL
w/hFZs7QLAc96XbnMqpu2D96f+A2d+/h3FvteQJf4fS2+LGH8o80fR8/HdhsptLz
7J0vCEj1km4XtEP7sQG4r3FNIu7jO5aFf7N6g/ldN0AomHOF674lQxgDLJhwNECe
Yc4Go1uMHsK1dTbl2d2egSv+QsURyxJ0STArZTvrsYagqDPQaTXk1MCr9gfV++0q
KsgxywWKrQYcK/yDismD7WLp5rOh6lTtKtNAAorx32vG81/eIEZMXgMQM/p4nyUu
QEIaXMQj/+uhc+I7fujDqgwXg6wExQbS/We0Q0q8QpqL6zgsUIwsIwv7JD6yZ375
B0VKJR/JOSRBmBbwG+CaUvExwIaOiRL0MG2dYcdcvB28nP/sC1nHl1v0wCvgiJoB
B23vnWYWpHiO3oWI480fz8CmWZITTFohvSjkq76dMfqtv9v02St3tIm2xP0UZjVj
xEyI1EW3jtuIZufqbHsAkCDpSRzEAjOB0kh8ggrjqnj44Hz6rrt2uP3V2hA6EdWv
HeFlyoHByw2IILBcPlhSSa25tlxqKHkxcBqZNsIWThzZRrCIA5eL2MRfbUi2Gpa4
uXWuq2VhBnWFoMUTIwHn+T0ZeKYaxZXuZ9lz5w7qXUitWrAjhE5a+tE2eMFTy1Xz
KM/uXGRlB7CzYkNLxdbGPzYy6feYF/On5QWnp9+pmjMIwxlpyW2ZrO3DLIxaueTB
xM/xVCoq2ZSt62r9J65SHkdbA0C+x6ypj3njWTYzqIMP43HN341SUQJ2YrHbpK1v
1h0Z4Jc3cKE0y0b3kxWh3VY/3r4qEiBtj1Ns+BChKOEYsfnmtMVPx7v/XTEc7OMn
8QH5uY21endHLxu2IIWlEbtV/WNq7tVy8iA7/65ndEA2WXUexqMvAXjcU6g2G2YZ
UnhY0oPHo+I0vzmWuwNA+nfQvx4Kst2Oi0SYNlZ+v0ByYGKCzM4Rm5Nloq9+9i0v
rDB009ebTMykCGOre3ArYG3o98ZF3jT/hVZMxYfAZYC8plA9FTnaTCvkFoQn6kFZ
RT5UlQEjpxguGinMpTzK4pm5HA5O9nlrmI2U2kjwsoJntW1Eq0LP7eUtU019KMKf
MufFmUHdYnh3C6Rtz5w39C1OjVYL1m2BjKCRbHd7TAXdXr0SUZgAIhQODB4of7L1
wn0mXshY7vjEB29oUMOK3lNCnc/wr6UTMlgVt5GSjb9ZeXmIM7GtVhAXK2YyevpW
wZfTX+Pib/vkyDciua6yJ+8z6K623gwrj0MwO/mO03AXvHie6Yyz5CYOiN4mAQiN
ZrWKY7zuOJjc5gykFA94djHn090n7wNVbTVYZEFmD1OTiLn742NyStc5aGoJWXbe
dIJRyWEo74PGGA45IiQY954asUR2h/TY6LJgozlQvY3Dm47Gie1B8KUWTD7ky7Xa
HxXxZ5PpiRXlscaicvus7twdTo5VI4rS0anA7iKc5QKte4O/Rp8g2YfZivVx6p2R
XK3Fo6a6IthvVH08vNRnmRPWsNnG8FAZ9Rd9p26Az+6h8ea15xcxl3VYZrU8v6yr
kuK4AlJN8J0Ffzo8pPfkAE/e1y/ZW+CR6ia/1s0qrcn7v1y42oc4nUG+HMk+KSvc
z3aexrU7g4tvXbwvhyxxODsPNEArJUdDCdpeNU0Q+hJagmP+fu7yyA2b29fr0k/m
EUYUG93WDnm15q/3M3on9b7JJ9L5Rr3NXO8y7glg6Qp4E3acEakgTMKn7wql1wXG
6tMaNEenNtY498+xmP+m8i3vqnWqdg6jXgRHLv50SWMvHK4Cwb+v5xkORfd8uN7/
2GVXP89+FvoCceOddFq6Z9yM3go73g9xHodxl21IrxXmr7olorlv19pTWdGjUTqN
+KPuLJRhQ8hDHGNLE+BKKSiBsS04Grd5+VTC/cdnsB/6cy4iXvlwfNP+q5LEjlNh
fXnF+HWscRpHDeN2QDxiVOrsdq9uIZ9Mm1mPvYScVPu0iJ5WQts7n1yGpqDDOnfw
MMR+Kvm1DiKFsrw2WNyecAZh7jLsiVAvXgQ/mW/lWm/bqH0bIwVO0AAtSuhczdn1
Jy4bbiCMuQ6oMCMcGnFjuGXFi48M2G/xdMWrHXtREkPNVLYW+LNU8N+W7igOxWKb
G55nxAoMjS+HhBMgpJ1EgEG7jnxOwxoBI0LXjlAZl2d3Nx0fQDoac40QxzJbuyo1
6reCYcVFH0ZjqukFxLuGMjvJ9l06+f2ltBNBwIiBQ7B3YS/mpc8Nj/PenQ9zPV51
AFv+XKSz520LXnJiHK3Ft8UReu+sfoq/o8zi8qBhH4847IqSTHU3aXDO01hy0h3b
FeJ47FsLvEXS9Lm31A9xAe7BmQ1cZEKNV2d6WG3MBSr/I+mxmH0PEjeUZhHhXsKR
bpnRl65L0s014Guw91mCs7CwafWU5+hCmVYccP2OGcGxvPTdHacE7hSE0pd5fFLN
zeHSIyGo+IFPQqRMRqqjAC/jPqf47Qv84oIWHsxVH1t98bq3ynAeTZgk1bBUAoK0
Nxp+FFjn+LmESFyMTYKkd6oxqfkwC5DItFXGZ6E/yDovMwon8YJgnULAnSM+6wC7
FQN28+h7eW95bva2Qv7tmAftTikM4201MgvjW7fcJK3yI85iLCVP3rvVhVNJtpav
QjwqXrZxdG5Unu2TFwIx00cPJvwXDpuVN1rkk2waDHp8a+R0Resd4Vu+LnZPkVXY
fKsJ+RY8iwbz656F3beJIx9VHkj++75l0rCL6QUO7G0ZtGkNHDhijzUmncpDWmjF
Hl+hFuV4ildsovxsyeIoAR+dsUWejt2U4YSNZh1AToFQUMbwDc+tHbrDrjbLwFya
nCxMtNSb8ky2AM6ZP/Qz/oEmkggzJVoqaa5u8mw8ckBlew/lJx6pfM9duD8IQFqe
4sQKoHeG/FyNAfAh8d2kznX4Mcvdj4RqPDXQh85G5hasjHjhfna+fyAGMXLiBUro
VW/IqhLsWp0cLUolKl91Uml3NpBzXc6XKrMnwzgSnh1WPcl8L6tzb4W/LVEm3fZz
cbaCNH14ULdyzszmeGJwKeRTn/2BZSxcMaTGAmxae4Kl0neAW8mR1KSU5BQoY81G
+GSaY18dtVd4g/FmTGwzTQjk62YFySf0fZ0q5sAlwfgKnAKA3hZR+qZ4SpY2zTXR
Xxk3HTl1vVO6K1h6v1yVBm2MrUWx+cPFVoeTQTiTpHux+KLb6XPJH9EGpoO8o5Um
ZvdQCs/48spGCPTXafYBMAoYXW0WKahkB/YvNo4PR3jZuHLFG/gCaEarl+h9aMWN
UrSCgT7X6SRAfx+zLm/3NnfZYYM9PeYworAsqxZDKABEaEQjpGnM7t8cthaYG6te
B7n/Wq9AUu/SBvPNlawZV/2oNQpCP9hnz3lIBs/QCvTAQbkQj87+jPuDWKMedvVW
D3Gb8slLf7bf9A4HgRjnitMB5fOveUyeJaZMHCFybw+0Ht+jsi1KMYjUMJpX2PBb
QMN+9wqownNV5R12pUQBG1VfZLBjczKU+CNnc7X02SN0lxeV48ymp8kt9ODnjHTZ
K5IyzuboM4qrg174CkmPpOy2xy8HhNSBA5JCYeHPUmKKsf94t6EnL3kZlTIdMYGQ
DcrmjImuZRuBSKExyTu9ViO7JpK9OTYx6sjfNyXMoB4qsmfC+r0WaGvFNm1EqYpj
fxkbeVpMYFFd2P85KzTO28frMmt60SB+DL4oxZ8ETENSiFu76gPy/hnO5xkO7+De
g4JyT/jgvnXPhuoV+dNZMMJMcQaTtPR7Vg0rkD5ty4vOknFErSDaUORr9mSAzJBX
INnHU5wBAqNuHCr2S711rbdF/30KKFHf+Ttq0EuUvXyH6+kz4/+sOLVRCt6aGowV
undUS3jIQ5Jq5IOF4twMakMHldglXGK4Ql2ksDPnbjLOPhsISs4QYn1HD8Izeriy
m8d3N/PxNMIdQaEwppDilgdqtHtbT1av4ZkxfCWdGcfNoz8GzlMCfTB+rTcJyPjH
R2f7i2EWJdhjfPaIFG5j3yeDw/pm+8sAGKvBPpW6jvNT6UICnpcHe+S5Iq/5MS9W
+/I+8MRJ++P+cbeyPOqVF9uI8bVRM4m5vvGKrapgcOHP18jO6sGp9PJMijvk+UHn
PU4YYvbBCUyjx1iyY2xviquf3wTtZwXrEZaABtHAGr6j6uysN8S96LTp3cr32mgE
UgX2USVf3dO4yrdq7GWh3mAXV9P3MXewV8cTLYdN8q6VaoNKClJw1yclbS42n39B
LwYmOQ+oKECLUHrmMBBh+kx3wDxb5jx7XUT+u5wCVUnEBNO0F2bokxCR6OIo49j6
c6Xj/8yv7/oimOISQ5nB6f4QSHyf46JTxKvGbrUv08xfteUEifwHMWfVOBtXvFss
PH//f8UTQFMsvMGhTzAHUvii2Jt7lnaBWosF+P+QfnqzWZofzL6rIZ/3lq3J9kY2
7ljTnecUoPPMDU5kqDorHQ1iTleFey95BZgONLiJSY09j0ZPT1tjbMtm10T5zEwK
LZLvKUSSom7IuUv8rWrNFsk5e/KG3Fnl5jP92U8Dc5Kay06t9dcJkVArSBIhMccS
88qJ/wHZEFRvOjQ3lgSnYTMgmFfAc/NMmP4Sv1osMQ4Gkjnt9Rz1gkQviKf7hf/Y
GlZz4HYD7frt3gfp37QWpeZEzY8t1g92/t0dgwyBAPSmF+mItvZJOo1WE0bStyKh
h858XmSnSsJTGQ8ZPWy7kyRu8FD3qGX8pnX0i68inrOiCgqupopOtQ1lAAYDzdZ8
WEBohO2Pfq2Z4u2u8wrdFN2wWEJFs5cdkCLeZlKl326Ej88m5ReHhWXTI4FkrkaE
joS45MXXvBMknWZ6sAavXxilT/ugPEJEDeyT9jka1/pjunDvOhD0bUKvlrygSjDq
elEmrT9Pul5qnS9klvkmbXir40vEby+GQ9I2pDOaRXptvWKy0WTVl/ws8PeyCOwp
Qrs9C3OQpzHlY7I4zFQ+vzJPxvKRpSPZzSayPAKxEALTK0SOhuFRxWiZ2j8lQDyY
xZO7PQ0z1DDKF/qJN4th7FPOUCHHyCJPv8RUqhS+Wed7rxZ/Bk4RpXK/mHBLPdej
afqacF0iMww9qwD9AQN84nDNZL9kCRTRp5EY2qAlg/r1j28xDZ+SI5Cv4DpDGeYz
wn+9rw4xK4zihQY/APRM/0gCIGb7NXgh5VYhWiva7jhjpfh3rQBvyE75tReM4LlN
5fJJ9Kp+W6WCO7IrQhQnOwcXKG1oVjhklJrwwxWB3QdokdCgDkZY4uEIvNzxFbrz
SgZsvA/7IzWOp9K7J/lfTANmdyJFZGGRpwu8yynarIKUpVZcYRSi1f3mwciSF/TM
XwtRJtAFvIlaeleodXkZL9jEQqct02uMDsD4kk9jiIV1FLgH6bb6pVODUcQ9/JAU
jXKBgPOg3BRO9WxumirBmEnBckfT6rzKfG0WGrVYRBZ2YMhYxgeFxeVwY6MGBBk7
V+7RFV7mCUsjvFwMGRuQX4noic7E8SV2OKIzADhF3SXTRjjw4OsC29pl5YhLnbQs
ObivadBP0YgzPKhf+oa/jH2Rj+15AiZc1p/bMP9K6w5w29KCCTCWrcFRxRlmvJmH
iPMie8UctGiKJtSRV7mVdggdSupgaZudqRr8qaQE9UrX3kLYWNAFk/FHKljHEmNe
l3E7D+TVeibZHLiPAJRTbshN5uogtT1zGfx4zPi4DeJrKP2/vH0clmcT6jTj5je0
RAjt+u3AAycIxk8mFx1g7+GIhbwUwFkN/0tpxYxHFl9dzEs0ntXAxXBi6iT/1csw
vu5wtEB56Xihtscil2nETj7qSS3gDvJJPCuRGf4+t23yoeVju31dCSHu57rGPWWE
CEJJfqAv4k9/EhXDx/+nke0p5i3LeJ768usX65u6eKghxaTDfT9oUy72oN3SRo6f
tXOe8sjsVkjCopyKzXLK7fcDaBfPHL61CQurH78HouHYJJS7aokp/BNG5uC0Wx9W
jUWBtGBQ/nxnuu8eAOJPmgqbySu4tU7uB8PXd0zigTDbRvOmxpSNJblL+WfpKTr3
4Tmiinsurt4moht7rMrUfPtaErKWf2T2lTZjfqwuM7mr3oFoBWNlfE/CV5DBsn6V
LmLKY4RIYetyp19r+mQ5eS3L4JrObTdXg/OtO7LE0M7dy+sMN2XZEx56c+i3RDzR
ZGRbUHfCuGHFy0nNtJ9b1DB6qL+IxurgF5Buk0Kmbo2O036jZyeyJpuOza7LCjS6
YvZsk7huGDJSgMEUtnzBxQejCNjTVMU2mKqShor/iERF3fRco8Rp6yOVa7dd/RuB
1rw35puwDGzqtWBJLLoaUzzpEdF3goo4hd/VXcrWXtTv4QMoV9PQCrkPSoalN7LU
OIKfLU4fid2rA4OsEXg05JpqH4vcilGOafs4rhnxKaRzY/TxucgL5rVD/n4MrVFm
a4Ky8Ix3Nx03ujtD+dw3a28P2Y4+obZXHqg3tSuYGoAIgY5sV15RQyBdmfQzOdDg
O4sIu/5NmsLCbZzkDqlKvzDHdnWFbcTGfHTpHR3TROAhgA/y+QkCf/pbj1QhFqSC
z9w7JMw43X92ogJ3F+71uwBhxHO/ZvkSBI85dZM3re7RTsk+Rlr8Aw91hIhAT7Fx
+ydhNCrjyPjr0aU/0UAd0b6nwAC+778zn6YGkYT+WNcTEHPxSUDLPaCYC9synxz9
4fa82+oiryP2H/MVAIMaKPuMWNz7ZJ3BscuqcMIXiO7+/aU7w2Hgyuq5bTBnojfB
yXH1tG6FmiXtFc40NHGB9bNVhdMkmxkA/r9FSRRqgjA0d1zHY1vS6yQBzntGEUB1
OK6cvdy8DPhi8pSChh6y/r0SjdDrz+Rai2uzSCqgGn7ViiPAkTZwkPkKyS2rzn4Z
gdq9W/47f3IQJeglRos+vwF/S4L6AYVWngw+wvefbeGyDe/9gjX8+V6Mv9IUflvt
8FufiNZZ7679QMX0SDoTLNaQdUT+RaSUBglMFNJmatkB06WPg4P+ElzgVCnBM2ev
PsQj4iFOZ4Cijkg1vC95cSDRVi0O1i+Eq38nfJ173v/eKFURTDDpz/+AXB89I5QE
Wiu4JDIFqKbC/RQ52FnbmkyipgFZH66zPDs2i8Y7dwB0892+4frRRG9CJxiOwCqA
s+uAYvlJOdpk2UigsdK5Mv3quPie+QG4zSDZQnTpLjLf91oTHadNu/UaFvetv+BS
xV95WfT+Y0VD8ZT09tyqp9FDx9sKZ7myNYCZ+oxGSaqwBgRCxUzRyU5U66YlKbfc
1HktcngLvNta91sf3ItlGPBWdPNuYlhLXIHWFX31yroUk3Puj9Q4B4wVdEJ0/sy0
f2Rua9MchTbEJzS53qE7vAA4E6WXnCHl+zEyWj4U1F22Qlo1g7l+lpN9S8IO4GGL
vpXly+35whyWOHvw/7y4rIVAkC2BIgSuHLTYVFHk8NPeD8ufQ59h3sMLYeEm0fH9
FfqQ+PWTHn6jeizJKmJBUL10lWi83kZqx7VmAoLksZdxALJ2KOZPhpokcyOgGeCt
AFvlHz0kSzgUUUNc/Bd2cvNULzK5TOOFfQ9CTVfZ6VfJNb7dw0Bl9X+rS+SyFdzy
1dIj2PFv0f+Zd1HLfnddUuXSvSlqReVdr/V6iriq/dXdfekufzJrN/XpWIh5ToAV
NGT8bO7gPvQIroIWmBnnV85StzI7UB5ZvftKGJ8ebVYBKLpWKQYva7InDM8fOMQX
HNUKID1+fAVCVLvU6mNgWu7ACvB/3uqDsMT2K5x+w476u2otwiDXMynem02t1kGK
DTako/SzzUNrRLXdeMcyE4FhHQrdCnX9IcBYvsqIOSx9QcxkLCCtuJPu9X1Jz26s
NRiV2OZJfb0Bck0/1nTKt0BREdXBT5vt9kbgAmTamfYnowI8Iy9UsaGphliT7hfK
Q4rabUn0yC24EtUfQkDAgL5HNvb1XJogMgRhq++prZwVMGSU8L6xSldgMcLmpI9h
k7v714UafjyjXLry8O8l2x9Fid5MQFziYh2N+SexUvnaOyfvbtXnlE7zl78W3lUi
wL16qSSVad6WRw6O3ue7qMOvNLSpZvJz6Ii7fVewCt4wudtaA48xv8KIHfX62thg
c4IwxMLm4mpkzVnfkt8hQS9BZObvbJPfuStWHSS3bAK+oS7ib4sfF6VUUD8WDYB/
6Zb3HFwuWD6c7NzOohAwjOcz0YZjVMLpKT001X1FkmWO2MLdd9sUu/QnzqR6LEir
NQdlkyLCIlgHfiPI1cFwtVC/KEZDKLZFrz+IOvdB5KHdcXpJzeKvi4HEQxFTQtzu
WJatMRJrWelEDizm5m9CafzXU1bzaN/t3aQpZrpztQNLQtlInlw7TPHA3weVPdYA
9ye4fvo8GE28+Nn0nyyuI724PsITx9BgHmomwbKg7Z97m33ogDAYTCiSggqAnroZ
GHAXFuJ81CKRlIIkaAGUgIla7HEWIslNCfbxlGBa1mOS15JkTJ3FjZtXOCeQgtR8
PdEZehlSjZ8T36J7ECshmlF8xs8ctUC7JaARMrNBQm/ihkx5xX3ZrUjt6yD7PUGq
Uzk1UWkuLG5Xtq1IGTDC7UJRDfSlFCnJjJPVCnwcEQf5/S8T0imW/eiyYqxlAefA
LJuamT01yqULCOe5xYfHJU2lGUzU6et3TPBKzrWgfkmSDdH2sq6weARZwSD/2KI3
JxmwQzd3PbUq4DskPpfao2KN91HwYf/l4cS7EguWcLvr5XTGo2smLpYKH57YOiVE
zg7r27N15RyVg2CFQxnb5ScTy3toyPfc6+675bqDVkRiowFd9QDHG0itaKPMP9J/
xHGMtd20nf5jpOX3lmsKwVoyEx+/JNiVHAYgysKPgC1eA24Ka30LWePXAwTrz4QY
jHa92KUAc/XOnlKDj9I9gLNSxKucSaeIPzA18T+3LytrkHLNfUkkXDkTmGbpOFan
9dJYpYBWF5AJeA+ZeqAZHkI4cq0voIk7DcyMqDX3nx1nEioV7keFoui3skcAr8T2
DJI9tZhiM59qmgoA8kgVAZ9hPFMoMTxizl48v5rvSYBpDHTrPBi7dsixrwTTg14j
oBtbnAbxGN419b8CUNrs1G6VfQ1kdrN+Cbzfb/yjn3XJmnb8mC/haJJTWOykyZbl
HMPwUs58PJaCEaJpxpPLu2uJcno12O9aNVhz2/kvyKphNT4W2g7Bb6J0TN4dhPhV
YpL5TG6QkfU0zDyBwSZLS4m2tnxc1TT6iun0sogRwE876mYZ3fLOh5embaj2fHXU
I2yBo5LBXkUU9MS1qpW2GEfJvV70UShxzO+p4/VFIZI0fby4dKRkkKY0M54D6E1G
BLn30r4aiP2jgTk6gNLkO0BuGcDkIDPK6eMAF4ljHNY9Se5dwRn4PEQCqYJs8jnD
ryYB3oNrOBPpgACrcyNox2kyeOy0C/4yLY31HLzIrptX8pKCkWEqJdGoVgJeXh28
LegQqD/9X3FSfFxJG4ry2AYZFTXPDK+bKo+5Wy+lHPMKxXRZMd3wBAN/6UgNP/Vp
7O0Js5NhMkN5s0fr6eYUx2nLiBXpHlcn36CI4uM3F6JrMw/XRjm3Og8jXvXGkEC0
/oJnv7NZdQ9Vy9l10hCmo9KN/ePThpYtJ708eJOVh+4GPdzEBmy9GVXv2GXwLF6y
q9X8Akwjjw33OcsLasW3fvXbzTjy/b8ZTq4lPNa8YHay3v4IK+T1w84vqe2FnZpD
mGYKfx2C6bzeaJvyyweTriWqz4atyNXWCxRLrlrnH7oPqo3uEqNdrv0v73Bo5qI/
4j0ruwx85bubUMb1yOaJKyiH+YqTCv6p4DD9ximUzuRFT9XAOc9lA0CBE8l+vgTj
bp/ums1b1FSdEhtTpAvHPx92uSUaN8hT9Mni9afUVak8fcawwxe56/g92I9iO7T7
8C9hMr7gLw4LhrgkA6KbylYY/nbuxNsgA/w9O5qf9uztyALqI8vAQdNyGntC0wRm
HHI07aa2ftC/y4pivRwX4KcTBh3g9XR7/DBtRhwbgU+nkPhqVF1ZA/+XDJZlK0fg
W4Zl6mZHRrRnQDdK7PqqWzmLZ2TXHtztEWC5LNTbkfJrc7cjC8wSg+w/6VsDc+wq
KQ1B76h12zpihEfZrkb7JEPbf/+72A9Ctnd9TyWFopPEv9eKH3wje1FYaaITlCUo
Q5bgwiCy7+nBZkujDy5Ytuya26kNDnEgHBdZy8rhQPCmCfkyn4dp0qNvd/qL/O+O
eOcADl9PxfD9hfktvdM30RU25OSg4rYy1AmKJ+g6LzyEEg4WZU8sCIRGBZW1uO93
Qa0oUhYPpihMAqiCEeDC5MOiqEpzAiqJRASqdJr3n1nJ2GeXR582cqxEBz86EvUD
5+loitbJ/euOTmqssxabEp9daep7HLwVfx1MTQYyY9RBzucPM84z4BUWDhWnWAWS
wkZ760Vnvm2puCU2YlK+riFUe2Yt1peuAjh9GcoyYYR/m+7v4i9ViN1/VYyR1lqD
PrMIfhfkuUVHkzhcAwxjmpz3OLvJN7tVU/FgEGxtZbmXeJxFs55BJgCN8Zh6rOrK
VPlHbiTbyF1eS4/D61FpS2xOEzaRv0Wg1ZJbp6DLLcsmQo2crvt36//6rem2qccO
1UPlQXWB3pYDSc8PFNU+19NmcFUcxzSgJvGvTrjEfI70xycr8V3BzQh6IlRFJnJG
k4MLkqAG7j7TT3BCQW83TtluFhwGOkzE06dylU+dfPr82JMR1Yl5IwwGnmq9XyWB
H3n3yOteYAghXat2clt4tnN/OTrP41hnSUPmWRpNTlrnp8tIJJxju3i4hWTuU/rl
RroC3BCmZCF/46WFYDQu5mO6KGwiwpK4lOE1b5tQFEmWKkRo4W+9DyUXQ71Cbgk4
tyscQN+SOfyRRdDPIz9YaMqf/DCdxfftVe+NQ4MNBa43JIJqds/t8mAjPUg2Ukiw
TaC/d0D1g4lYR1xBuOK1gYV4O0i66mTO4afq4eVbcyaXO1tYNsOK+apjx2H/2NRL
KurjfJwWRmrBZ0rKmIoiKcMLm34+/rnGi5jllr2Q2LcUeApNfFMdUGvgXE/fcoay
A2nIxlw85Bosp8Qf0rUctUx8g/sVgflNPEGYxB2eDv5xawQtbZMkeZQ+cqhEl2GR
V7FrP+Za5bw1qZzd03a+KDt5g7D7EDebpHxneIZ3mjo9/TjRwV7IpS+2bcZemLxC
+xG768VLh+hclf7OKAFjGSslDbkSY9Gmy8JcUHwhuH4dqLVB/gV+UlBBOtDjvwjc
AXPJlI1h6IO5TOGO0jGCm/2R5ApOlRYtpEQAWAVfhn+RodqCwU9rsWrjWJAW7Lnq
DccaTLYj1CogrKlaT2LrGxleyH8+V3bXLNnU+TLNER4C3WiW9Q58jDJncIfAAalj
NtkSmLVAvsuTedw5vm+UGwA38DL9DAsMcLF/ZfRjBAE+Bwsjvak27tX90VGLSDiD
OtyYy+q94CAwy1mffzZ0Fg5jTutOiskmTlazkcH22onl4Thm2kTt5f34NaNkE+hs
Cp67PZxwTrhamEywtj6z9RkZG6Yyl2VpHxGfe5cqHf44d6dVtd9rIDGCGy+vX4lC
v6H21w6f7wqXFmKeeBySb1ez75D2cLIwUGnOkeVFFJWtWDoVSv0gyPTw6MnmqIUt
obO4qnCXcEnUc0zXrPLiiX0LpVT35P9bq6AFBSSlRwBohc+W6BI8ZzRTRbcQPUT/
RW6+f+ljfTuuz3KPqweMoQtHE69GLuNE6RWJmBIsR2kXKXvQQuJfhHdugTFLpqVI
UFENE3yd9mrR4G8Cmd4bY88v0571eehaSFWIj/wInRsU6zIKj58eRFixDHvShowc
8H2Boc0qu7plDycuZf3n9PI94PopaFcrh4L9E6Zq9o7fHf3RIrIClBe+KCk+iwHP
5c4tEwCrOG1bRrglSZO4AiDERJnNrmSuZI7Ygl889SiaEH8tyn4Yn/SwqLxTERcK
Efijue7YQTYl40HxYeTIhg0JTfeAZT8kLINlNYOZNNdmm8+qvCsGs8yDEyM64lyV
Xp+HeXpFKyUOIiVC0C9NYm1sw/KWN3xpffFgvmbapX2OlEaqvHHgbA093HVUtmiU
82IckesxRr7MxSKgjRUH0D0wHNZVahSFeAL8HTgZtUtKEADpq3oyEJb2xovfyZXT
m5Wc1e6HKrZ3rfG5pL2aqz1dqBAGe++gm/xZbAOpGrLkedCLMDAK2KVNJOFumXux
5rTRyKx0hAPaBwIxOkUvTvkhlhud7/tRq4G6tgTuCXpbDj1CPl5WRRwqhoJatTD6
t1gJLmujqbea8tr/du2L1Pg5Lpt4lF9gY/AHcGYShHMLfW9xjcglo5XfNYuJFF9t
2d0pcVDNUslA+NcDT3anxKkKPtAuhWvNhGFDF29Rj3n/OGyqG5g9B/dybdmAIuc3
dfTe4o7kJ/wDQW0Kf1NUBgQYIow48R8rZG8+L4k+Bsr2ozHAgAmGKVwwoefhL0td
9MKAnPQlTxUxk021fBfwoUOGg9YKG/LOHRVsDJjDt2tkTSkYcGdwfJv7IHV2lHMT
gNp2FyIrhDI1eCGsHz8etPnPtaLyktwZIVg6+svAaOk1vtjzaqaFmnSF9Os7Upwp
KVbb3p7KOUBj7ek7C9DE+XNi0/bgGf4JuB0ATD8xo9H994HSmLG4ani8n6D00k4Z
vwjv31Ihz9NhFV4fG9Cu5x5VDEphMLWdwOORheaGHdOcHdngAUQ/w8iOmKb/XFdb
LB51Fsh3SumZPPcMZHWq59jT0ByipKncQAsGno4eAf2iC2t7mBkwPQERbbKlnkdw
CoMiBnKrxdHtxw94sEEN6Ne8gKUF94yGUelJvcRUsTnipTK+6iH31kRFMnde7kQi
ww7wzo2QqTfvlRAVozuGIynh/kQ1Qkp/sla4EbSLAt3vL6pkd4iCWrm/fqsKkGYc
r7v+cujdTWRnGw0716k1ahL6Cl2ROfPql4YlRJILCGz+BVMXI+WNozbLfqO1gRG8
sG4Y2G1H5mYXC/wFYmsVJd+zo0ej/6w5OHKzKHi7cugzNUIrMY/d18ghctvIlEuF
r96NP1/r0zLRr3b5xrGJjRNt6iQ45Yf+9G4QrKh7/CdTf2Bs7GSTyShHRl2FPJ+d
x6CbmypgbGh3tU+V6XDw71xylMt7Bb46Nl80wW7qwPsl3OKpv4XpeoP74zFdrr8P
+KOCdK+msEaF7Z+bGxb5+g6umg9/yV0ud3EETDYxfveAuNS+kaBLRWn8h7BJtDwi
CjPwBghvsni8rE6uG/OZvPJ7O+9ZgkVeHqv9NNaVFShP/8ikWm5fWNLnnHQYvBWf
qvNAHOekvBpqggPXMaZBsXztEhp35if0DtsyrdZlXIHmniNLEikTez7ccmI5Yv92
cxgQmvcfj9QVd5ZHzfDPvpbYvDRTaBaf7+tdF1pi5XDDqiCrqj0J69p5MyAMerOW
/ChWep/96iKL8jdXCyCutJgd/Nrbit7niXr0Jym5GO8MUowP9fBqsFpjuswsg6DM
EsNPFC3B2VLobz9x7JKZFJJVDe9WVbdVgoTKAJktzsqClnsysQn1lCoC4KE4F4vY
QZIfWtDrXmEv7ZWMjEAs/s6IQL/D8d6979C1WHyUeXQdjO1TWtsuIDskJHMmjZya
sleWY6PmNVFvsGSDT2lEywFBAbBjk669fI7TLqTBVrRx7gmFymtXOLUHBQxtr3Sp
nPX63z2I5v+HqOwxt2loMMQUxDmoX2O7FFAbWWOVhd/4DA0hkn8a9/wfrm3Y97YM
6UHJP5FZ6DI9O33esQAGdX0iZwbE+2wLVyDdis4GTyrI8lXd5DvVGnWlFmVDP4Xb
hBCeWfTNDozsYgR694kFQ8jN9nr5WhRWG478LQTrJYvQu5A8VQF8y2picQkUnsBg
mMmkNfmrYreWodUQLrcDzrR/cyI3xmGtcspQUWUuRVT+FSaJQOPZOk+X+GXLgtdk
KtPCvzyJk1Y9Q2ZUEGMPclM7zztX8TbxwzYoAeFmzcrXOJZaCwiAd884WIM406XS
YVANvnw/kmA3ONdor6KOz1nmLAmzXevzWYH7i3bFor6YgbetCPit8W9R3FyEZMkG
ruW5URJAtORBJppa3Np7q5MPMMzeXbuAI5Ly6tHETdlAhs7vd7gRevDZCdNLGvyC
byVqAXzF052dqb3f1es7HjckgffE56olhjOvn5WMTtO32/NYlrK5ifemF+v+1mtR
nUCiSqxb6tkDMi/xdShfNfMRV1FxHzjwnEsigYBdqcf6Glp9hGFR56pTxkRIwIxq
8iUOvarbHIDmW7u6IuOMzq5fsv3vq8jTjEnGqhRSFhUP/b9GEU8sqICXexoHKAQD
qsspKMXQ8ZvqAfoH/3RayESjK7hgqwQDb83pzrS56mzXm9s4ZfR6Pr0toWkmAFWg
62ePzrwu4bdjyt2O8132AvRvtx/b6FzR7GoDMfevl9JgXssRe7dhZRVE3mz9YRHG
oWF1rxZSo4+WnTs/HMC03BUSQExYyiJFp0RcrIY+CjnbrWJeTUYCu5uBg0yyBjR9
M46IB4Uy9K2WAJJaqwgI4SCAiASmA+R9BoiBRbsTBmxWviTA940AgKHFLvPGqGGK
utz1MKiCcwMvKbSPmVKtItdPKiEObVnZUZ5xnnPXvmEFUBJWSg2g1iLDJHfXz+OO
Mr5N0vQ9FodOeL9IBymKgiJve0NqBCEwbiSC4VM73NxpTxIApE1DM+20tkdmUU6t
eQ01e9xZ3hANedmuWDtyEU7D775LKyLHrOY12lzMGmBEs36vrfUNBpQkxp36YI5O
+bMoPNhwukGtAwjgNUiMhmAzZ8ZS3ZhYjYSe9HBbVwlkX6OCOJuBCInaZtwHYFCi
gtzCvmrYkKb4rQnOLaCk7nrWt7wf1OYPygfBx5i990wSYY/veY8Q1aNLq31YJ4op
QZ2imXitY6I4jZo+bY6qYXdfiZVnoKZVeO6sIWPBqYQWMzMPPjt3AhyrvqxeF6O/
RDXHfk5ZW45agWZt9/c4p5Sw3tqQbWUm64zc2ytCRR3aFTR6lTGmC++uy1O+Vd3t
QPzCiq5HjKkU0azJgkjDtaJB1b9ERmpXzEBC+d7GvbSSlVPhGPwA2bfIn2ak62Tt
W1JE6t045cup3bUTU5pi7FZ/ud27jmJBqGA71/3qyLzhmwpH2EV3Bq9iPnMayydT
Yv1EK8G4PU7Jds5kg7rqP+HPZo9Sw8rUu0n0+/NiAIeQFIpaiVpH8MQBKrQR/4Wt
I1+it7XRy42EmJvC9mut/WHXr4DxT8cJaKSHGDBa8Qy436m/t4H8F0EXJVmPyXYg
hRezvaOn9bjcciKIze8a4Pr9GGTCWOK328SBOQRvSKEeFwFQbWJNQxEzFRdIReut
PDKfxXc7fmx3YT0fPUTIE9ISwHiOYUOcWdcxuDPNw9NeYxxTonGcvKeQeWf5awWJ
1QvSrJN64cX+UTBXZ84Sqd8ZgwFB/QnawHgB+YQ/l6Odhic4XKa9itojkoojq4Yx
xkSlOvmkTJwxWQwbioxSESv0ZngQZSfwd0zf6totv1fXbPKMi4DYHCyByZxLEllQ
2vkNGwGtiebo+47/9BUIyilGDg0lzRCdakBCWx2DUKG8VqjYhsrWbREgnBMKWh81
XkCkYWSmFj9sPPA42wDjRfxWH8sKwAKYcAHP5QNf4AgimfEupnImQu2Ly/q844Bq
QoZ33QUAl9jleCxUCjQupcADcp7Z6+ampYgtZoaYyj4y/0zfC4YdBclFDuFuuxh8
Jy5R47Bj6vG2D6i6/uc+KRmziEsKh2fBvxBJ0Cp0gR9Bu+K6Qz4EjZfrFFIi0kc4
dkLcPxrR+Xz2824smTL8qpK+VBLpCpvmXRx6xbmbyUi+oq/4IZvWW2lBMsvNy50K
yZMagVURZrwkutqWRjqnCUDa6+XPSsN5qIWjuz9R2LQ7T7b81VVNYp6cWWBOsa7w
Ll3Q2LByLRstfBc96msGqC7OEnewylk6BIfhTfvhVHTp33iCwRAe6CmaEuXICTLQ
qZwfau1VkSbJd58euBQIcMXelW0jLH/UVTwMGfbT4cPhDJAQqHSVNzCNo1XZuotj
WcX4o/lIY0FWwtWx5i6jzCbCWAywYRFk4FSOvDiBcc1FAIBxjEybKR5Vktn4V+XL
Ig6mMD5fR+yWN82VC+7hCPRGVBRUat6Pk+gIxz2RjgCeyTFw1NtZoqbssoK1r3u1
2Kv86gHn6HE01IM+ryO0z66qg21LvuJE0nIg1wd9xeLoF1xqZ2tmEFHS4j/HxPzE
fQ4E4lNf6dRwyLq/edIDIIdwnS4jvYW8jZ9rFvXqzusaSAgPQs3iRkAh9FJuylUn
xBMR21wP+qgVWpAMqbC6kHxSAp/EvhcQNO7Gdde+3jmOefwuyxYMKsH9H4Rq3rtw
Gyv4KP6ZKzb4tKxr2/5sDYVen3REPWRFEc5sEgfW25KkcWKYb3yy+Okc8XmikHGk
dYx31QSTX/Afo2fqwLrY5m4zGmUl3mV91kSV0bombowsPp26TKrJZr/kzGsfHMBi
cMVaduLaHhFnUTuMVsfHth4TtLAdLAMBcokzxC0hGcV12a6DGC/wqoXqLCrZBAF0
hUHAvsSIB+Fl07Utj38nhow+CSRdDcLkB5qr/iZZNtLZSh6zAdZ1t/+tj/OO8pOe
37R3/6t7HHodYTIOa2g49Q9aewmESez+yDSxSKRFqMJGMA4B4LlBGosiMGi1afbH
TSOzOEM04o7vBn7h0bJeM/WfqQ53ZgcMtUSYdfYSxrnWHk5YplrNaT7JmaYwGFaF
GF7S0t6ewyXFELodF1pIWvecJDnQNPEyXFLyDNcnuppHoUKzWkfIReBBuJAoS+wX
Slw7qb8/9Sr6i9QxiKWdXj8cbo4qt7bPdZIteN3VeKpy+CxWvJ5Wz+hIeZhTRLQa
d/LEd6TnJwzn862qPbKnDauuElyCdTUDss2AtxwpwIGKlD5GqXcMhvd0KtqE/8KA
8IAfY50aMlcte0sr5IBZVNygZdaE6YugwMh3o5mCn6xwsSEL1MWCzMmF/ORHtfXK
ZnbP3fR6UVuuO/AqItRRLqkZNSdDLRENrs8HEY5I5VHAnmZHvsmDFNVeGVzZ+ex0
UsVdeTIHX93H1B8ebopVpFGWBI392YUgkKHPF0sazfXxImGfQZ3qTJlYbnxq6Xmx
xSMvCrEnYu8VX1PXVZJB0WzS/iQAJyKE2l8SicyQLtXupeBPGvyct0m/gssI57tR
JDVT5nUv7wEeUsiraN16ORDryJy/lAPB8DFT4ItUGFyPuxhhJJWqFEdhh3fCdYIQ
QpKcHR/VNZxTCyZE5KE5Ab2JHVHf06tSAN1gucp+QZ0FMhnM5M4re0LEP0FsgYYk
ldeKZp94ThK7afQCjx6YCXC3RWEdu7hK0dVZhEj7WMfCnZahiA8/vjErzzRvZIEF
N+VpdAXMCZ6vlHEBRYTJvfWKhK7mJcmpVO5kXXiPJDni9BduedNQHcimg2eM/lgu
/fkq1QEcjYsL2xSrW9adNifBCh75dT/o4SD/YNvA95+lHc5K/8r085wW6D6filC3
kC543kbwEiz9CT0Nuf4foU2wbmt3sDwCRYw3XY/qnBnpTkuzxuFW5nsedPl1RInc
WThfepn3iZ5uFdLFyINUmhKRNP7NIbU2e1CaUC6WeS9Z3fiWNW6FiYDxkxpavxVf
KsG3z3ibgwi9JOJh326ZxZ1jDeJmqESgiC6b+Lk6qG4fARAErCZo84fN37+iLHkr
1S1PjCH4uLNz2hKgL69t93hNlrn1LzEaq5ZnNvDYpAC3T/D9J0O4+XhgLlFL5PnW
tm8K5UZ1if/Al6ikxn1nm/+Sn91q6fAFHLx9GF9A1CKfHKj4IPUEEqnrWVmDWZKI
3Up6r2HOO2zMaIY/Zf4fBMDN0OECdQDgs8N8tEOCsuU2eB6X3oxw0t/xJGfY3RuX
opgAF6zw0vDg5siqN8+MhNXTGN+ROucG3d2fHLIWtmAhMdB+IMomrhWmQMvrSP+O
t/cfHZaQ7PMlWGGRygR8NRsaGs1OunDvDl3ACuU8CXGFN0isMykVWi34OIof4pe7
693+Y5XXe7TylAgIzwF3HWnLuqOZ5HiCGO+jgMbMoOiJAFyd2lHIBcMXReUuyppt
nLoQDe+zgC33bH0Lqut1Jq6En/HNkupPpnKlZgxu5RxXOe6BEZ9VEX0tAbB/yGJs
a5mD2NcY22YoQy3aX2BzLnr8Ej1UzBPw7OmMFGXjMgHh7lEUP3X0EM8xXbHCDtIb
9GB5vbD0/mWPUBGjfEkVPJ71re+VTBmNl8y0T2poEoRihVFqBEEV+jNOJS0HvAes
UAE6mdFuxB843iSNv7XoilvXVm5Ro6NZg1L+HWV4DSM4QZy7KTB3Sdvg4CJoD41v
RX8iSkChXYotARW0KyHMt0Y2I6jloYimGcY17TRDp8vRhWERt461j8YMfMTT6LdK
XlaOPVppll17Hu+4lzJncOpdHbd0zDfoU/415cTkcgQ5d65a/nKQlC5JYA8qd9GP
Xy+MolN6XiPiswavHHZOaENYLontMB7c5zOlzTd5NkRAINDLuZUxu61HMnu8mBiL
u1RPnZeIdwzq7FLrLmgAikK1aIovsQvDPk81f+ZlCBt/aYd1fCnnjSN95dik12Z7
5T9CZLr5vCBK27vSBAXc0NRlvmjvqV1e4lTOoTnmMxR3FBp5+6oKOyKpb4xFNCoy
C7hRQXsdMYzwOpS2odQQgcHTH2l2xZq8emHWjKaEkKzagCgOdGp9z8Wv7nTUAWse
SAxEyCA0O1hpY9rOxLgORIvu9XhOlH/lyVPAbDAi9Cz1RFerGYWfb/VOROEU9zV7
npje4QdG0BPfJ2i2takrIPiq6vTgH6/Wtq1TIMEXNM+xQuPSZLdGfqGu8Wg+xcgo
gPaz4fHQVEOETag2sp84UZQ/Qd0u54Ef7omYolwQEAqvKrSWw5ZLVwjf8YWAFDRs
w4/01ptJfKdZBULy2ltHq4a8yAWC77vE/ljthjDeDo4rCatyU5Y513BxY007ZMit
xujcfxCpSQziz3rCdfSiiNowqgPNpLXMuhhDGwVYix/vkLTqKleGGWwll3eLLG4r
gJvwyJ9v1skjJdo+6shyYHpNopFMg5M70VGovGG+EsYdnQG4amRT0tpqqW5syvX4
N1kfUh/keYpCh46xxIQKXIvGF2ckDKMj5uGj1ZNvi/nPxOrRt5Bo6cNUr7XjBeq+
Us0fYRwOcB8G5Klkd2SWm+wOZ/yMfP5EeSi36dZ0TD7zT8/7mm2fJODrTKjcoi1L
BEuATPSEKyIv1NlQybKMcmIYJ+f8xD8wdF3niS6BiM/0EqvaAanRsYJL9uNGTWuL
i+jEsezTfvziW7Y5I+unc8JgwKanL8HvVpm/9Z6jBZvMp9DpwNRRG1quuNO5SE1L
nGpTORl8Wu6WyqC7YmjGqY8S+wI4sZPlAGHsEdIwNqE8WN86yjS58/c9pjoRISSS
7JGd3PU7q19wlyCnE2qEL1O8L8s4z6eWxnb9IjUHKH9GBA2MdEOOpLo9fVTvkyV9
Eg6NZXXwT3JnV4yd/OXlu5C0q9rFkNupM0k6QyWkiBB1YzurnN6/1QyxwzE8WulR
Rk5PFZpINRAHDuYnNMVf0QPEuMmNIKVckRXF95ZbUxQ3a+w0pKIEl0CreC9h+7pB
QIv0jc+qJNzQoO/z5Zy31jeyrZFgRi42SWc4yZTL17BhRsB1k41ObbyY15RCsMy1
ReNSuWAWBHTcH5/jY4WNchs2Zpf+twMzd/FIVEbNO4UyMKTMvLCX2kqN7CzHgf7F
UuELoGGhDQBt8v4pZdjW5CNZj3rsJVs279Hw57vGZ8z1hx9RJnzYdU3qKigZgV/6
w49woogyGkG/VmsWGuFYSe1WzX7inR7O9Iw1GD5AmKLD9Lzb6Oq95o7qPL/m6f9a
wpOj4xE478M2qOMSClMS4+7USUc0db5C0fbV1KPLg9kIeSi/sbtbhot8yHS/3N+L
nnVrG5zgGM44f0XOq2oGLzdzI2Gdz0l9HA2pLwBZ6Eqyrb2qT6Ji0SNnadeHLi/K
L05DTZfMkTcBbrUS3DBw9UiH/vUqkGMAar2K9OF9xZ1Hsf9+gqylU/qq/67L8xHx
syUXYfJ2p7u7a5TRy1blp9gMPCDT/ow/lvjQpGSQqYaTjGcQ8zpHf6qqBAIKCrOQ
oyYr8XXtcjaQiARhYLJmicsZTAmYd8ihfqvv6FxwiA4adjklEO53L5I4t33LeWD5
ewi4ay6mKEJLGG5B/YJ+nm/vpXCbtdPcBQifuIqP37UsN81lqIkV2xbxAxYMiqBD
iFMSYvTr91/xPLbFArW8CmQmKJBOoXK3V5TykDsbxs/UIOGZY0KJik7nTi95bw5e
lYopSQeEgh4NZk6Xbr+J3LuYtdddMR8ezNevTm5hoLbM9Ep2mR/gyorqYE7QLLt6
PnbWFT1d9UAorpF5ffyQVqF2538+nYMY6UG7qvfAhlpNkhBPuMMhZGT4jRNMB/QA
rKvw+VAQ4XNsAzzhF4Q6okcLAOube0JJ0WF/jAQyCS4JHy9S/njWPBNeGHsPF6z8
7JctCQN6k7C4Nq5vs3PtoAcYVg6gs8bA8ky1Z5QxlNfkWHkJB20VYN+cyplGJ4ve
2M6EUtRlUb/A0CsJjrAH6BZSB/Su6lbqT5vjlwmZYT/HHMhDCcbQV+3fl6S/zaXi
s40eG5pYAuD9+8O/0JJ0fq3DsmzDn244U8j6Q9Kbr/3rpz66Y4PecjP+sPpRfchs
8MQhxMH/mo5xEaRU4+GsJ/tRkbqvwNfTrcpUmChuREYh4ytCuKK0fn76mOX9xtwW
/hub1pFfk4CcztmN2U8LmB9M1UwO/RbciaHrFl6y60JIL3rQNLbeI7ZFtNBzmk31
a61qzNUjs+jDiOU/9nKlrZ58G9U8ibY9op0Jw8fWi9V5xPCu2slpnO2ssajDK/sF
EN9cBJwn9SHxiNiOgyVQxpKFntx5Sv53hZiX1rnRgIDsrYU1MPGBnZovL8UPJfe6
5FRgxHxdUE/huT2a0aC3p+178TDqoKlojiwuXP2j/l8dvSwuKCsLkv9kA043GJJy
OML75NBIhi0vhZSj59FLUhM1gKp36vZWJCl7f/Zp9bcGw3wOvO8Vy2VgoC0G0msd
eTtvzR9BEaQwRZX12V9xSHZWILJpO6eQq3B6vMk+vUrT8e1GPJldZ9lu9+o3RFNa
98COItZSVXTbcMPxTqmavMyhkU0wsHFKHpviHObMVA/33DuFou4ogmeGGDJJcGHq
9UXWjAA+xp023CxqNpyckQJUDEE+WA3qWPFtFEyUkcc/SXBwnnKicoOK5NIzjz1c
vtHkkQAK+pxApQ/0jNaqFXF2x4SHEm8okqVaVRmjHwWnCOboejLJ8rn6vb8SPue7
do5dZt2/2zEdGyhN79RkiVUQN6EcRURdgiCoF0MGhrHjuCLE8xeTOw3Vmj4v3hpu
XpFArFd93wBy8cPfxgnAtnYBbeSt3/pA7XiqKZgtNKhBKiKa7D/mCPOW4mDGV/ly
B/sXeOcRZtjHFDUKUAbHbIXk+m9TTh0Xqs8WZXmEc5/JTpHADRjYB1Rz8h8cf1PT
ByUMLIIoJRm/IhS6l2Of9xQ47QmCJTZ89IH1+bKYjq8SrSz7JVomBSSeNq+xLYc0
tbiU2ax8GTSPkFFsV4sji0AZuDFh/FT7ZnPb8X2OL/BHiFfa4Bmw59zoQceAQ0cm
HEP3I4X5FBeCi7XLRy3BDv6iUOOCi6Vn+Ry9zuRUaAtqQY/p44kYOcewcjKrK+/f
qUmqy/NJLYo3362lhkGCsNQUBVLDTUD6Gb9fwn8IpcpemsGT9Jdgd9ESBfGT0Maa
1C7fZVniw9Bq6cYc/3+6aTn1xqnO1fKKQ+sE7Qp6vJDULTlGyWI5jfRPu4fr1mLs
+W63pxwYfp9pTBweWP6CFiZ6BSeeeJH2xwUxEFNNI333eGyQIh1U4y25yblBcZ10
KI6FxJ3IO0A9f+2IQ81NqhvApp9zRyMSw6iIkElkzwhisKGiV8Kc8GLxZgc2B7+Y
EyPs5RyK/bmUN0qa+56SlNVp8er+RQOFkxpCw0HimyGCmGr8uj3SNR7pSAqWF5Wx
zWvPHeGJtCXC5KXzbVMjf9iyyZT22XKuONn77adR727O1+L/vJ/5ii9rr+1ovJUh
tlBkPELN0TY5WQMzG87+9Oaebk/ZYVtUiztnFGd0ULuC3JUS4b3/zx7vpT6a6ksM
DwCPtFB3cCm5Q9oxWORho0ut2sntJlDll9LMFam3cmySuoDVUGWUa1Zu3mjkotm8
58RoheQHZ6dBp+95AFKhW2u8ug6cZ1yBclfTy3zRksR8f8tQofD6ORdMorKhbOaO
ZzEd/ul/nfj+Lc2xi+YbFbTEvL/jtc43j/sWI7nIzYxz/kmA2wOyMooOIsbDFaTI
PxJKQryaEl1BK44Z7d8nmstAA6VsCDJzRETEdG6S1+8pQ6G6Kafzl4XvcSBmovFD
mz3t2mkCtvGnCFIXFvY3LnILEROoojp5IuUQEp+kR/Ln4lQKfuCaQIs6C0HpbB1j
or4Qs3UQjjplh8HZb6bpbqFg/qrc9GnxWvZ5OZ2Hbz0ukZAo0R3ukF4e+mDI+0Dt
jZug89NWiEPk4WP6WVKcU8JnvASkNWR2PoXrhFLGpD0p2ltlgmKNMtftoCjxcdZt
Sp/HQ8bsEmuesXwyG+VMUxr/z/4/HbdkkBjJl85yoYwX4xH37eOwaIcU3QLW/Ke8
fKWYC3Sz9irvCnR9g8T+K3900iGsJCrduzaBIzCFUgepZMaD90gKse0tuCBglWhP
nQ9ghSOSecH7ffEKp9CnVw4nDv6L0Hi5id1lKKxtI6Iobawdv0xJlmtA9YOaf2Sg
9Vd3SqglUDcCCWREuan2X5yfIZa0xWcpAVtmLQ4Zg4WvursSoX18zbAfptWg/ORN
eBxg77KVIFvIdtlbEbd33BIiC9O/PZZJPE3DesH8V3bNdZ3UOCnLilcyzMBo5X7V
7BmIzeS/uBCgo6iaih3VI7BjFs9qZn2H2llnus4GyvP/outSSYAoL6p57oRMzRz9
3PipuFBma1q1cXiiR+0TuW/v5sh+GaSmWGyetJAWzkYn+saweNZ685BKtdTWu3UH
kAEO3f+OWbBwa6O41rAll+GxlEVq1Nzehp7Cr6ICuXXzNycqct6RviVmucf6kfxV
F58Pogkb+Wpmjnt52d0wMcXeY00LQ7cy0CCP0WgkITLvOZFPJq/cwcDXBMo7FWpV
Y4Uv/6Miv+BDTs2M4sBP64BA5GnJm5SN5PdYE9YDJ4XtgZgXDzUb82/r62OyTL8e
UImmV0PH2lws8isp3gQGt5/QbH+jB5w5YGKlamhUfRi3UBmTdsCY8WLcHi1Iymnl
o9LTY161tO2R6TBdBwNea0LN9/dmRQHk9WaJU0Dy1Gr7En6ksj5i4grToDO0V5Ov
BFecRejAJ19yHXkbT1v91Y9H7N9Zd9eJt6VvyW0wx4RSPZT3+ChIbV6+ToMIu4k0
S7KaD+ulFwKaxsgu7Ys1o/J6c9mD1FLE8eBskwk/+taqrjBN9A9y0Lztght71TGx
zBCoMz33T+ZF2Wruag3h1QQlUgxctNpozgWRhp4+40q1vWKG4ousKn/vgDifNd80
yN5NHebfd4GV7YPQz5tMTe8SOWZj2C1+L+RYE5J1yI7X5xYKGBcS1rzTyshLMMGI
EfSPcL7OtVok6z0Hgefh+LfzeVnULIzos3yMzPtlq2lNPcngprbC2ugbcZUS59tU
Snu4SbN3f1hoHzfoSoK3RD8fegsTGFURY3uLr6VDXargOUJ+eKN8MCKXQOF1NBO+
rXpKjpUamZWfDS7kRjf+nO7PGjVb4ZSarz7VGn5EBV5YRt9bMkAODYL6Y/ay3Im1
cR+QluilxHTCkSVKHlBQv/zC0VifdSnXvpX/Ifow163PiOZR/sQ2L/3tgblwNGEA
FsAvzwPp/ai28Yn4zzQpLDTA4a+//xC7my3W0WxYjI8HVz6F6h87L9BFJkfJ+59V
tvE+eihR9bb6KL0s5j1NCgNA2YqHEjxkULqk4MLW+XNFA71JQyr2OihulKtaWc4k
usF2DemUVbPdHWuhoZWvX05viIb/eAq+Cbe0a2e6cSmTKQnOoqhNG+4021b5ycog
KRVw9NhkgUYq7pf3U6HIz4DIke3p8UTJ69ptPX8XowFQLpo5/FBvNpecsQu6AmOx
LHzleJ8aBjCPV2hrwyXeWxl8h7Bzl/qaStvSEix8vuH4WvNgBByylUVwXxkIXuB2
QyI0wdEmSFWOTH2w/vrrdAb+ApdhqZSgmw4FoGtW6DkAAjI0x3Ge+kRagMCGMBR4
PuyHCcQ1KyLU/EYf99Kufbw+NtdNeU7OQi2aM/UTP5JPTUdGd35tqqo1ssR/q3co
xsNrW0fkv2VAAW7/h8BNj0c3RsEpY5NWT6eMYDgchRSWEf8HwiuKrJik5Zhi29E0
OAP6+W4GiYExiziKMpwMTd2M4EBMYEeKeC2PfsQ1ovaT9W/r5qYBScPF++5uIOUI
aXFiLTcLC5mldEeqpefOLb1NqygF3dPVcJPUqD8ymZ9EIFfVBne5shRftFZRkG8P
4Shc3vkXSPTl/4aUmuDTV1tH2JT2HUpNWy0zzXOwV52/uqrcEvKa5uewsrTby4FB
y5w3tds26vfXjO4tI1+En/9A1h6ADeE3/BiAUD8QJVob1LTAhlbbUTTOSXc1BK3L
fgNkqpoSJY1Wva6HKdSVNxElvEnsx4y+F8bh77tTUIR1ioAK78BynjIDfICmwLQm
/kYS4BMdDaQCzmkH6zmF9txn849j7hcakY8q3bWXGLUH8yrxK5l2Zy1aApN4Uee5
OJZm1l4Vd0bSaorPxwMPfAsSHn/FfTfcD6GX2ArVwA+ku7uxjOn082mNSh4yOd9X
v/pDO7IUtYvLSvyXtmiJz9Juc4lfJey5qFhnWpFbbBI8NMe/mEOAwpTzA5eV7JHP
jxeCpzk1EJsGqhsb4TAneywWruYVj9Ps6XZvXfYRjPqFQoZ+PEvA1TKD+axy9Nmp
+LMWsiSLoxIYyNH9gT5kzcO9xwudEl1WQeUtXx9l5F2iZd0t+l7VOxy9w1GAJkaa
CbuQCdOcrtHJvsOpTjH0l5Iy9q0fsgnTcvmNjyN6TzGvzZ5dKk5P7GRDJ//gX0st
zPDOSvOctuUyF0YEDmdYqhHCgCWTI69nAApHXCG9+z7Zh4iKCjtiglVsP4Lk0JTa
cO3W9Yi0Ye/OgRE1e8CSzi1FEqz9TZbye6/PALY6YAPSZHywF6tT5iW5zFFn7/KE
Ylw+ZRhzCvC+mF/Yz/5/a3nEbG996vJhEH0Zf12rstXEUHDVtGSdurSqCHmnQ9W8
upbGgC8wmIKqqJqmGaHwwGxxv2K0SeYwAQcwzF6LzWQ8Z1bjezZje/ar5+r46JQ1
CyIWw7W7uyjiJIg3/gmoIJ7NbKOPuA49P+NdfUQDN8RpNcnbwTtb8bzbPt6ed3pF
5PpPshdUlJuFVv7ocR24Meyl2CTKGHZJ9agiMEjlpROGeDOunHjYIqveJEHgvPST
FGeJ1QVuJVyBmBUCIXFlcU+8BVR2qsgtgt8IlczTrD0fNOXYkJKbsibFXh5m8UtZ
3UTN+QXHaFsaZngQEPRz7BJeXzrVdnNS0tMNT6uwSURTEmMZ6427pQPPwDqAT8is
8oe8jOiKfTxzJDRezL6ZnhHEC9mY4KqyIbXdrHj6bFsHKx2VZn34wcTqDy3h/jq4
xJA4tW1LCyYhWWDuYobG4qFceW+XlMXGAhgzDX+Ph9P2bI1yFBvaR9vjoc7eWHBE
pkU75O+CTAl1JRCHw3UaJxOjg92Sg0PndxYU+v1tyvfIOMNJjumkqVYqx3Ol6JSi
q1swibynYvVKz8qANdvg/+m9L5wxeRETbCXHlpg+tNguVouUYQLKZXf+IifeU3ee
kd4dXLFcLd9BNM1KNIuSgvObNISEJusts+amDi0xJUSWkwolKkUP31wYbA/6oDG6
PlkFQhoTuoIq11tBX4x9U+UP+35EWmbB/U14cCR3/ID5h6xOeJJClkFoWrlWexfM
uDfMv+2T0uNr3grQDLV0M7KwIZ7hCWnp6wZCRtUmyZC5skANn9mEy7qchIahlSDD
Odh6CjHgjyrXeRItjy2S8EFvQa0DXf9gxaqpjpA1dmd8vKmc1PUyy049c2d5+oqW
MMfY7KDN81N4u6DsJvAPeEP3tfp41DAv72Cha9XtDlp7e1wLNVFWVpJF+z9rwYtV
lD2E+BDMD4CDpEvIwoTjBgCmnbdGIu+7D2KRfGvgtAyxkjux8NPJijIkNBMFYlEy
lkNWfOTDT0bPUBNqnGjzcFF2svu+g6W5JK9rxDC6MoNbLMKZ5cFtdDBGXA/OiCtR
5LSepW+82uudr4rFmepHHTv2aHutDiyT2sTr98I/hM+bj3/4JR9fKn3qnkT5zH1v
/vQQsjH+CQyX1I8zMGhSyfiSttJNf490nu/HH/i3z+ChaE++cNlztVvUi+qfiiqJ
TG0nZRdBlN3xNhVI86dFXMQvpkXK8g14DUFobF9crFcbbSfapLVNIT6akX59bhFY
6qFip6HGDQmjeq5G0xPnGjiZdhrAM0VqOtqh2I/30b137lpAtjXXwOOmehNEL2hX
eLK+QsWiAab3liLZDTo3Z5bQfYcuiDFc6009iFybolEvu7AuYBY++X0qF7Q2hRX7
s1ADBD8SVuYzDrBuFA602/95INSWBPnamaCDi1fCWkEo6yNfzdfN1Jb6+UmjHRqG
iHoB5tDOZkxjI3e5OPd/atMDo2M1n0yncM0jBP0yMY1lP9teiYffLMQmrwh3cT3E
n3+CBZAL7I/VQ+VRJOZnMjF7ZODzIteptzrmQqbaGOE8OZU6kBegFJcz8byjDlfs
tVx5jWeTiE5iUsqQPKciiqJvWz/o8TfaHRnWXqBMQiaKL/pePAae2xhs2oAE2acJ
V/RL6iyYBd0caYXOO7bZQ/1IXvhfsyo6yrPJv5V0GkgVxnNaj0/sOWckrFa4C3Ix
xLKGGeCkEaR8atKu3q5u7sMtkFUreyfXcofCvH7nXrkrpBxhSlZuLwD9GIal5YTq
Nieqbm8eAmC7CqXqp+m8ZBQ15YOF8vqVgqbLiJe6ucVpm/JzCgAatVuR/XdLXbLB
r923P1Jgtmuo+aUUIgfosVgsFqoBChNEv/x4ALJaFlFxsfwjMAtH4CY/pE/SPcR/
hviuuVqOn2o9TjLCK2KCo+aGdOZhAY+LnLaDDSrh6iVNHgJhvYQ9095siFBVniY7
A6Ugj3sc05jyoMUkR77lAmalDopFjR2NoRKJVkgd1w5t6tITNoo6lsWtMK14Iai/
v9ThwKVnyU+1I94NwMdQE465gMo9rR10gdXzf0O8EDc8WNP0nbUb+DOvh3mls/U5
WARq43Zt8Vxl+K19ZQyZhLfySv95isRsFqk3bI3+zNS4ScddWWuQq7ycgj7JIGxR
0G7JvdVPl5bEFoN9JlzEWQ/TlzI37gogHVbAeJYeGAUYdrwYDxMl/TlSK03YJudG
CENw0Irkiw+UgvvbiLdIyu6vGtZ60yaX/6/DGXG1Pf1a9oYamt2NwsbsA8IYwJ/u
WdCqMUAInI5S/K7pDadR8gUNnjB5wj/pHXzN19YFzwszrj6Q3m87c28z9WStTPuN
P7oDc/FePH3QCHoyzkEkEZT5+U2JFYpTg1mswtxjoQxRmQjIyhhtqgDZfNMMMixg
Mn9u/pS0BsaWCV1PcAHfLbTp99ZvZ/XARaq78Jkzy8uYTgq7e9U7U9Syy/UQQtbl
wg1UQO+tMN4LXPWaHbGhYA190BYKmr5GtF+5jb4XnAtlAoFFQFtlpCx/SJoTl2lq
KhT3sqhcp04coVxSYVxuvMjWe+gPm17eixQnDkkOXR+aWzEBmxSukRFlAKtctX+K
OVCtujM5T3Xk0s9NDkQVR/gX1mgFNQp1ipdEkGxnpbchWdb5KoyeIhPfrRw7t7tW
75WWaY+oEfNLb+SXZngjTNj9XqMgJDjxW+i/ZJT4g1uintM80ctXL00dmNIyDS0y
8LFCfu55k8DU9yPtLVYhn7Ugnaaekblw5GrzxuGHOZpXn9XN09A2Rc6oahYcItP1
UwwzpHuGO7eUC/R+qWRyRoTb8ZbPn0r2OSqz4dZ1QLGlvj4BCN3W8xKD6ud/6x4t
WGYNlcELJurvKEfHnkRz8lzjjI8InqgNIAgcdzcYHPCfLLM5fInwn8bCfGGiy3tv
lunuI9rrzJFFBaiibm6kNzFWBOhLATw3d9YMJ2eIr9KxAE2ZcCka+0epJz18PLn/
QpbIz/dX49j7trjN2r9xT0IKwQ4pm3ixIgC90DU37Ii0MmnK7z2ZccnTFmlbStty
jNTOJUigqyf5lE56ATYbib9ctVyNXrqYg9go4BZObQNvZMtiX1cGm+LqPqpfqDWh
n/C8Tt/gQIRC/Z6kjzOHSug/gJL2T1Uaixe9NyY8AwOvJQiwM1TFA4lR+6sNtMjy
iL2PhnQsnD8ZlnP70s44ypzoDm3H+H6E4/n9WjINV7IPWJiFw5XI52ufK+xq0R6Z
K9/J4VstVQYrj2Bwgk32NSvNJ2dIVDrfN9GSrqth3mqVxGZInSK4rdDIIQUxzxuz
LgGeD4acU/xRM6WjGEmPL/QgFZ3B37rIT1Xyb39BgZBx4HwkNEEwRYkQWpSy0OpR
fjBb5H4V4HqGi33Zdb7I9aQbr33eG2oDT/V5YC2aOzsghIocIPEM7VeDw+PjQq7a
dNdcBrsGCJLug+jr2+aY+r1aOo1Efr7Iu6btieYb/PeA9IYTjhMpY0bXlyBkgBuD
ZHZiRe+XC3SFw+nzgO4F1IcqkxhII8VeX8q2KRcZoE0AJdSF9YaQVr+EWl1O1Tpu
rBvNFOnYGcSHcChdOswsv+JL0ACnCeM78XFbIvM2Gd7qbs3knjwaUn6J+luzfxZO
vJuKu7IN5uf6scdqMa9HjTD9XRk7U95iuLwVZq6EqwbXYaiJAlNr4EaEn6hoOacE
Tozxusqst2bQJEizdeIs/K/sMyDTlkUQZ+xuH6jVPjJc6R84b9+F0I3EZjausePT
R4NzocD8eIDkRNqh8BmAOs7EquvH/5J97J8hwD/5HDnY7qgFNk5rn/r3HUlX08gV
iKOrbNnR3f7d+JZArjncNLuV7wvda1s4e4VnIdW8/F6ZT2QFtholpa7UAYgxePjs
ah3O0/UDL9UM5g/3vK3ZIfhHIar0SkkkzsAgCavbj1m0S1I4vV+jxgGvHew0vHug
khIZi5D9wLFafBxzirzEbgCMs+Ui6Iaqvho6HvD6sdGUUc4Jg3uxoczLUUS3aMI0
WBEa4cJZ5spcu+ETgySo5V1xu/ujwnJYR/1V1fiQR29GyKUKRutkD7u6tru98Id9
UiLQaNx+texKKXqHebzT8v7F//UqwYip0hxTHmmgDs3yz0STSvgbqjsBmaONNKGa
22sR8YsxlquD7skHmiBI9aF2dxCXYDJWCW2t+0R7MPG1L4XCE4wkgOXFEK3i0RY8
WEhIDRI5XPDq7b93QZ5PJ8rzoL/Oorpjac4InoeQqEO2JAcknT9kCPOM0g2PEM5E
o3q1wS22II5g3mQmaLJchE9lbUDPeVivDumA3G34zlO8dIA3Mn7fn/GV5VLjbZdZ
1Wkoe3EklzY1Dt2AeHa0o7bLzHM8Y7ay1aDKHPHHPS4cqvNgsij7m6aTSN1TijM+
vB73m5+zwbJQYwglU9kaOT7qJZtPxPpyXGja00jbDH3r4mkU0QF7X/3K37S5T520
54PfPBZKBY/MtuJeP5vC0e+fN6GEvx1EEb/FD+OXjY1Fnij9lHLkoevIBf/t8EnW
eNWBQ6uM7AGUizaKd+PDhb6Gjhd/KG8nPtXzsWtuXArwf0mGZFWkBMcKpdIsqLmd
oQVSCln1oTcS+VgyvxkcPXsT7VSn9armaU4/mOcA1uP6k+8gdwTnWfAt+VYSGXyx
JQEheB1zk4KVU2vptFEvDS7JXI/AEIx7gOMyvGcgzpStUZlCxPIRKYJFmCTRbxGI
6QJJm0Duneo8bF6kWtzNQxw63c7l/fT4qmxtMdtyCdHztnJTRCYSA5/wXoJWWF5H
65nCu0SiL6rWjNfRctjx3kmYtMYEcuSUnyqSOYmuA2QGIvXaMyjqviJXhtFQgo+X
d/FviVYiexZAASB6VQs9ezz6bb8x1j8HwqXVQHuX6h6emdIFYtwqRWuJXsVfJs1e
jFpPImbvtwx+Z8odYL4GowVYgJB+qAzKRNAbmIrrg/D4+WIDhcr2jF4YPXNC9H1I
Qi3Sb3f95GrinG4GSaumoENUd4NnKghJkzleqrDnOxHJPPUg84XZUk2pKo/asIa6
sbfev7yIrvBKJfBe5RAc4IgFDA27LODxGA82f9SJai1uHxMFmtLg/WRQ+KU8Ib80
qh9jthSpBMxSUzrx/+sbHVc4z2dXLGte8X3YRHhC7dmQOpEJMvUX3Wl7Lsucm99Z
bToRxw09ZnXXstdks+ao4QzFZDN/3c4tq6bqBNrd9ziFlJQ0gvJ0XsE/yOz+u92q
LZnWWJUMkzNW0tZ/pcDx5mO0ymyERKB0RDLYgLZq0Zf7uAY9GEy+vgLe+2Ls/Miw
YmLCm9YFc3PPb0q3sT8WVSh33Ep6LCY0OPUyAZyhwOhHtMKX1L8fJD5qmM5eF1Lp
vf61jWMNyTpGW7rsWUCgUjZoF/0h2XOW3mPM16TLQJUgEZhF+LFErnpL2jKjK/2R
sKBmSXVBIRBCKR4WwjWkFEPo/YK8iEvUVVO3EFtSDPDOR9kZjdU+jDF5FZPmDosJ
JSptfJHtDZi7PwsTXzAw2vhpSUMXhBNP6Gkopwh4DteCyglB+32isDukXEEkbhPw
ugGpvMA9VZCDS5Uk6K8CttkeP/NigSjIu21BQvvorPo6MDLoA0vVyqGGqfkORIvs
6B/MSb+XEPXrpz7RDWXPcMKsZSN+e78XhRuIbmx9vSXIr/hQlLnwOst3kX7E+doX
4d8vorLxBEUqrhpcHxml7pXlImeprm/Oj2Nn5gAIF4t9jOy+0+r0ceEEibLBXfr1
XRr7ntGUCBIOZudzOsHi1/dNhARwsOHpXjrvioevcVTEwGT5fNykYJYBTNQ/Ahi/
tFwTaJ9grDGFFukfPWLoyP5PiIuPNIgibAUptk931hL36GcbtKF4uWGAxrx02Dtw
OH/AbRYaceL3MFh+6kOnKST8N9//SuNxwXG9tkEvbST4zgr6q5cH97IqOPnW9SE1
gGPRFlnuN4YOosXUIAG2RnjP+gWIykaqTYdiOhahNyguPeEQJwlZFPf8+idxyIVP
CwLAkTtzDcxveY72xYy5dPgB+P45IX0T6v22OeH7ALU/mHVxr5sdIl0rMGTFsBOC
Lg3G75p8wzsGyEgGLb1vethxlkPk9BAO8I523duKzzacryS/o5ZArQt46ukzRP6K
PmIiZ9rmDnv9g3dz83SIRAz67UjE6kVedhrWkY3HlyRKGw1dqRbFRWc2W+MXdy9x
8q/XMr4Lg2eWzdl0jBCDYjc54cowMjqpn4b6/NVb27kyVtYP3NW6EuJDV5PRyxX7
WaZr9S3hrk2gaoUAIhmnPSf3dGxE8Bk6NUxzllLbnGDUwBb2fDI71FNuruzPobjo
QsS2U5rkapHAUSLQ/n/MsNuGLrHB1jzhxrOePxUfyVN2C96wlqtDczX1k3mdpyl5
kTqjUU+Fa6+maIr0an4JU60+PXPSpKWc3njWHMrdKGM6QiNE0bHFkwFSF8dzlam7
8qTdqG7KJNEvFPShdnbnvgm0arVuA0zpGVvAqjJ/vxImaJ3xDXB1lcaoG4xRvt8o
3MUrqvSOFN2Q9QChoWGZpldzEABUGGrJnlLDalEFZWFwR7xR7gEFhkQ6DZS+mOlL
fjxZhOzGTWbjaUbnoX34wZ1l7spb9fybBojzXqJDbLLppeN5Qwd5ufdmDEhCWkDh
f+o9FMIBHRyeSMgIB0yyQ7QiTSUVGEbnLSAuqxXegpn9wsd9wtmo1NyXHiHrVOSy
0s3BJJw4qWDho2O3mgDxmObqKtt8JhIVmKWv6fsY9mvDhj12Fl02/C8xQLAftzhQ
NMrTPXvh6Pv7jC00AGBUiRQgGqwQ+VziwdeKx07wy0xhnKMLr71xfwmcYXYYYIcV
nyeau0WwWnZv6gOjQtblloo8pz1/lcA0Kg0uqG/22Jls4d5hw0F5B8rTtWgq6+JW
TVuqiFQGiM8x+qXfrRzrVZLa8F9SRhomQp/63M2A8a16tHVTEUExun7fuHJGaC32
byg6X32PX0Eps9BBxGknYM+T5H8mrvQM7e0V5g1GRG/j9qYc6e6QagUokspIG5Gq
/m+JYip3CTLKfD09rqoR5cNom1KDCdaGbUBngz0inGU6lgKmkfnkd0L6gvbEkRCl
2WeKbq5M515+4xupqSEAZELTAFAKhuV0Dj8rRl3mpFAtPToLH0oQX2Aai8J9L+gi
pNRfX+kJ3LLaB6C7UwtSg5YYRCeG5+qrPjUmfMT9o3iFaG3v4I9hNvUaBeuxptMM
V5c0fq8yAckEoYdtq/ULg9hKCw856L6caAtkvl9I3l9+9nKze2PmPj121L9P5hLo
/bXV95hXr8b8+h6XKtnr+Huoqwor4FCQHjBfbfKDD+IP6+ADQQtQ1NxkP8ro1w7D
Hhp/hmUvicxszA6Rg+Wp41lBlzuAJwqUkys+8RUEyCcttzLikRkwMp6FFjPm7ID6
RZpDYyudr86znZoXUFv/A+0EMPF6b43S+20c/RVIzdZsl8zQ1sTo1E8HpOSKoAPr
knPYMUSjyqKhN1WtL2JieFc1KJetq0o96K5ATzeUzeC45ciYXUCOCsCFk5954nTn
NZXatyTLkrkEfZbT9KucgXV3KrHG1URlULk9ViX2Kai1DYffRW1p0Jkp0h5bGvej
cRtPUchoCvaoNcZrk9MmBR/wJZHAwkdPULiS5M7N9O2lg0dHjiJScpCFmdianNqY
LNhqAbU+I8o8udc/KBwOkcIl+4pyKZRzM85p2h8DDWZ+5i/c+Jb3lCU2mrin+ptG
HmwYrkpGz13FUgXDkwaj7CAS+TmUicwEonpzWNHjWhrDU6zqZXRqWn1thkGemaL1
WVKM3EkuySxQ55YYyi0EK9R7t5cw/9vcTiVbfz3ktGeNRqhKzE+9w+7ekW9+R35P
4Yw67YSwUOsUqdCKa3mHnHFcQ098YbyLqPAv7LKUBqMkfQk99sinpZkGwfFG5lxn
qTZhW2eyQ9cQXAxJb922UzTMBoxl5CNQiFwpj/vNoC/28L8ilk6gp7vAEoQicInN
2a5pkeZ+gPogLrBy/LZOJq/1xdENqQNlYqAwQ8YNFKexq5uhvAHTzO8LrOpf2LM+
H45PyRsvYysvXFfhP+b84k2jmHUIL2vd8eu6NS30JAuwHoscYH/So02AJ17IIXRW
iu92l+XIJB8XnMyZLT63UOTepoMwm7LSYDxwPF1iH9iSg4sDRDlgpOcIjqYJH9Wi
kZY6NX32lsVrP6PKt6sOmbY1c8miE45T+LycvtshZO5yRWR1iZX5mDHizWhx7IL9
AdTpGkoTJ6KGCMyRxmbbpE2ldKs3Fa1fyaFYJTzP1mPSsMqjw02tVjXP6SBGjOn7
Phjz4mafx6DG6Az7lYDwqGAr8g2rq2BS3J1P6ICR663JP9fDnkniTZVbru0jHBIn
Z7w+fq7wAD0MZfpJYLlkvkvgxQ+fVBiUuq6XIM59644ZocIfkGRCPkzv3g7fsITK
y4GRSdhyWGKctqNMNElAyZTOW9Oa8PoNC3VYJeMe30p4bIiwajM3Zyq9QFu2W0RP
GGmkKMpn3Pjq57WUPeJ/wMwSW7h1gIL0yLE18MDq84wozgdGTtrOd9Twf3Q3KUc9
UF1XvGHQ7rPt2qjJyPWZPjkUVd9onYPzt5GpbQnvFYke7hYaoCSKvg6hp76ObatI
QHY2+RO/Zohdun+CJR3zoV/4EkikGhuS0ScRvTO0DvTlIOYvKSjNErTfWX8aJoSQ
KPZvhGkX7rcRRXCfGDGc6YIruOa9bkx4Z7kW29ldL0tTb1ehwr5U/18oSwhz+VKe
0IWof7gRAdUzrKK11Y1dtA1Jo0CsU4w7tB24F03lCPHmiClKo8ydPeVn/P6ZKFRV
pZwICekMvkcHSubYXTJxeKQNwxmXH6DWwdyaJaaq5CbGL1/uIHHCAXNTpRAwLV8s
eLQafGtg13Q2ka02+24zqszsrhIA/oFKMVnXZkbQToF/MSCgIY35HbYlGHKWBoVL
7cmnSejJPntiR1SGzdbHiPZTKFqBvd01eBxubF8R4jnX3PqnyHO8jvkEQhgnl9r1
Ugaos+zWGuw1t62bsepruQ0OqXkE6dtaCMjvDz1SysmD2Hrc2JstAqY762sC5ydd
i0U170Avb7AvIYawp6Hdtq+Hj0CnHpfNKNeL7v1mZGetzniBQ5V40Qr7WrfNBTFA
Dc/1beT/XUe7wE+OMBgfotiBlhuTankyvg1Ye0+K0yfrxFd9ZvuYY9YjEtr6TeIT
RpwRINdj/dzjzQfVk4Q4qTuSxInd6SRaPGGAUhVvmu5cv6nNNEb4f0tnwQhDz8v7
yByrfdMLDMMZ6wvtxoLgGkq4YA3JaPlUBZJcg6xAdaqAhewT6WLB314RigYS02te
XtqwOGwA53yWADPGft/VRxZR2i2JteSWXTW9RWmJVO1XSsaHBKijdgOsk1/KzojN
iU2ufT1TVN6MoXgIwp/eGW6+zl9uN+8TohccDdOoI2JS1BtKLyo0hMliT+QUcIcq
Yzy4apUna3q/nnBUzN11e7aPZ+xEu379jJLsf65nxuyytPSIwi+7pluVSYIIV4u7
UnWtTaS3RQvdH+taG2lAlgRxdEvIu7x7DVta15yZiloljeQSfMBzFwYe9vcuCVGS
ghr4B29BYaFPE5qOcFWLPYqG2VJ6OCyWGSQI1KgmJhOMDPCTFArfUK78MO9eotDz
IesFlUvfZM88gkJbBxgQ78/xNe5wtGW3EaE9EkqNJYyFf+wLUh0l3AjQipLnvA0r
K/VjiMR84jiEGY1huTMrzRFW2qi6zbauDKEuQg9q9zOZTAOUG+0KWMTmBZFQdExr
tItUxMmMx2IKYvWiDcH6sgUwtyb6CApAm3jtLAzTW2cLUa7tjO+5bW8mRc64gXpc
IbnuhYCqEbzZroRs8TDZsbFXHMdDxT3K+cIdON6aHc83hQavk0Eccv2eBSukauLl
rfvYFOfsQ3+e1mvBeWjGlX/DfIcxPHg/lPdn11TyGjePj+UeerDiTmH3fvbEZV+g
EKhy1ycCh+AlLaumUYmaaZ3ZIVg0z1RqmSgL+Zk0lvm7KXnMjsrdpnYzCVePT7+u
Vr8mOmpbPekbChsZdTOhZL7Y+BFmCt5X4G+IlSglDMkXSmU0yp4yMHm83ZlaAfEG
/QppbIDBaLrH/hJL2bsZRmfWUE/72TI7JEp9f8p7MsByqTK484dcV+QN7y36MLYP
QKTCZLXaZMbtTE5X/tYIChXZq7Dnd9+9kBVakw1Cx8EWP5v7pZ0eOjfJ5ECxcXBo
GMXa6hHt9v5vQANBWWBSwqKEsS15sgsBbylobmoo+L7ceC7AUboLt73kZAwoxief
WecpzJLNGVPltpQikPK686rhKPC7Zl5wyyghxPrBSoiv7yy0s7Uo4V6hPTDOVEu4
gS3Bi6PznzdAPD2gdQCc1Bg1lyiUFOoTe5jYRII2QybvwG4eFLfClg8R7fPkRtUF
MrFNQl2mt1TSZbOot2R+qQgl2qXAB3HLsXkKkmY9Bn78Gm77H+7R5BTxmMIM2TQJ
VrED9Hl4zZUhC2ynelKM3JRBej4ymms7lslxwKeA7wawMJPNxsjbN1rCXIiF4t3K
kOSkB/Qvmcqb3j1xLEo14S8HjZX7MtmmT+0qv86aWGSqqX8tHuzCXPP4Ki0I8hoO
8+zkg182c0CDVYQohswFFrCwfqUEZpsaVYU23NZsPXrdQhiGYa4ddT/S/Z2dQYg6
sODxkAoABZyJFIUEqgDYLowXQ1euvb5G+9AZ9t7cB2st+g9BFAZs8HZbcpK0DSOV
A4GGK7qGv2k39BDL9RSYjbEmN4VQ3nPu+//RcNGvdYljJmgbFajQSXeYEJSz5IAG
IwsB6gA5kzgCLnjC83K40Lei1/lWTbXN2lvRTO8QI4xkREq0gWOowvobt3d0xBaU
ZQJ4wZMXiDCsXS2QeFKRP6mAot278qIhDT7RSZwAUIsVEFOZMC9oQprVfaemBv/s
5aUUSAg9IXqTvLNl4QeQ+hUkJLogUL2CMFzAUvJzkoKyuK9sWm5yEbpPyNqAUPTE
3z8GniMxPNW7SZso7HNrv5Xdu79KSK1OAHWd6BWvCrf27gH6FmNJqAf7huSkXs2d
7xj9nzu9M7lN4G5HMSjciA3xArIg2aTD/Ar9iCMcYouvG/SGkdTMn/sCMfrCRUOp
uL+nfAbBv09eKhb8Kpmt1DmWHx7NAPeBqoc+FeNYPemDT9+8hTu72OPXoc7JFsfK
OMxyGopDqN1hl58CEuJe2hbrsfNg109E4OwC4y3GQm5pEpadUUwX6B3Xqmt2lpCD
VPh9X9SQfZHIEdQYbjU8dBTzvCF4SPGVHXZMPVYze0+DGziIXn9XE4VhtoSjekGy
D635vt1cOgJHLvuYuH0bNbo4Kvw0qgWHtCy313grTl9OwU9VTIJPTo6LyYwPWDKM
/RQjKgZ9XizPwiXTLZPx+zRIvgQdvXNn+beAdIeLZnrgD9eIY1yHTg0BpJ7CgONO
QJyDf1+Ciycj488RafzF+C/hr4i8czMvY24Ob1j6Gh7TysQv0flizSTqRhXbLDu9
MUFVTm5Grt8srcQxnZENsUpwwRB3aQlSzkt/gabHke9OnzrFwf8onY+McrqYwqIl
hbHOjK/nBfXYIi3F9I9BSOQyC/fdX2rBebjuaGCjSkHtEZg9RZcOyawEM2+ZHM8j
rBwqQJ/3vDSHSZQ5ERmvXP9txWdcZsw+n9B6ESuWDU3h/x3ZtXs/+cg40wz2JSza
9NAgQdCXr/kgLF/uVUUvgIk30XvAFU9Pzbx+aU37xWguF7TBSO6xR+aDaj5gyoh2
bEdUq4g2IZy4Uc2SFRlMm3Wd7haU/kSVm/8BHYqN1L/cznHm6ehCnnwzGnrSLBDA
9EhBLso+G1XGrmrozNuG3cvdXu3lTyJ0Sp92iHh0OuiVa0nAfy50OG9AZwc//JZW
5JbN3O7BlxpbfV9tkyhKQN6w7NwAO+i3PDVz6pCWirh874xuX3sX7hvhz8vPYpVm
SkTYM0CatCnupg/a5mQBQSuACsoWWrn6ii65KtbRYZkSDYDTBwLb5ASNlwim4sDZ
7Lae7RJ83CzVqv+Y7z+zCOgC5PpAM23SUQdFtm0qDr5UGtFqSSec5bFpy1eiK+HY
vrGQKXzP8XwFEH5tE/7ZlmSbNc0MXKPsAVWlkXVYHuHeLW4MmsYAK3hMSAG4K931
WxJ5pbcFdVTIs7R19VQpLOp9/+YFH+PjRrm4iKDOlkHX3CK/nubop2htsib1p5hw
RtnayzbJZscqO1d9GHQvSHqAI0cliR5Jtry8Pxu0IGNpY0tiQ4CdTjgS5dlslHrg
SzxZAPgB1QVWvZ8SH01LFlVFrHLs9Rlqjr+UCPC1/suDB9YMP/3yafKwfbEOdcOP
6XgpeAqM1+H6PTLkTh6ZIh/IobzeL5dglMG3i/+1wwWZw5Gf8WYTMDKHs4xdTYfN
zL/JbhZr2nVqrjq0ZPpTxFvgwUpKb6JPBoki7Qh5HYI8RnHZtdu5roOGHO78lID5
Ozkd6/5TFwcfP3IbbdHC+SczKEVWCB4xuuNGDWYDaZc5REFm1PMM0Pz2+RUKRRKQ
7aEbHF0VwAzKON5JR7h03D5RaSeQgYyPjP/H31fVef6s3ZfU8qnTi/5w30IHq9WI
qUU7YXgoktyu3iTRhnBnmhBq/bZAjT2awCevhfNSVcDNi2dwjQoXdjtDRTihDBPf
1ryUoZQa/J2MKTXOHDP4CefilMehBttZzDpTmcQSZXCXN3PDdctBQ4aZpOXFythn
oTIKyHHeCAuL7pEWaa8DhYc4rzm1FBwMYifirFKB5tXANI0eyWqjqA9M6Ri2Bkeq
1g1saXXpRt2KpECbk1d6Hwnm1T6RTm6BtXIgS3nCQG2JHAn0axs5UrCa5CMKXVqO
Fda8MIYP5L/CDvPcWr54kYeOdGrs5FaSV7+0qJSGPKpdCyk7J13Whb3/aSXD0tFN
6UR3NEsrJfHNIkFahNqKtkyRkL4UbFAuaTsQnOtXakQ61MyCeGL8vBAQRqaFNmBU
E39UxAlN1e6AAo/HPyiQUV6mBks5fDecbSSaRQEjik0t/ykyR2m+UEszk+PrbTrg
/ag50Y5FNagj3MVj3rMnzScdaXXYoMzZpYgUcRpOV2xcQJt+6rYzQAi09VcDgwUZ
D/HHX8rOYvV3hxxSRkc0TW19kA5RUsuyZ5ht/YzBharYdMrwqDj+kxGagxePcH99
piRp4Z5WVP5ItnX/hhq40FBd2playvi2o5nx3kYI88IXKil4obewJx+Z+ATBJbaA
4HVjl7L6pmUki+VwWkKCptbxGZRt4QK0x1fZ0A60RrV47wqacbMq7kZwZr9VNXKR
DLus9ZZCIXY3VQQHXBwOa+9y/zFK0LTW9HrLfgt4ZEgiLKrfGla8TzjIlq1BmlBB
ge3lITd8NK98ilHOjb/5ZB9/dbSSUMAoFZJdTJ0FcSxzRzjUzr8G/zS9DsCRSlyt
QjX1oImUGUPzfrwAqa5LPjtTHQ0C4fQMcz7g8ObdLKSE/sOcBtIYwRK3bylKoup3
pFku28kQ1eVkf2s58AxRVVeMB+M1kKQl2vHjXIfhsONyCiiCE3CsMpYX/E/CQRR3
HSMfY1yZiXMuvy/7bwOts8BCuKTKniXwZE4c5e4uWXes95KaizluokgDP0LCNM1j
jyJEsbfWGkHyjYXqwksr/gO0QkiqgIOvyyBE+JjcB4B5gx8zaov7jq2h6Dph//FD
YMPXvaEqhf3W71+qwwktEr6S+3kzvuW6Q4AqAnsisVeXSNj59bIpTtoUJQrw33gO
0qgCkqjwRYD7JP6xpCFIoITJrbscZaHK1IgJ1YKAvFoSo5fgZlf/MdsZBAHwlEQj
iZUJLxVCQ2FOLcYtZ+BVrrL5QygUI851IUljiZEevgKMeNDegaNo3IvC49nTQz7x
PUj+XsCSTTICp8bWoHolUgp3W9Kp64QvN8Sht7OH5WS9aRoj5N6jS81f6VPvD8zQ
PLaIrD27H1KYdohIapXNvsLUfLCFuCi1hUiZMSxfjWtKD1Vnt4GxZ6Y7+iR/G6QT
ajW58xfrhM1FSf0W6s5YB+H1o1p/Qh/S1KFti9IUiUdK4fsnrMl1dwiebm/xXhif
A3yKLnmtPi1GPMr1MYzctjB1KywIuDgazZVjee+9lJLOV8+5D3pi/WhWDDRwP9Dv
JAHK0IMq7j1RYbf42Mgq5rZmbE5SrYyvFcSn+MjmVcLVDPOYGkxMcg6jLce+yYlG
IUtwNWIbVcRlyMAX5IZwDB5kFYeISEIc6a9dPOiHRssHQYqbc+ugznHYNB5F+AZ7
zJU93f6B3Ekvm1d/MSW5R7JYPs54IopK8ixXXoY93J1U16nPcArwDY0k64immnjy
+1kCUWgnb2UTGeKnOMRUlz2ElfPnm5s1yBb345oUBoMoTIvxoR37VuKSR40x+U4M
cysKY5hPNn89EMA0b/m7H6FGaV869JGRugM5Cx/RcFCaQUNjwLy/8+ueOv/bqwu4
qYDC6SsfixTpLv3Cr72GWNrROAtfvb9FcUmUputSltQNtbNbg8TlOrHNpTuaqThk
svGNACQrKaGc+vkmbngqJz2Ag9mSnPcOd29I4xx2MiRjPw86KXrT+jLGouiRTguB
qH9CCbF5Z/dnayEuvmJDLQOBrveu+1nIzmbJXD25aMXyHMI5tdZ0vFIA9JKerV//
dvDoSe1+K/+CiL2thaX2Io5hXgs0OY9VE3jb+VYzuDo9qT+MoRqg8tFScQ8iuz/L
fXsU7h9AB8at2gm3qUqhtJ2xfx/zHEAXCc3rIsbqlR4duIIYEcqEf8AYHfgG2oWq
b6kXehvUWJATS2BNULCiplIc5FLtpkbbgPpWO7JLTTZBiXDNepRi7e7E+2aL6MkM
A6aYOG2FXxQtf8qIXifoL2LH0+A9k5EXBh7f+vVfTOu0vhczkmun480K41qHah7q
siE03pO8ZNZhYjvZyXY6ZRptBfRSaeQPR1Bb5MX0FSH6YR0LbPBanMh3CNbmVag4
hOUlalm+ii/tbLO5UuzG2Cl8ldiLwUjjq4xH/4mm0tc0iYOrvwDD14LwTCwymSww
WnEjLF+fbxdn7ZUdsSjwGloOVdxnY/II0+6D4SzInlwXfKzg3uVmo6/uAHHr/ewe
WvP8ZjpDMGjdOoTlVMimH2GVRLCwF5uP01FelGaZ1dbIqllVLLeZkVkjqXyozfVd
H6zjsWtwyxtwAMEadg0s4psf2ph/B4L4SzCc90oPbdZA0esEqhRLYWJinZq4a8sK
f0ZkQn+pMZwodpH8Buu4dxyvxCqZyci1VMoNBIxoGpLJYdd55Goj7++vsRh5L5PB
Ut++3VMZ68J/4pcL2YgCRPq8cjlTIdzCoEBENEpbW+5ndBGqSdmboSaBBEycb1XV
Zf9JUopjULp0UVgP1TTGDL/jZO+vGuTRAXrKeZhsRDcTmUIgSu8qIkotHaaPU4LM
YM9tZz1xJEAyjjbuRkY+Mk9Ax2BGWFRm9ansBocurPa15DVCd94k4fpXdpt7GUf2
lj4L80nIuSS+VCNMB46ramz5cTFMWcjHg1t0bMW43Ee/pBdH/Y3mX+n4Q+8aJNGE
zttLIwP0szoM8h1OcgKMQCYUxMV98VnbW7bgSY5mkgZEF4vBclduLNbIJTmzBym0
fWp+gWc3Vix36B83GTeh3KbPSF6bsHH8hPvqmhSyisIHGiS+wBb02Lz7yihnT5Oh
XAzolMo4ljZK47J1FboVrwye3khij0qsLC2va0NRYeJ/g+fTtjNHndeWesqol4Hk
OuW8nUR2PxC4dTwhLxeXbB2PCIoETOXK85igTPW9ImQzlUIIoZ6eOj0533ErjPa4
HrBRdpGdqKSgjMZyds24hk7khcRyEWH228r4+ZGdKYy3Bbk6T1WiAGixLdo47gBN
4XH5ZTCnJZuJFYSCjoKQYgWOlZrw6QQQzXK0ecTGJSJRC8vSHR/8P6FsW1UvQ4Cl
sHSxGzQRg/GvVbf35XaYFP82XTggsmruxbp5LYV0AcR1UMHeeGGcOgp3FnzongFr
x1ZC/Crg0o/LXntPjm/Cbe4p9OooY5neoEKBmE1SmWMF3n4GtWdmYcmU9V64WBp3
Eqrhdbcd711enA90EgrhalalbpwddH5uKoxfbNIG3oFQtMezVe7/g3J30pVTvidV
1tTJMpavH8xRuvuKQRaPOIbwxD2L3xXEtKrsoWbByL+WC8oJczDL/t9+Noh/pxhl
Hl8/DluA27PNcTbRrdztJljlKk8iaYP7FUqFCVdY2RQRSKhw2byeQ3z6aMhZ5wx6
RY/JnLW/jga9TZv5BewsfmOQbZeQwpXPTEs4Yh4CKgLHrWthrpuLD4RGVq0fOnAT
6FweyhLi8mt0FGpWFE/QvjzSrrSTKBAy15mZJK597tRQWOSRahqxZO6gCAcUs0yX
ZvgJGL/mqubKamL4wyqdX/QmJUTK7WraLsGfOYwlhg+Tl8ScZlvjcsqX6hQJni0N
H0zajT8RSHy37k/rGL+AeGD2xYRHBsk1LlAdhX0t/OpXYzircCbybMosNlwckHWk
VCinpzd2I9Np+eB3b2wXpiWxaP56P1kvfHntYNXohN2L25z9k88GWncJ+9sVP8f6
m1uiTOelhTKs2hjM0JAaMOe3GrmhvvjrC+7Udxvd74u6I2H7rhvz5IsYUN94kMq5
5flWwjOytpldL705yTzOSCTUBRvu5iNc7hvKMFXdxqJvEXsfAu03qAn6fP5tiEEA
IV4b+kAXcnxXLrFiBeY1I2JTr0NG+PGBSfpjKCXJNp3tWSwhcgrQCI7jJonl6+5d
EunY4TGulP2SMmK8zCWiNW3P55eQkp8DvNB6CJ4e/iRGA5ViKNEB76nLWUDGIULd
ka8VpcsUa6bhfDhUeU1GQomCz8Y+S7R7/Y7AnpAqTmFI1HUf81vTRFd1iMqAaHWg
AGsYHWAYFjR+/aJHqJBpYII+5HnhMHAESsJPunYAZQJ8SlMD5UVQ+WbzXnNFppEq
pdYTOg4/RYDvNATcJc19pfqfpvDH0lQFhy7XkJQ9hOh72Gutm8xL2EoiqYt3QClw
qC8LMnzf148/SXI5qqd/nsZu6s6UoXZh6+jMe0MhUPClQ2aacU3DNGRn8xZ8kHFu
9oH0ZklinkVqnWAmuuEFXzMg1ByjSDNecjmynkCxsUT9NFUdqvEX1H699BpD5BzU
oN6jY/RlZGtuGL1/TVgirDiMOAtvhBXzzoScAy5s76tKnKQ1i1cPSbs9U4yZ4sDP
9kGVwFo73+eGdcwUHRJDTsVfOZ6tUR7uCCHJ1frgorPKBWafDzOmBUKtiZLDoRcc
NDRelHGRxAgC1t9s+sUoX+6sFxdWAjVJ7CB+dYqu/zCCK195qUbnMOSQVvG7e1ZT
E5g7f6W0MpaKeQ6Ta2HGnY9u8uLcoeWboDhVQI2PaAgE7stC0q8r/UbgsRU2mWVA
0oYNQamAb7MItR/1jQmjDziacZZHHxUxc5MwEA3VyGwwrBSJT2+bJPwTW9wbdGQn
tNpP33EGKL6+qHXQ3JBTZtKzF9KJPUaeYQey1g28ftrLymJQD5kbcJQlaUPswCFZ
xeZqgPNkvG9q8d/+cZbIk0LDzw6iyu1ciZm99eaAw9CNOsFU0jbU5GfknFG6H7RL
geTpmIYLEGg4PqEdmZ5T1ADEQuYrJxY8tQZb3UZufy52LB9pMsYYQ/nggfRUcYGQ
jJIivd/bkR6NWrnfvExw1nlsP96nJ0y1giuT/UmwmvZua8iH8SsE40Yy+Ag/vT4y
/8RlUlruh53lSXAeMsmuAkkAUO5LkZopzViaxjoJ+VoBZYVjlnlRNtMQJs2tQY7p
7Qqm/00BaG9Psv1lirq03POMU6YjjYW75B+R8i+dM/fkYzmwOmTQaV0JT+IuGM+s
A+wjCE0XYKlrnnrXFeFN6oEX/sq3LJsBjw8dw+BctaYLOCFTOwWlAUjsGjy6fUQ4
EfvlDpdiEYCuJpjc3tq/L6C+PAPcva6viyIyNk87o7xAoHcHjIKMYaqj07VvJQuy
6p5IIJG5ThiAe2tpNv5oJhqXbxZH4tKc1SZwbFl9MjlJS15DkKO0vF21kg2ggYhX
IpTcVnOUxs5DYjJj0eDWYVP/QCxofGYg+Gs21Q3pT7MwdKz1qmypW9EDJyqZxRkR
xA0utIvAizjjR0EEdMgR+KsTvHgegLh2X7KYQrH+cN0TN3HVkh5punCEh5k2J2vw
loaO+M3fmbnMbhbdAljoAG9bQ3sV/HSw9yHg9UUmOclnSRWf7GNBnKDTo0AljOKb
M1Cwi00gUSTo/1XSrIFk0E173lnQZJxfIj0XoGpzgiOoIfezEVvqSXTxiatKoDje
6WcpSD+gCd6OqQxlSP8bAvg5vPUGo1MZxxeiHGSVE0ZXRQ5w4r147Qe1H2DFHfSa
UuJxesj1vALKhj3C0re5WXUqcfOoF2aoA4wyEOe/411YCk5I4U5eWVM0fvXG/SRc
FO1X6rlaw59W8bQ6xAJNmoYuhJfu+kZF8eSMzHej1B8RKkryu9lM5d/bsJrQ2Ds0
2p6g+aKFnx75rpe+xkbPUGVO362FXOvEj/X5CadzO+HvKTzopyKNYLB89kPPbouj
8rpSMqGW0BXoMBLMSNb60P+b0GY1hSYOvKnrdB/bQ9m3U098GJa+BUOBfFzrSliu
GERjheVj/pYSFNZEwxyg5sijqCrITudef+whXPTXJjERkQV7RyPERo/Yxu4LccVE
EBiz3Orn084vw3lzjxZPt2KH528rGq6rJm/uV/Aj4kx5lmnBBojuvAKgS/7EO6Yg
R4r3UFzZvP6FLl1h0vVB+Bzj3pxhjYBx21hVqWsfsMv45sqjkQO6Jzky4XpmOig0
KYSU5+IbdCt27y6PuXaroyUhC579xUteUzUMZJxd94L6+BidwUY8kQTdwfqcrbTk
j91Spbx1ZWJN0gjNmT50ghD7aOZcsNRI6vVzlC0KFETKcNV9wEw+r1fxT97eayHt
G2xLsynLXwR80l1EmFHKoIPA7jw9Z7J2Stb+I9+zQKNPSd/dGAfYtEZ762YmwukH
PJ8f56/K3Fo5vFgnObwsvQgCHgv8v+fIp9XmvAAKCXGZPc9MksF+BEt2MGJVzlsS
oxLq0xwrjmyBQFGAiwN8cJld2cRI/yQj/3Mp/f1n8+X93UJ3HkNki+t7FR/RTnu/
IFNW7x1cBzv+Wu9NZZXaBi33vDI/r19pVWnewtuFNtq+fEUdVw0oX8NBC0DfS2+3
3isC/yn9TF+IIqUVRWCpp3sUldYfoOdYyed55xvxXeOkP4NWJXMTQ35+FwSVjo68
XyuDgor7xkU7Cprp/vwRzcZ6pM/VYb3D0MdAbJQn3i9e9NCdBjZ3d59W3UjMjexa
b/Fmotv+hv9l46z99KPzdZLkGj2GI520QqXKxXwd7JUURSQEOaPgUORCV8M5FFqm
V0auINoePJAK3sjeqDqQFJ5hDb4i5UVGLSr6CHiM0ES4NFxMlU5pLKeRHPmChaci
+CQUlOtkcuLkWkSfmrrTGukRkzTwaVeGEPdVzTYD25vIdPQde3IR+yWuucuo4Phe
ufHQF7yfv6ETQWUySSDx9kHaF4AukW3guOzKBuqJQUR5Ds4/JE7x1ibJa4A/662Z
tv4yff7QkgDLqrvAS/jpLhgxnGLjN9wRf/6SNntk6yW3amZWqIqSqOMKs4qb6zjQ
tQMSQNhCmDJ5rzA7LenkVCXV4lzQNVgDypoHlsk3FViWMOWgqydLYMigldbjC+9E
U5AMg9KegZXDkdAERXnG/qpjh4GtXgZBH28iVm/tk/K4m3YC08vQHsdqamrTxZ4u
90NbHlvGPbj8J6MzrhmQuG0kbsZjQosolo1do/UrNG/QDGOGeJYFwZGYV8alADOd
XnlnTdIlfa5SOtSDZib/M0fdhFbmidYuEcTATH+pUHqro/Gbw428/H/Ltv6eETK1
cSXSuqhlvGssvaMTwZAcCG/Acf89raoWL7UFCIRTfkIlAuHnZQuCfvK+9BiRlZru
a0UlDfAV0A6yxLz7SXvakIgSkJxp5H6x6z4NOyO4SjDSf6gKq7p26vvbwNHTx2UN
g/o571w23PAdxYXJZdNW22dhEHdvqVEkdPAkHIBUvj8bu93v66uPRhvrc2s6c8MI
8QPSNMTApOPZXgc0ShwC+GQ7Jw10+87mONcxoN965zHW/dZrHJkbXz3AMH3IPqeS
8fKXqtJZ8rQlV9v6rxyZhzmHqSsKCiPb0wLlz4k6Hi7OXBE8VmMoSi7vt5qxGG9W
rIs5qoRShgdQhMGd2bIb31j8KIKgVcR0trKN86RyhCZsM+1E9lKFTHkrR4xPswYE
mr4WedGOGqmJtBIu3mTuuvobU9a4yIs5Xt7+nfFhL5FuKV+E84hLHnrqkum/HZY1
hHK1DDXqNjTz/hzPGk8PssgDILnvfQaKjEkfHUiZmAwC6r60O4op9x2p7CAwXyIO
2uUgF9tcSfcfkqm3Wsagy0kBQMueaj0xHQ3umfETSx3+3YiEDU6248xHBfajEL7x
RqolIfH3ArkRmR7mFV83mmhWhWRJnEFhOBMcDHEWN7C6TA5XtrQEYET01IARG57L
JG/bLWiawDrqVOJwif7kamhCVlQvFbgipDS5jTGdQfruF+ckrU2OQI4alNFcKs06
jIS/vC3K57StA9irDzd9E+OF5Ov5YUQIPXDYu48JHZY6w9P15NSLMQHBC4l6M2/d
H1PPF+wr0CGSJOAhPupkC8VgKMOF/70zaqrUD+uw46+UAlmeLLFyxLVR9wfMTHHe
BgalI/iVrumxvt1FG0X6DJXb6cvKebdRQEAe1ibTj7RpqDOf8XonaxzvM4mqgYz4
m/p5ycuiGthc0T1Bc8aAKztiaCH/temEUk4kXAtGcRAEIpp38frrrkOr+nsyfCh9
wLHsNTp7HMZJb8+HrXLysYSjzEybFwf/49G8uGzC8xqOCVI6YcEiNs1uJP69Taid
AmTKvQVvxyLQ/Tc6Rka+Si7wRAul4QhXIUPbmPkV5yEPOIqcRjQHg7uFjIB+t1Y5
DQMu0hKqN4DaDLLnV9euHIMfAiY679DkiQ6mBMSbY+3TLGfCYD7k5hktTize5I+w
AIEv9qgQ7WypRB3b3D377ISsYw24BqtnH/4yzkhzv0AhCopL5zegH8Nov81HF9G8
mKa4d0m5UUb/tm53MNbsfprEUugJgjXkgWDp4tVKuORx1/DppyhRGseXsxxGkExc
8QMJgfvFJ+20daegOrURG0lUSZIsnxYRmhh+ssT5LRdssL82i4B7OYRK5YYN6PSR
VgrQoybvAJxf6uG+ZI5F7cjNPxYHJPadJE+lzNDTdLnPbQYzrwQV9ZnmqPORTF0B
CDcdUNSb/bv/iqCtF7egSXaX8OOQu78Hj/TjFnoznl2TK2r8WX6X17EeSiamPzBY
LdBwDL9n+OEGmDn6BZrCoPjcO6vhFH28FmBQvfa7RZWFKZj4vGe+wB43vpIepze4
yeaxcRA3QjTw1rugMPrMHHs+PnkhV/HES05YMMicUfsSFctxbQB21MHUBRjlMo7m
OTostkodstb6PJ2gLziMIJppCEn5L2Sk2kudTSxuclkYtUbzy8J08JLfqaE6gK4O
g4WLK3iGueXV4CXAvuPxL8iieAFXs/IOsQYDcLKrmRNzcBUDl9K+evJiAttPTK60
wWX+KY1oVJhJWcsDcxGLN7/ODm9swKN6Dzl3nODtD9yx76Jf5T+CNy97EtMpy08o
pnRL67AEAHNLT4hzt4GHKvTnJ63R548DJGkTIx5zLzOG+BppjLQN4pGLLlNRI0Lz
9pAr6OWHLj8yCN3ep3kaybbvjkjIYQGaouiwUjPhDZCGvIw30/ApBp4JL9XYT1TD
2fG7m1guSwFnnd3YgvJkE27yUrmo9IJYawogVvfU0XZTX0Fek/TioEWPQAE1Mp8Q
UAQ1hKiKKbV1gidkcBSMQFd/C+2BfcwpkMSitbXeQQgxkRPm+3y+QtYhxFE3/ziu
foEcQQyKJ98WZzK7PJVADfQ7Tykhuab+vGOIpgOusohr60x7H37YgCaafphhPkys
jdnsQR3wRXG8gnlampQUrikIW0CtZsSvMGFJtL5DbFYr9FsW4qU4LN7+QXwblwnj
fMvIdlZoPQRYbYLchxoQRclrpnPSXNbwklLTfgXzJQ2zGkyu9hJxSDKIxt57Ubwm
+HJIc4eQGaod8BGhvk4dTbQKk+5b40haZkJln7DBiDrtcEmoQDhyD8qqp/MzaCvz
bdRAIawMs+fH8KXDtWShTIoFy0i1HrEFFd7Kw962d/yKCzoPP1d9siuPI14Y4Y0r
HKLd9sOOIaU4TvCEdwBjFRvbWOONtGCP/WBawfuNkaMp3nX8rinlkXr3wZjOz/NA
oUhY/qEwZvEnan9pzDyS3bEoU0SDtUV5mPdO+r4Ix9WOu9/WZL14GRFpj6FKeoLW
fwQluS8PtMRlt97s0Ym/NvXVyzArfbNXXoXhI26pHvoP8fgqf9eebhr5Cl7tNE6g
4+5ZHs2/ISeZu0XjWjGKu/BLdhg9zy7BC1WzXEWNAxBSvgaAnLHQcUUhf+vKnerS
BUCtWtNrwfImTV1Q5f3uubAk8MCqjKMaCjNFNJI4UYcZF8ZOLd1030NEc+5FmVhU
20wU1Acwi3+tqjtoI4fZIzfzOO/Se9mFAkWvREZbN4JsxDmicHZolKjQ8+K7e6tJ
ke2iv9NY9bU1i+d4+pod+9QOnhyzhAd2M5XhHwHAfjVIkMNHTmAaOvIT4epzoFl+
bTAS5B1F7RNiPy5eCyv5S6II+9+pt0NuqvSdw6ZTODxaiob2GRab5tQe/DYO77Jw
c2uScQonpTUO7A1BiCKNtyIkI3b7euI127pkp5gyQd5ngP5T4nTANAcz5OxJspC1
sG/WGqTCefOd+KykbUFy57WBxQUY1djgCKqI03uP99Jp19Y0XLT6/DbwV14JyUs6
x2G1oMLK5hbFE2bZhv80WgUy1IChsKLu0H1m3WRbC+z79vKDLo4CrMCqbU9haPM8
tn4QrPbFqyco5q5Fx3zDFEqLjhChTNGajZmlSMcm4meRbThOogyLrqMUmfGtgEJW
fUCx46t6R+nggT25cl13+T/8Y+UBkmEdW6Ch18D+J8DzQHINswau8oIm/w00Yg+l
0ZtzPly1qEvaNtooEKfbc9eOItZsWHUayzhIKlSRtfwasRC4q6urx9kcnAv7vRGK
62x/IxuRlkVJkoyrhgA07kc7L+yslA946c9z4wrVyEPB+sicUsXLR+iYOx+YQeZ+
Dwir0DIF0Yi+6ldaUooSdwWigqtp7q7yzUQSqWzyXrKhPbPIIfsH04+BhiyG1B8d
4pRpYzyVZJUS1Nm/x7GCsHYCwRAhFsc4MzDJzAjVUbcKBW3v+3HgTQziVaWH/6xr
R0jPGPr3MF3rJ6GecNhA+q53cszbvStbqcYznIJoWISHTsyCS+2Oa659wlZOKv6j
fWYtJltwCnjZdbm2eQJE2mw9tAfP05Qcz96YPxmtsheDiLZibERy7qEMT8oKwD6m
FI6TJVkchvCp3FPN0bn7wrAV8GesoHzHuJLZlrnaG3gosk/P3cGY/tCrp77oeJHe
8CnBE0HwU4525g1VoXhqLLXLDeNR7ykOFNF2Vzb24qpzoNcCElw3GwSX75dFlTZM
F+9j4lUML+/i+cxmH650Z3jVU10eFhtBJlUJuN1rB0lIWkkQQAjUXG3zcqB0eFEV
w+3LiJ76v9In+nglMoinUrKNKh/qmX8jrOKcxcUBouUjmFsHHe9bR778TmYzUDX4
qoXc1ROd1nhYTQogbH0vD3CTnk53V+JFUa/1x2AH045tQM81SM13J1GVt59PupyS
GYomlofr33TpBubYIWkq2IO579SExY7sCsclHBS/opjL3GeKd9iK8KV3iSKZyELz
ECcEIlFy/OmDmuIjMc/Q5t/FG0IM+hkzJbgQC5pCM22SQfKSP24P16BCmi70BetR
oDBbUqtkUI5DLBOd84NO055Qz4Gka4xouoabozAuDEGV4AvS3z1EnG7TWFCkSFl7
/fekN46+IJzfr5BefWrTMzN4N3NIYCYqblJ4E/B+077adkSJeOMCBkdFatdIcPYL
myjvimv7yhLhcJDF1O3WbUZsNsDrW73Cu/KpVenMfqKkvggCh7b8ws1/ZxieLw2D
MaDLdGaDe/t1TzWYEaV+UKNYU6vduuF62LYApGQRX0WukwBMLtp9LnACMkJIfdmB
jYG4Oa0zH6KmG+Ez4YuX1sTQW/Kq2/NvqsPLRtQRH7p+zGEFISj/aRxX/hXeJZdl
MJHbr5WgmN3TN+GXMk62NEdNHzryc86NLbiVZNQTBpqJgEiFYZDQ/BOpOdkovDSJ
BsBF+Oo9IvjxVfYVuHkHsxzWRSjP9NeQm3Dznh6YS1uTr9besU0fuwyWhgpJhqLp
Ykycrg9IcwfOPPR1FcYBlcZqJSCl8RbhraiVp0M40cg2Cj9qBfHakql9KX+hEI71
uAf9hw6QiZ4izlAUDq5SGy+W1SWlMRIh5ue4qPTJxc64mZlqqCEmuVw/cHnPSeNQ
TEME3EXeHfem/BjksC+oIIulqX3vBJrmyqpYc9mzpC8tk2G6r/nYiKP2Iwctx/r5
XVTxw5qYRkhqOHAwPAc+K201dxnRPT8b4wVf08gaQaAa0TbsGFL93h7wzR/Sad3U
t6s1/kXe/lQLQSLopZ2ipRuBFIf4zCLEtd5NUasFfT8k8k4n6wP6AoVIuam0SaqN
igdOsafFlkTPCDxd5+gsPocLCSz7Zf1cV0qxGi5VqlikxxCuuvHNN0g93lnUl9jB
RuaoNB1OsHtlDqdVORMtaTjtpj971oDohqlM6dnDTHHxqOZHVRNSEnHjoETnf6qq
EQ1YbO/dAB2xkcKO1V1PshV1OO6xsap54mGB2rKUa51bw9DFJRlMxrKVcp8BKbo2
OpKfXSXw+xE3mG+C902adVjLyIjTgY8VBDBgoLrFv1IAh4uZi5CmTThwEt7Z9kQM
jQ7JmgJZbA4vwDXFa89zZ4V0Q8MXVtchgRNKlu9+lLWYvqVl2Tvy45A5Fw0TJy/J
9Pr1t+HwSo7QM5F+9r8kv74bd5iLOV23o7eyMRBPnqAa6gYYRQx1g9q+HaTklm0u
vHvgcBlpU8G83nYPZ+C4dDUJCqo0syZMnFP+Q2dds477nIS/sjbe4fhx1yL023wZ
V036ZspP0OLV4uymmV13I/4AujTFmrhRUTBuvz5pmH+UfVnarkt6BlufokCcbw24
TJe0Pgy/7I1+17c9DG4vfsQtW58CrSYu7cBtyH+05d/Lc7ZF0b/Xu0RKvQthVYKk
vtF//nw9tijsns0StyZgPTKwIryB7qZZHnlfDC2CxKlFy6It7GHSikdhYfRgZTDk
DPLRLVROjEoi7+zey90rvN/lpHkwc4BZMBy6bsnU7K4nIJu/owW+RJhYYyavqmLk
v4yEZtZ59+G1TyldF8qaJYWjB9CPfEbkj2IhxsISAAnTSu0G3xQJGIf1r3V5DbmL
usWeLuLr1X9KnvCJNycjKLOX3aM+yxSprRUqCksxnVtpwbVvKInaFBAjInGInoqL
KP9p9ld2CLsN8VZyMOaKPueKaA+MeP0GRuFClEZ2cPdCFUwaYwkuutBVXxhGGqIb
S+tpJHLVqlbjByzAWnHBAHlNzy3Y4wVE5tiUmNlr2tbG+c1zwHaj/TemPLk0/Gnd
G8kc92Ov2eDaNpuaakObWyi7ZPZGpqSTN5XSX3emwKqLB5KuzEGW+uGP+7F8276w
jCOnECcg/NXYPxfsaWSLt+myPLtDsWH6bTWBVPOY/gey+OYlgplJ1+4qPhbnN1xn
kRYrClhuK47UIWwLqz/s71SMp+ovJhe7ccaCN8UsP7OuSJLGbx6I4qjfgO0lRwDE
jmAGk5y/tb62f9cQxknidQup663X1csp4mbvZ2X9ROS7W0XjDyxoNV3M9XI5yDyK
nbhOJt/qIAB//KTmXT1RwQ82sq5n7EVIQ8PkaX6Y9xtm1jjO3CNFum80nwDvQZoU
k/hRveazcdIhKd94vwWHiMyBk8Um8jMgTHN00mIiOWed3taPxe5mxucTaXWz87gU
vdTvJPBDVSgu8SDqcE3Gy/qBJ4C1qxXzr1enXXeFdKCnkg336J2LhU/poR/lQOoF
JniRd0+6hg2EPzdX7DDcW6PKWX6k3ZL4QQy5GhpoDx6sMXyHh+FZQWXO0OO2cvll
Ym0r/vRa8OecpyKQNiZAmLPD8+GzL79tc2k9ex+dIFx6xt1fUJRo97ewuMUX6ihZ
6K+7qYPvP/Ll8n3t2CQ9zlw1vpHBv6S9pVIyUZFH4zkEEbF9bjFpKL9pUVjtDKoq
qpegEvKhMr+i0Euelys0/E0/ybIW07ISKb6aAwCtuOQkDfcXch/LgvB7/5YSjvZ/
FLvHolWBHnVzGEHgVGz9F+LvfAkZISxmw97QQOzub7STVpCQRqYa5piwLtXcjJsa
Ng7oQmoFsRn0z7Xqc1R7tut5IKszhe+GPDB14jxZMegug36R0VxR9j8MSbTtdiS6
qRIAo8MLKzf5SR1H4TH6rLsgLWbT7rF8d1MEltkr+VbiZUrXSLcPdBFw/BFBZiXs
OMW7/IpfIujj2jySFaeAzf1KMwm76AT26hykDg53JUGasfDpSMv2oQNgYsNa7o4T
iC8mOm4m4tzTXTPqSRrWOOHkU3Oz9Wd89SdIDdtKGoqL8RIiIeEn5sZF25vVZm8i
C1JOjXOx7CM367zXIMc4iE7x/Zon3vPHGDfYOXfYK78fXo6jD8bV2XKWGnx1vtdZ
j3pl5X2LzewEqe47RDOjtQ6Yjg1q50l7hsEUtejfW+xfsZywhB2/I8uiFJAxuclj
4THKNWtELoJeT+as8pxv46gugLYzzY04HnGFF+Ll5Djg2SP29lu0HpSWNoI4TKF2
nYOcjJFpQ3w/ksYeQPDx2ZaASvgTBZP1Jkc2KQ2Mh0h9oeH6qCB+zQsJF4gMGsUt
/xrj6Ij70JoR9v0BO6VqeOlE9wqi/RM18+LD2OWzhxvlw5sEJQMpRuEBTMpUnh0y
wzEeS50jgmf3J0BkH77sJs/h1aATpdgWqqMpKAmas036KdCQU4uh+KPcJqG6I/V7
nRlcpiMQ+y5P4h0qEyJKgWaZkF6UV7brLJB7nzzJAXRkQKHxh8auHiEheUYOlPdG
Hs7mnwxn77gkWUCsqE9PvvDuVLtsz8m0LQal1I2pGay5qhWMiVlI5ePre8AbzRcl
ZeMs7wQPeJseMw+eTux4IxvURe/bJcH+WYAAMmu3Rp3QOhz1Zj8uKYXb6p6aqvNb
kE4fAkv7dRP1T5uo55834pRC9T+LOEfcPTXfU/TU6JxiruTX1McrWzLn5oHBOSo6
gDQbJFnd/RMg9PAbu8dwEXgis41g8ZToleiRW71vv+59oU84X334ei4qMiKeJ336
srfeXYEeDmG/ERKgzci7luv2i7M9mo4lFUxq4tbXrFJkIGy0J6cxcGw9aqxx1stS
0yy3F1NZkAhvedvQwxM3WziyfO9HN+rLlmS/bF1Y0eGP+QrjVhRp6X32IqgZJObr
JYsEJq4Yt7WzK6eWgk1CqVyILF16MYO+nVRQFyD3NcffAVhGNkkrWxJEL0fv9z9P
9HyS+g0vIrb/okEgIqKKqjImJFcrWZ9e0XBCS+Juzsfi8VPrEZZpfzXvO+Cy8Axs
9A2EfKfOqDHpgDZO30PZChWNCqsLrmAtnQ+W86ZBXob2cTEsx9IbaLa2YSpzcYIR
uRuGlhWB2vjn7Q/KA6q5bocbe6FshR+Yb5pZ3Sc5tT4KBKoXpR2siy5bLvImlYY1
dbvA17V1rXm6ahW0IWzipHA/UWXlVUXxh95+gaET+KsTHrw81iZ8Iq8sqvaa/lJF
cdqkVSGqJwoC6NQmSGlFpSKZbUV+wcCxzVX8ydhIBZO2UlQml4hFjTU7gxdKLWXO
CSblh4gzYqocpTgjhCHyaetwyTHzcYflfbLE+ogbA6/0jdHyXrXe5yCzxhv/l6zj
ROdrzfLyZ96pTJw6458fl2hCcSAWePvUDcxOJX1688GJY45PlQOjxtVB00yvHIp1
ZIfU8UoSxCvvhe6vzdsmPrN7j8yia4CbeLuMSm+1swP2h6T955CXCLjoDTBxmMGv
CePVmFLWryjueEW5vRpLo4x0ZjaRogtwsKRaqglf8fYFa+K0gd/eA0SVf3GuKCFg
g0hCNBafFLaiHzp35VUzUmZhUjndVli8GABFlpB7QOZtIONznZ/r/bkoKeiLe8Kj
SxKbJutUc+J9xuYC5h0DqkB5oQUbk5RqXhUbH1H6HZiaNOw7guPRE6cihvcGa0Gh
xb9eDWdVyF4m2P32gAWA0ZQ0jwm/huZMdD+gTbVcKUOY0SMASNYzhipyVlrb6ZSL
NBV1twfppUlJvWbrmVP+PvaOJI7WE+9myzr4wsMsOphAPI+MxRs+qY/TY5iqpnbI
OhC/emdBi9CGft+ofL5p2++o/0Hr7ClywE4/tS75fT2ETJM3X/7EsjllLkKCdedQ
pKn4tT8MlzHaeoKi8c2tQXYdT5VYwb1WstXm4qAOwwkZpaOXwhgGAPx/Dbbp3pY2
zq+fnt5kNOdecff4FTi1cvWlRXLl7V6YDbcrvEkdRL3VsPEo6goG30p5JlG4iP1h
X3xvlRvayOlHx7shunnQ8FAi3K4sfff1PWUSK0080rau/4BbW1IjyYxAhPq/DXAG
liz0q5W00j6pHCx31uXMeBH908PUip2WVd+XW8eKH4bj8zmBDiRofXxNv9ZecoB5
4Q2QlDn7c/zpFZvKvL2h2MZcEhuCdYvzUCA49vHvD4mYlOhLYIZRO8sWxnVUH/qt
PQhnzpxSJapCGlei4v5radI9oJ59FUVFG1DZR1LDY0s4KM0J0HHByFRuWFy2Sy7W
LOGTRLt0VNx8YlvAesOrkEvl2NEpaPVAe2SjfxexFgYRolrsPbGetF+4mU0U3Yw9
OcCkR9X9o0jR6/N4gtrQsQn44xUS5dMTt/DQt8E43DGEeRtC8sYhgos1W75LKnMQ
karznRpPYUHnJDhYVfsetqbHkAqBzDRPerx/1nhxNG/6kJLyKPDZtLWGWH0XelrR
4tQmoHdQCb4T8Vhc6jWDif55jqlSJ57QElvz/cEAt5bp8ss7NYxD96AAGqhSeatD
lTu216GpbNb5/YsxRbIV3r5kgWayEdPQjmK0A0Kq9/1xoW8BTArz7CFqlxkSuSI+
I3apYqwfweVzqiYM7Uovf0b+d5ULKnCOuL9jStAAkFM0TZE0bvkKQfUY10Se3N2M
P3PPOyVuuK0prYwip82h+9BTVHJ/txGo8B0FjQbuSgUkOjGbhm0nRXUzWTzetibx
HBA/3W6j/xvUt0UEaLNyP6Cih6wEgSq+71JKHcyrscg3spk4wBb8O+omiDZw5+dp
fXTrXPXxwp+PyfQpuw18khvDU6ot388Q+KCx0v3AXc+yVUDYSGVYpJQ0BiQkQH65
AbqJ7Lz/Ei0gEKPyliuRgBmrfqRObSl0o051WDK2iNOXoPmF/l1p/aR5OmJIf2NN
ZLlcRoFkQT5lwJgbqPr8CXKlEEW0YFEdo+XNQ7PURDHnwC+mwN5kFnLIXWuLPh4Q
nwsuQ8D9UEhO8YHm3CzWa6e5SzN3iZpfTwyyjocCjFra7ALBT1kM22Il9ir/lvqz
tUk1RBp5VQwEYMoATVgeMr55uFoIGJq/38d2UdMSsZ1T0e+LmA8RfQ+Y2na3JjZT
tstbHFKFdhQPF1X+I/0pCxovOExhqCxzc2HzFNwXAyHRDx0+CRexJgxsPC5KZw0G
tYa37aAS1neoSgi2IkOG87cZRaDPFuJvcIFudwjjqzfx0+uMPUNAKYCbBDfwC2BV
K5tnqlKtEDAbaFM+Dd4vH0fl/kI8UFVzf5GQMnx90xBSw+PB4IMd33ebTrImLFyX
tGZBYlmtKsc3tc5rYYkqiAQbz3861xO1Q8Rd7tzVaIwr96PBufS+oWMKiq3OwuwB
X5b8TtYpjQSIne9A4xBbDxmWLy+GxzBKCVsz4G2DGIFWMqzn7NuqyBWXx1VRzt/8
/Q/1BPF+mq5LqEFxDIWWACSfygFX/z0y96U76m3l1xtpg5mT7tRRfmDlubTm2pAf
VwogwdL/z9nfJeDiIJKTz4bgo0oaFChtoN//4czL5gVw7YwRs8UQSUtgpx1Avdti
xRbE82fzayDaq7bk/Q8fzhDoTErw7P6mNbtGrFZcOlmLDM50bUI9mHrV5Zrcrt3V
h+6MPylHAhhNOccLfNJBN3sSGc1V+xmj6GPqjGWyumcSpeKrrWjYGa9TMO8lPJeh
colLbj+bvorsiduzz+5dn5cQcFl0v9e7GNQ64hyWINMPgIRiBgYZdG2TukXbgSgN
tvjfBFMRT5T6fRIYjn4O0ii9Y3CH9+DoN8id2hJGqWjtfVjCqbJHKtSFNz2Bqjqu
msKRAmzU5LdTrNP+3Cl0VY0bHoOtPNV6Mtu5cE9wShGBZdFTxeDYtffoLX8cUIoY
O2gzhx2EKEvQTswFMBVocHAm/my6Lzy/CnLvVSgwhbtdCgVisFUtIbdKTXL6I1tr
AbH94BQfZ0OBHqocJEVxCvoS28D/0zoW6o23rin2ES3GAm7qZIX8aYkPswsIMeXP
aL7qzucfWR3S6oN1qiGGTqRBqUws17OJUmQCNDCCBJ+IqnZkZjEIpvH0VXiNTH0c
cZS6DwFv7ejKCoLaA8wUU/kb9xq+5kFbQDc7fELqQ++ZemaVmHpkLGhTGLLpfjlg
pbCSKWLPqo1nDIzbCrb4yiXfxWc7YfleUl14lOndTHrqtmvGj7DqMyYzg92Vpc42
tJ6WgB9Vfge8G/9f/cTbCy41FZUsEW4VDBqizsrBbCaMsttE1tJLu80cuthVQgy3
V5AoBGlHygMCZ2Sj9UzbF4/Z9QmB5kko3nycAdrQYkO3YXenrZ/g9QStG3lwHgLX
/E5g/oYO+FFaNZ/57T1qZHKq9tzpAyIhjoCSWYI+dEvyyrMUdu8boKiD3KliOa6N
gqZVenTNufYpIFjTU/YMYzp7YVRz5Faq09UJ2ir7ZS24jnuYyR2Qf+6h8KYgEiiE
5nOsuTpGlXqSbUh5RyxknpkHN1HfivUIJstbvGEi9c2nVd6Zt0nyQYt88inAi0xI
A8DQjpQpuJpsx0XMXKcMnePz67ZSLPumBdYyDg2wsgf4kcLKRlVclOr0e4PYe1fX
rXrR9MRBssI3xUZOmSOjBnb1R+LrIdglvLrl38zYtN8HF+CheetzZ3QOSbCmtCLl
36ADMjbXpJgeoK+NcHf3wMYdlApUFPxQEIDrcQHnjU3tzF+eNg/0hyn3kyH/Jz/h
vDONtaZLLrNOuoKg6xm9gUKD8jNURzGNcOPIQvVilJ0/vuYfWc6j4Q55QLo6YBVU
/r6dQ/+Htr0/61RckDtV9PQ2y0raTtzWO4gLBDI6I1FmpLYQhEkJTyH+eG5B0rga
1VC4ujyJ1a1xUhYVujrXzxEr9/yywpHCg49O5MQkGSC10lfwGA98tVP6qfIlv5l1
KggvZdGP1QFWlvdR4wULp0WKBa17eXHDYzrOiB/7hOPXvLrsQ1WYrLvLEHfkzLDi
1sQLoechcO/ppYKl1TJSMtrsRumSGXEzsCX8jObdNlHCX8Oe7M9P82RHMkLvDmlB
xdvNDOyPDcYhIU9Acfz6EYBtjE178Ke02S00jjJrquVq/e02RdV4bt8MqRWohoAO
L2QFNoofDV/xFpYv8G2Lr2Fs/8caTMja25sbFs66u0tGSAUM/FRbaSiPj134vJvd
d9be2DCxkEunZrZU0RH/GwcWmD+5aNbGUJ2yxTChXJCH1JsMINVtxl40DxGvepbv
XzVCcB1K7K6b8l80CJsTlXwjfCep0cMXjamjP3xE6wr7lw1WI4Ts/BlfO3TtEBLL
UYsTcaisy0umIa63Ginvlc/AN67BPHrRQd35/FhvmjPVRsh9h9w6ocLBhMMa8guN
aSzhtkJ7R94traygcGdZrDhW9FduDWy+z7Rhu2fYOY0uRmu4q8OP6LZ+fGVCwnkB
BhEECNKB/pix+V+LpBeIv2c6ZCo1N6C1DW4gtkOUHrnbxh9dQUXNSZoJ5dD5HrSD
p22s1tnFzdj7GxHluJ49yJEq1uWt31oTkYaU/T38MA6li2DPJ3Q55KTEHs/fXzsQ
NGfHZbwbEhNqI1as0WKapsxVmTe36ih0JVHNv+VoIW/QBpzovf5rJCR5OG92/lDh
c+LpHt1eG0t2T7nlBuAo+SH3SPXdN7qzTEcy3sp9VUMLF58X3Zlh0pLU44oTsGcY
F+ny36DeqiasyiP074WmdlS6GPebJVZz/l03AQGRoHzF1/RZb2DzS58954m6s6NG
dxMwQSFgDUxIdW04K78v8fqsgOaDu0FvNZpAjQfla6oW8BJZrAZCLruIvASNGRYR
u56AO4nSI1KOTgp6xV3/s3QpDSHGK3QNxmo7whGj7NPGqM4ekWXd8AhVz1Du+X23
fJ5Pu8Upt2aQZWni8vErYyY/JejxaLq7OebVYA7AfvwnqloS5fvbVMvgxqx38lbH
R6+1gjFkdnoL3HskmWUVHbfqSVlFpC14pLeihSube3ggM1OWONwvRYl/C84jNHv8
u5DBdz6Jcvxmp8HcFBThM+dkXuOKUqS0tubKRL83usb0oQ3h0RILf25nW7BU2DYe
Jq8hfiT+0JYn0lgYAApHu+1l1MI7LQF6bMCKlHgAPeDG2/o82Xz8t29kKnX+TpME
XZs7kqzy4y+AWvcWDf9sBQ8KljIp/lhVRpTAYELf5R14FHO6YE/n3dlEJAQF5iUc
vhvieP86LbVYE8Ga1rB5T0ZfOA+SthkwEXRfYl0kLaaGnHH/Rv4/fHnU/NrhgYHP
ndWM+tyTxDDGTLsBv2GrYK9noGBEM/LWZ7Fgp0r8muOX8mrXAejdJyI1WW4LmPQr
53XRepAPUWbEx0lHMgqwHBmbM1Z0X1OKyFxguRNiiSkl/sLXmn/LZggUHDi7skym
f9MU+dTTKhC6i9LxfBMmM8h8TIbrdYuzyvOK3GynKBT0Xn4Hwv15aaNwMwbB/iqH
3X6OUop8+5V87NBHHN3HyBmXjZwis3fnQx5nVKdmKK22DQMZNYPqFXusUETIMU5C
z79OCG+mU+Psn45SUSS12aRUOnaMXsjGwJ50HqK2RZbDsfngyeePMrcgYfM3bwLy
t4ss0hiyscZyt6+L73fysMzE4jLMuto4MqSLnxZLYGIYT4hTQXbKuWtIVKSwBkVa
Wrr1ZgcHthfMzWqK3ih7oIzjLpbFVxqWdIpTQYQB6qJgq8Mq1ol00YkWRaoa+BOp
qMOEnflZaITMxpAhD9mRtVzk+18KmlpbKAq/5Z64AiUtD0dCVPLzRGjb4GVNjc54
/8s1WBm8Ax8gW9WnZwTrFd58og4jV/cl5V6O2vpmxFYEEDmEb8QaPWJTjsdvNlo/
IrQq8hXcDiiOyFjgfHsfTcxdtyEmR3VdaoNww57WUHpB965ksgGCkVIsp7pmRadu
C++c/j6ZgdrF7HAsBotZ+/q7z8P2VZuKjMhRZKzb+xV3kfdtRRFLHWi18A1VzRV8
xh46FIU73b7TLKH1D0hdJWOgRPaYYjuL/bwIou5EU9VBB+KU/otG8n153IjAQ/Cr
7GIbqbgr00ez6uyDFDDtEUDlUSKF23yeg0Bu9FiomfDHI8SRPbO8NgdFzULBQ6MZ
WXAY0cAtsuChK1JBJjtGBk/JcfwI+aO85rUI6zaPFSIjEYuEybFbKET5P+3aqPWY
NsqmS9KQSHNWEwKUSyL6KcBBZegqNHuaQlMiuqDAKFn3VVyw4VHdkvSAfMkzqpJb
6dPzmZh7Dy+3amzoLHJSE/th3eqiizEoWZ6YEg7W3qdbBG9nGEG4XAq/SboSaaZB
b5RxXgDIsoP69J0SWLZhaokkWCyDpwD/66Xpw5h9cPSRaASK6f8hgUyLl9qqwUyq
+E7+lFwR67EQHmfjP9Nc8S7ZH7Nz7NCbToRJs8aYK2iXOZcfl2OEA0YT7/Ot7/sH
m3xHfsxjzvkpJpt4yZiNjZPSZNsY2cEgxTd91bbTtkGS1BsMy+KMbYHb9fJ9KNCY
kwSgUrrV+Q4UXgvEAwoVNcvHd1vfzXLDykb9N62eq5nptlgs/VsfaAGY34jsPYe7
xXiCjGD43O39BvFc9gXxqpo9pFvmU4Yio0vA294LDNORA62XSr1vlXliMe5YZDIb
BCH6+Vxry3HeGythCiJ9O9TTZPkPmd6cUOS6sd7nUZGOwxli4Q3a6tQhcSYa+P/k
4eq590N5M8Dm2ARnyonzv7nDWxsOFv04GvkxJk6Tf/7d8f1/7YjfaoFSwEQkvyPS
Lh7ZOs9Kg//IdTM5fqIi9MxrB+EbOUgQdR7zAzW/MYPbxoxZBvCyzZzDvaR/Zgfj
/lKAEgPKAq9m9WFa/Qsr+tu0duVbYm3+4l4RUH9mgQRJFGPnZSBklPdKzJ5kLImN
2WkHMO65rznsmzjxV61WZthxeP89gSOTbS0VUImPbCJg7840vPR4yHPhuXI3tg2b
vBJeyunrDLFMwpOCNaI/apdDS4Rs43P4m2acwhnNbRYaGdjgGLV33S7sRi3Rk6pj
RQ4z7cOJEVYzPkKKtsuQxDgRvYGABhHIq+O5Dyx+qt54+uRbVvxLfwNTWvkFISBH
IadGXAiiolml/EU6Bh7xkJWTygo8zsgGC4LqNmn/3PeYwyb+2G+e4KC2gsAS/f44
zTI49uXjTeT+V3Km0IM/Ck4VS6rysaV+aiAb1BRV0zNXjjHdWUQlM8YDu5L8P6Ti
8YEUZETPlax9S8I/PjRlgrVlXSHOMStqcFJEdWCQ7iaPs/0Zzj5i6QGDFKg/4Qha
7pst80HVVoi+himHMgKKK6CBJHi7JgTv7opxw1G1fYjtBmIJ9hemEa9QnJuUtbd7
dBiw31JJq+tkjcMT9GZWhdtSxsSBI7ZNiDP7+YmEAkqpvHmIC4rfdoie5w0Y79Nq
LY6If3hTWUuPW52XarIF5cbvGPmO5GtfhvYtI9YzaBd21I+AdjtmO4br8oflh1j6
5CGZh6Zi4WxCe2DQMQogrF0iNHsk3/zx033urMTiIQEWGJuoegMKuIOBCYV+H5zX
SUTHoj5ZtvDVkE/4cnGNJXnIRLmpkAz0J4t/U9FNYE0RIFr0uPekFhPpQ8gHcT6b
5Yq8JavdqJed3LDQ0kLcNhOBnFlTgSBnESGwQT7cRkt6rg+pX3T2MjY7hEvt3MlN
HETbhJLI79fooUdUAs+1Yt3VOn3UhyQN/8fcu0v/0ZJRbrlJSzxKMoSjXr18Cs1j
hSPr7fsVtcifyMjbyai9Oe3bi+bx8pW/i4m5gLqBgMqIqA4jMWSvS3stLfCcMBbl
lS3HDyyaVYOCFxadBEpf6HjpQCk716qqXPb6pstNIBsDCWOtaYtwwUZiicDq2sls
0CoFT/Vpm2WWM42EZf7CWYiaLN5TmsODT67ymjtevSeEdvEaGq39zyQZXl0mHS1E
0At+2i6EgYT5cM4jTccRBUGbboRIqwnuvTXx+tLsL/QH9GY4BW4WRi8E15pr6MAN
n/6oMwTDu6T8XL5mEOBqrVyl6AuJDe5/7wwlbPoZUs0xTuhk0nLEZL2v7utp7BDW
KwSZFbrEGDyXqdVXqFGq9kAXhC/4jwsFdmFsvjUg4IHVcfMsQrCh84TQtGM+WBMO
ykx0Or7iB65bGZsqnnb8bdGJTOo6hXl+yNF43nSYeMs/RVXvdueCZUZCcLgc6VZm
XXp0UekWA4rkj0fFlmJsiUXN7pDXzj59v9YitI3Uh/DUbdvehCVBz/D57kLVtePP
RAojhjByS0kz2/ot73NtMUkv71m+ykZxAcD5XXmPWkcyBg4rPaJTLRcFuajRVU74
m1dwBuSYVCM7yXFZndqAMNLHhnWon/bzcBX7dHa35i1pdkvVafqBpV0bOa2s8vyR
VVLCUJZ9mY2NQlttpSCLbBat5DeQQfM6ARVMBPjLwsG8AXyb6Tkjo4NQwR/pplKY
k/0BT1uvm/YCWnIjMaKigItprM8mRbHQXmQ1M+aJGpDqwK54PwleV3T+0ik2ucYl
ojZBC8SenY72g17wzFBKECu6QCI5nkOQA3X0vHmxr/9kekQobr2SH+z+cMx8DWSF
rQvDsI5cimuoX/SZDhqirrme5TnK2en1R1WWCDPlH2TEogs5FkPyV89bqh0bGA3i
JQrtEoyK8WwP4vmRlj4/v/hqmRM53iPU0Qs//T8lFrcP3FynEUIwaVnA0rBOT826
jcp4saKkFQsbAHPePKsDcBqYq9KnruCa63JFf8RuUn82kK5Uru7V8ZSLR6fdq3iP
0kYUfJyfavI5e4d3TbVTgUve3DbG4aHzNkZNWaYIvGBK7HXMvuTuOTsbzIUvBqPP
aGQFYHtreMipAVATcTsOIMR8VKZTFcFZwgtITEYT4pE9NlriFc3YoNMrxDx+Q78h
9kviEwguaOgGdPZ2IxGprZydg8xMV5ARKrXke3ztQ2SMnpOH6gq6U/Q3RZv0iQhH
rTw+HLSiwmKFu3uOhmgusNLtEWldxbwiDIcpbY4uFcfPZGcmzr2gy4XFGb02fwM4
ySXaKgneQ3Nt/VUCeC4qrNGbPP+jqWjeccpHbMQ5OaONoUfOzQKLw7UcBvW+olae
Zy+V+beHg1FdxOXH3aiLZHBPhMzrP4cVEAGVNirReNEm87Pmlm9WFBgNpN4qoimm
FZDTfeb9ic4ImbzoamUyGsunmGg0FFBarPeb3tpTdE2WKzlTfdwhrSZ0iu+99q6E
t+OfFUGS9dZ7nwGharIdGctWMio8d0J1s289HlE3RlON0rLsWRivgeUPbafyrmgP
rb+5ZtaTrUXG/4dRfaadA/WZLEtJUMgfHQRteljiI5ZphAWqhYIzcU7kSp1TKwxO
qN8WO4HblzFtRVdZbPgYZzORaS9opXpb8NSpKS45gIxY9RTafnUtJYhLwdAs9wlk
nrIlwkCpdTx5g/JhVlLq1iRIyXl887sGZGlAezUwl+Vz5TxLyUvkvqcRM85Z2BM9
aw61VUM5Hf6aT0oEeS4Q2iBQkfaRA1QrBr7aDAixCU8HNWDGUqJh9wNRHwACm3IH
s+TSMnXg+6dEI8soBOTrqt0H6cVLwHbFPb5fWdu3l70FqRQAbno0PL7jwCGRGDEi
o6mZzgcqkIKkj7y7NIiCMoNJvvPnO0+FT8zSlnHYfQ4g4ZnV0b7OMmCmjou+yd8y
8qMlsTWH5I2gmiAqbo+FDYnDws3tE2S6b/riQdLFCIl8+7BuF6L/9VvXhSeApbfE
1uVKm5OQqPuuo4Mool1j4tSSxWgwQnFQxXe1NaMFXuRmPU65SCtxDTfsDpYkEQco
+bZRsEUjbJC9lcYdpS6BasvIGLA+JhSLEMwiq0d8UrKFViIDhZFQsrPNxlD3Qj+j
+Xrlq4fyvFb0ebRQA+BPUl3fuJEoB0FeugHKrdw0ao3ruyAIa921jUWra5IdkjE1
SHmFu639XvnnA1l17abvWK/JsBVFkKS0fdGH7nDIu5g8dMvUz/jB3a35P4enspLq
W4d0OBU3wWKN8dpZkXfpeY8OV5T9Or67YXsb+jAFZejAlDjkcyNo9xwz6ELdkZz8
0q6cKIbUwxQhCxDpmvxBt4vCDNKpkhaeXgpDf9eeQ6xPSoQDVjmUlKW54JTH/gD5
/rherc8rq00q+uwSVkVWec8y84i4YpfVa0+q/MDQ0hGafa5d66keHvRERX0E2HH8
cyT+ReJqTboW4PI1+M5/Ztn4ARl5zo9QcWet3aMagvf/QzFC4YWsINq5EVltWRol
LNc6WYwzs018NkMrw8OETq4GD1cxawTE6GE3sHyfUcqfbIEIxQDlLWoXBdXh/fm7
81czMGnzwJ0iKuCZGFdzJqUMaieSee/LXLuwpTNsd0jTA/xpUEY9oTYIU0qOipxY
Gsm0bkPWop7qhchnDZTiKmAXeZxo/HPM0UTBTQYncDGDJy/RJxDxI8T2HfzULoLq
P0UkaZrLirOf4DR8ouoG+7DHQANiRlKvL2a37ad8cxfXSGPL0N4HILpV9L7iPpsW
xC0qrmQikVoEhBfWfMPm6sAjUv6E7925PWeFZ9pMRaM1BD7tXEs62Yqb4hQNvoBd
EXAS+imr6Q+ufQw4xFZ64E8oPGNc3PdCXa9Ejx2vFEmDwUapP8LuTNhI1x3HEBVC
N4ENSUNWFhqzSDY89L021pk54NdXfl6fTwSRadEGiatp0xpVN4n5+uyguiKDTYor
tbS/JL4neccXjgrOJ2daEUFlD+29Xj+B7dsKMPjlg/DZNDBc+cmh0m0aBfOngqH3
ksjN82Vf/twKXnCgl2xG0Mz9XKYrY3we8IKI7EWYM1HsgAqkMGC6yvIXXWgQC3NB
cMinJbMrr2QeOVo3zn4ZdZrkYACD6xVJT3HgwHWv6qth+V5cqtDkCUdCJyMnuelr
TMHPrRh66F3BrRsYt5mmX6odGi2m3/clcriHf0UTWI9l+PQ7KVrgDo7HhS2XW5yq
X9uA8Rft1cfbHbRCLz2au7/0rM6ZwBKCJF79TkIfzzB5vg698LuaJKYvslOj3ShO
MLborILw90jj5BTLFH0E2gFEI9Z4VWrMKgKoThenHf8veb69n3DV3WQKWPSgEuax
uYHDxX5ZVf7GOCEnM1p3VE/84kbA7CexzV8UEMG3P1pQOJO0mA0Gntsb17mbx0BO
RuUAzfZ5QXScgSLIg5QnFYNJLo1DuuzlXwlbjoyGzlm5OMLtwonz9q6XyrxLQLDn
oPvdjn9Q2ojhBo70E/NpHynJTgNuaVE5ckNIXvcz+fNjtqnu3u+s+RECcy+jN/YS
eMwJdV3o7pb9LrLJ89jPLZbcSof9V5v5YJ7LgKa0K9/2eI/6igskEVHb5B5j9c0S
0Z3meYcvMU7YsXpCWV9p0tnv/Jv/rQu7yXk0yYDXJCDvVxVQ1kgEijkoY/tMrRpe
8cU/FDL+RjtPXZJ84nYBjvrEZ5O8mIO1JQY9buV4Jo3lFwT2705V6PVnCz9FkWfl
6+Pzrkjl+6UaFGTCIy5VqTUrp3iaRrvTZaYePMeNbyuSGgFjSHADdgCHv1PVTvH2
Q44y1B5/Y9znWXq8D/jmEWjJJsT4IMTKs9FgM7JojFCrDr+r1Dp9NNsiMvg4lhZC
QXSkvS42mpeobBAA6mTOTOorm8NnO7ffwBZCeNb7Ro0zbaONUK6BHOLRVD/x3eLs
7OcQiAOXvv9B4y2ub+YZ1T3PN7P8vMZHHq3LmN5OHQH51YibYYEkG07jsCRSH9ZY
vrK9M9xnsMHuFpDr658oKPDoS/u1h0gEoElVG+n+AmoYegOkn1qLwUa1tTnicaJD
mkPfIcJCXM0KyxdYnILxRu6l5ECsFpE/DFq8SIi1GWinaRfVhgd5/mFl3K3F1Jvk
JJk2Ctwknsz+efNIqhN+yTnggNOTPCRdK7ODfQE4Yoo1mRhSug012wgKVPhqcoPl
hLkh89gnl3JGE9hJDFXCOhUjCYCCbrl6or6y1mB4C8R0a76+kx+iHCTAh6GLikCd
3nhWESvsKQfHBIarJXOFRpBJ7225C7d6M7QHnBkSIZ1TGfNCUfq0MxNtijBeUT/y
TmuWIIk35uUru5jNjiNQ4yiIkU5UxeGPPv0IxHRK3HuZiymT3mbF6GmGOsUrekL7
x8klGxLwEm5HTdU9a7OAk+QW+G3GwOKt8cEuqrAW8RfeQ4Q+Qdwhnf//6lQaIayT
6FmSomkKUjfI9bYTKuCpDFut2lOtSBvnZKQVeenYslc83SMdsiPzL9CAS5wqt1lK
purVbMrJJydxCp1V5fRfipJA3w6wj236lQYJsUC3jUz8jPiFfHiEzkyYx6fd+zJb
QiNbTo6Qtvr4se6yc6MRyABpUzn4wxoJGOz4zkqET9f0B6ydnbHCjat/q/bP5KEX
kLw3bp0cPMvSfmb5SSZFyVjegtwPV/7FphZCIjLbatKC4eLX8MJJqAOnPrpMmOJb
zBU33cNt+56xDzreIM796wInzPLCQn7ADGOZf9FlbqDLBj7BK+gPZFtSjzJOqlyZ
PMUEkIE22RatH5zUNaIcWNGUoB2Tu9xeXLgFgmx4M9er5DxycLkQZZtHSjV1IKSs
u6E89xH+5R6ncY1tG/CcA2S5E1249GPqWolG1uEUHZkx4YBraG1Qx02OtkQDXMXY
wW6uihZsqoSj03kOBps918ISn400bIwpz3lqvXhxyUNMHT88/H1c4I54uOsgSXnb
lrYtlrrWU5pnG8EYTgDDesuAbWnQhvYYDCdFqM41P1P6diVKWi0aBN8Dqjdgvu0Q
QkHBfUKij8wlNO9GCbdcF4bFHZckxvgUsULJncA2sUhE4lp34nS/89hceRGwlhq6
oo3i2oldLOa89NLi4oIp5+G6bGjz8slltRCmCSoRfArFAoSonZ/8pGMU7jNkWxp9
Y8NnDfDjN30JJCjqzzTCWsiDYt6nY7ch/veI16VFO/A5nMbS5vxO8zH94cvyQ7Ho
ktMQpTty3dVk6TOPuf5RqB5RleWDuPl4z3GTtlfvX1gHMOCh6GfmVDewalwC5Tdc
fJbNoQbqnxeSZrOkVjFre6W7OJQw2CWzGaSXrevByYrkBaAPIQmHbva5bZrRs7Rc
IJxmcpvRT6dfHYoS4p/oUNGl5xT4SGRJcipFw9pX731OpwfANKByl/03O5FKsUwe
Ym+yBihC0qBBkPiF+zIgNIfzQx64yQcpy1fJQmBCH55sCLmeNvgg3iNm+qmUWc1X
RJBVDxNs8TXKbN1oTCmSyaK4UHAIwDfge1ZWHPlKwlYUx2lDbV5T/y3OJv7edUxJ
vJI5dzcD7cQ/+SJEq4LdaKaaqY9M/QBR/09Uxyk7Q1FO30pktoSr9UyWBQ171yYl
+cC4BwWbA4xi6rlB9cqrCfKvjZNI5v2fyj6/7AHV3OVCnSxvxaSNLKXNKptPo/A9
dvHw2cl+cuDsjCW5TPW6ODhHdh4NQQYdMWRDeuv2iXoHKf4wJFCUvChnmefdLZXH
FgKuOiDVT5rklaJ2CNifWGfMbZH4rMXO+9EIOF2hwSeuzIpJBCHsIlkRUdDVju5y
KTww7mWskSRkytQqVQvqUU+sgjLgNGSzc3+hqStKXz2U1QL13NPthpdRsdSE4xP5
PQF5jKHDoTo4CYtco1vIzpH9LPQo9IsCkUfVu7BJoDl9FXCxIUSqSulAAHny8/BL
sT4RCW0osqVDnfwfGFoy91R+UysdyMDUIfmltTlAx0sgPXtjc6V6zeMRqGJs0AJu
D7DOYDJj8Y4Drkm3358ox0438DMu3VWlujhUMENo0KpeuAV7Mo/4l10uE5lbvfC5
eppIEpoVdkpilfYCo6SrXmQJxr3Kt/FTU5nTWmnwojQQ+Jv6Ht7Xw7Q1LaWcfUqh
AAzilbwscgIRu5K+ZY2+D8VUsss14viFgDY7siOZcX1z/9GZ7DGBbFaCfAT0nSxz
5+RZYvuRQVKknBmN2EQVzOAKEYmKokEFUdDk+jIXNeo9ZvoOdv4TZdJ/2NR3B8rW
4BaEZmeIhD5j7QAYoTdjSTIcwdW2mXbb5bvMNUYvt/UOfxqEy2dSuopmvNJwhvcg
UWo720wgP08a7mY5fsGKFdqFPKvYxsshU03pxcu/vK2dPIxHyMxXIBWx9m/OFNlI
bobVd4qDiFvBbpqRXfIdh/fkASNnMGGTGPbO5f6eLbf+IaNr7/s+eUZCUx3jJ5XN
jAllEAYe7DxfKbH+gI5307Im23zODo9S57gBocuzH+1z7Y+m5y+GbCeaj57rQG48
bnp6iICnCKXuLLqbI6gdpE2UU8m12xxGSqNomqakOc4pmQiGI3i3PfTOBk70/9Kl
k9W1O/xhxMFSMf9AxBhbnPdpIHOkZVBXyiwICyH/Oo2JAxlsfdusH8b6GvEoBgxj
ovyeIilHiH7N/BDVN8FD4jNt1nJbBp1xpW8XI+BB8GYsFCkm2yM6ld0aeKLbNgk5
XhatOIn2/Xej57ydRggGH/qn+bajK/f/odgUQJA901J8RgdikIZ+CcgmsaFST6ms
RCIeH9PhEz0GWiLWA1vahaQ1LYu2n6Ktl6EYOa+dLeUydT1fS7QlNxHAb6hm4rew
q8VUUa2dm5rNXCnRZbMetiNSdHXSxPC8EA0rJjseYvVbThW/HNVUOn8rjIkK5QyN
eIzVUST3S9gjZpSZfn6vKKLPF3YMtH1mc53NwvCQZaII6jEivnsrtEteh/ePEbBs
D8tNHWx/flBqhGTYQMLD+5zO2y7DegxtgMNAV6Au5jOH5kSDHNyk/tWOcpoLJvpu
mrkWCnxWVvVxV55V8wzEh1WmB9gBqvn79fLifPGQcLFYO6RFJ9fYK4pj31zb+Sl3
QczK4UExM0+yRbqYmtCTDoQkJlAUxjnIQVZHQQzglNG4r/dAFzSjMWGNjuBqiDH8
pOLSAjKyCmiV6E5w0jRFUxuJFVZJK4fp1b71VT3ENaCXTCIbXdPdmCdS08WAQ7UA
2NyBHMbULkQZ45xiuZVKxb4p+8PnENDF2rAMlzz/+CEqfdw+NKPRjUBee/6dKNVE
67f6vuZl8ejt7GpiwynfmWQ6Ue/G8D6NS0Ly7IAKBGHgfwyt90Bd9S+B4WDkMZDJ
2au9l7Fw3/AZIZ1n4hjRD2bzz6E5GX0pIEQzXjpVMX+mKR8CoKOVfRigv2N+EHrQ
/HH8BD/IcoOq64gm+heHpr9m0dIK7diAE9xL/Gz4Mi5EysEPU0MHNUT3hCagJnWF
ZGrQqmH1OXV+NqtFxj/PA+FRrVhqK2rmdlA2CQ7iHf2f/lvp3vZZTIMnAZH3FPEx
Dvsww8qVqJcBup/jYJCPj/Sqpe36lmMmGcSrroyNnFrEhFuG52Ftq5inOBCAaMel
1DgZkotchnYJUZQdCm+ZUJog2O5FeUqjcRcgZ7HnQUVBookUQ7dUAWK4sG+3A/1T
0aA/T9ZP6VoB6Q63heDlveuf06HfvOJw0jc3sWAgC+tbVrLslnkgIoo8wye9Rsi6
3eeawhA6gBh+44MKfUe5F48a2rK0M2VmgPE/Vu6+xfVrVLPb5YWlxgYqUz960nE/
Zgguk4xXZPZrY4Xle5wjRa+N6cBAcNT+WLf5fgmshj4vjHr/DIMtPvEmFgZkUBKE
CN2MaSdE99qjST9EyXh23MMPs2A1qaEkcBXvnGhGApDzIE1JkMj435hRyLIY6zBg
X5OMYRz0u+P2TFwmeOab0I2vKbKf21G1Vr3+zWuNqAgudwG2TmLnkp4RwjIyKzCq
H1gVC9sipr/T3+Tc/rAvEA0k3vfPryInNvSPQpfjHU+wahumM82QVCjxUrZnA/Dy
J69okqabwqI04w16FHLkdiTxGF0RDw9N1HQwx7mi4sWc3i+VoBnxUh5qqU8dY7Hm
yCeuCWiP3CuLLPxyEuMU9a6hTsEi8XtdFJlwQITbNzZogW8kYYZDWaYur52jGhwM
0DvCrpwjzTDgtNJVNQgUPRrxstzNCGOz9KYX1dyIvQRrc/ecrACgk3k/Bvm8EN2U
2VAEbkOk1ogsfLG5cAUARmo0aHQKTE9YM5pWSFKQNOdRH1ix3UhZfBdEdUnxS3ib
mwepdsYJ//FM1FA+iVFSOQQfkj48CQMwd5ygHc4Tu93rcu9iFz7Eufr8HUvqc8H4
uoVrRmMFMQQ4wlnnHFoD7vNmEexJyOaaWrZkT2xvdyndypmEQwSxw1k0bstIxo/L
KkVvCbVbgeIN8Cy7h4xWOiTMTcUWropbsnW3+8r52K3cqztFZp//BqOcfWBFw8YI
E0oKAhX92l6GFocAZ6FhUksU0OVttye5xv9qk043CET3oi6hIwz9nb5ccXA08g4b
y6rag13gKIFxbSnbjsDQPfDbcLDs6ltrsYMVuXcFgmvOf9JrKKYoQBLpo2G2x/LN
8yUWTq3rSdFI/IyAWJSaKnrWTsS5Kp3YFspdpC+/fI1woKvbmh8GNeax3aCBhtf2
qa7fSsPiqq/hYRnVcFq4VkLJG4uGxJjaov0QGTLyqFtYaJw2YParuY0DwbY2lAdb
+giMYsUZK7jwIK82tgBmnEUPeXaOvbl+cAunA4CAsAu9/07KwbLap78uYdmYmBL+
MTtkNz92MS8obEKjVssEMP1sto5XNlnlHeuqY27FPKrZ9nJNpt3yXqDhk7ok2TgA
TQbAlm3guf60dO/HISlWP2KtwyU8Ofv+FcwCjpMUBLTxLfbsJpuDqytXZeNYJakl
X+k+94KYCHQNwqCJ7SRpDWlN46l7pfk/m+9JNAxfrMjPa3ZKYe77QytT8u6Q/Iw4
0vV95IdNaYruB9LCmHkcyA9xh1WUGgt0gckNT3LduzCDiwvi0/7ScZDUWxEq2mL0
iL4QApjWLRPNaUPKLOl+QVPag/gMGLjmvMlRll4Fvlj7nUZTaaGf/Q2cljFRoGp5
zObLIgWUHVFNtF/U+AJ9QqnLZD6gxyYgcFlwuAX1mqXO8vALJngAzRbJ8EZF1x8G
FpBQkJy9FDzEM60NwFiKDNtTjCwQhN9gvWW/5PgvpvdG00FNoFh1jr+NOwgwx8P5
w5ywaMUKVSJpjeRKVTl4HCqzwv6v0LXRiLy1h5Qp0FJ37j5feOP9kqpkN22MlbHi
YXLz42oOhKpVFg3428sLfvqV/zvrARvHMHSZx+NeVBGgGCvQxp7BRwFa0kDdizP7
WyVzc7CnL3K5jN013L1JX4RAkQl5Knnx/mbOUIrB5KLSZ0//AROIUZX9vmd44sLx
bJvjhOTVWCccDqEj7WPTFWLO0rrng8pTAAh/iEmIuB59cFMcBW/D+zySNkeBT9TB
CFEvlMQnGXdnAyKGpD7lelQeUuJj8SwlO1Sk6GSyLHGGqXOJpOHWuT7XJMJoMpL+
G2V3dAAGOh957FO+mvO0aQeSSiGM+DA8IBykYiPVegJ0WE/vvoARWnUgtM7TkAxp
ilTiAcZkdSs16iU3xzQ1bH76yGhJjM0t/nwnR1ZUTyBBUqa5K6Cl2XboXCUZFomM
HZOLhikj9VMh6/EtGZe+DoknKBLIa8un+CE0yBSVapT+Si5A+92F/qcdDFjFaNhN
m6pRQZhncbXoy+mIpFCYymDgsxwkU0wPNe0dfqG5wEtu7+vXSLA2mIdQPLpOqz17
vbBAZUlVG1zY/NLtqPMXB7DPDij6E1LLkhS8iuTKaJo29AwjUeTaR39tOYhNibdN
oo9FAiMPWSw/mhApafWbRLgCv/7qbmaV5ltnMeKfZSxp8oHesQYcHsrzDZEBbfw/
k/cr2rOUu6U6+cJT5ep+GgrE7KgU1wFdsdkCaeYeGuTKYKW1Gy4bYT6pIJgLzqKK
ekuUCe+mHMZ0hJYQSHxiXMkLt6jOzJlFTLtMYZQCFeQm8sb2Wy0Q/yp16Fb7BonU
jEPXXJMUovGVGuBAPHC1B8TmlOz4CyIC68Bv57Mk254/u/9ezrkhoNkrhF4BZFr6
RrVtavsq6Qz6fzZAACvh2Vs94nBW/l6UGdYgLShgG/IQ7Bgg/7s5lhjTsX03UD0I
iYCD4YDqMDZ32SSTLUI0g7tby0mFqDE6P8szib11KvmTNf4C4/9yyKSfqfpYNZr+
VE3S4aSMUQjsXqpIfh55aTS3mlOtX+YLkrFrr23n47dsGnbViRtsugLGBQcxfO7C
Rlz+rbVrY1AKSMg02squiNauHpr7NwgE/NRJY+BOHgrM8wuiSZraD0PG/3SRz6sN
dsr4gbDjRgoIKxbpGAqu//w65DZRDGZ0Dj2JUtm+xA+C/FZSgl/Kx6zVdVttPCB/
W+8JiqbZeGmmHJLfvjjIR9UkLHr9Zmx4VBShIkCeQmuujhc12NpWSL3LIKTVWfJP
US/plTi98rr96qYXyt0NMwY2GOPYSkVX+ccgjDGpSYrf3/IzmB0euSQNF8R0q5oW
J2telcQom+Yk8J86IiDg02ZQ6g9REQpzztzI4eHwSzq8svVvmLEYIgeQGrRFPXMI
ycA2dSRDK0plfs0hBzr/AJ/OBsXFYbX/CoWFpzllU9WW9aeEW62EcCFm2pRZuiB8
L3bwXrSSA6gIlJLrz8XjfQIWmZSjXEKez+WdOoT8j4QsuQV1cquXefM/DuyMmfR5
NrsfjqYzuEC7uJcGou7oC2ieHzZPtmUJqiS4lCwBtBKwoDKdVhRXDXb6AlSu4NQ/
1KDGgquN2ZBDP/RbVuk0SvLagD3dEii+8zQWQG53TTfnjvTiPDbGY+iaEtAp+Cq6
2kCChxgukA3MvgnQcHUCR+/HtfObnO4clO2amyVSYVupzGUbliNpIqSC/+LeLsm2
ZRdwQFYWoGD1HYMA75djeeTEqVdImvuyo0FMuUpQDlAMMDcmDFfqv8eke7mBnpjs
VOOiBG47eYud0tvjPbnyP4CrflYMq6rS5OW8mCqkJ/c35TVThTv0tWiU15cgD3rG
qAGL2eawIMvKtLphgqECUGl0dUrguY7L0Jn5u9fDSc0glB69dsSGR1C3rTFEUL1l
dwITlrOvipz8fEe/VICHinPsPLbUvlMaw6mgcNIodspjk96EGrGuzE8+yenwPO3K
k2XWBV7cATW2s3alw6TGa1FX1mLtjoOv3FLR60TdBQ4kOaTONI+1iCJtFa3/FX4V
17GBOFYCaomfPmZAcOxXxiRy0pKaFYiMJbwjPv3FaNqkDpZuSds75RldljSmt+57
54ks6mLPLBOkvF1HWdtQS+oneOE/R/VZ8CfnnHTXgwd2TCtLcnOZMynkgXu3kWjO
rs5waJmfWT++SO+scIXHimtc8idQCFSTe9oMjM+IrO5UjVAkCmjernTVbzJNl305
01Su1erkQI+jdmPpFEqJ8a5/TMc9ENR3uDVhKzWCN+kLa2RiselcPY+E4h3V3aLE
3Q0C4eU9ZG6XBAkp9Ydpt0wtUB114jSfbW6WuUHbKuqVtwJ7gjvhBXGZsqt1uQ3u
r7f8mffBm3mwk4lJLZr9pIha4Ln92n8X7B4EmxyhRoJ5dikY1WugPtkgKHkuw0r6
mvo7oNw9A6TIGZ2VbejfFsbHpFnwbB6jL6AJihEfP034Lw+PXlAZu+i2acOsmmG0
s0n2XodB+R0Jwsnf8ssedEHC7REaf1/3GATKV+T28qqki7zzX1wQVCJnGku9fmm7
aS1UTnxRrcxt3qoB3U0DTB9PNPNl6HZwQR2B5fR5+KHyqGbI+kKAxlJYuv5Jr8AG
R4apDyIyMMdFCLvqpM73qb4DFhtLBV3o4FVAG62JQGPCMfd7+No5q/XXcoMjgP7e
jEB2ZksFDHURg1w1pvEhkxVSi5JtumQip5tI9eC2x/gJeM1Ta2WLKdwEx5908rAu
pCubSCx87EzSMUM4DK3xBljpN/+UjQ39asGB1UebPrLwsh1cM/2qyJwjnUtACqU9
BBUeHQ0M1fO7dMoxErw1YY0RFl67ZMHDOQU9Sp+fBDzLtRaqevkBJKnXu0Qj3fM4
IDIM89inyRIz5V+iDNVm4VDbRkKwF/kVYT5ynHzRyfMvQ0jjmTMCHKghNfnuObX/
KA6eFETV7I3uZYRspWHDaMSyYstXOgq4z2EaEliYMQ530/4qzHohG/V3f1ZC9bSM
HLCZig37zo1X8n//yNgDWN+PM9Vejld51HtGUytszTqzs1SEWhTz81GUPWsuDgt/
I+Wpav6bgm4MqBVijHBzAmIrGK2Od+LG0u+UWbuI+Z7zRbULhxjyvSPG/Y7D0Mmf
AeHASZtBK5/L75Jp5taa4nUxA7htmZ9RIgRITFG2zs4EYWJFpdsqYsLi9DHhmQz3
ba773zN2PFt4+ciNOc314W/RfBnrwBB+Tynxh/vFZ/HjqnLpJOpFqgYLFiS+XLS/
rmhSgIeNQQVW+73w0nOVIIy/rVmjBPWUHX17vaqhlwF25FbjbCudOEKaD/K+0cP+
iFu4VER1C7xPt/+R+SzzgkzuoLDMK7eZscmZQYIQ8fXt0dR6VGi91CZzGwlp/49S
NqMWfTm80tDeF+GiwyaXFZlP9/q88A6IIwZbGb0HaF9qgmtephfws8y46Q6EC1L9
UEQAmCuip1uZzZmyeq7V+WLCOtkulao1UjEP0acpr3ooFvOjVnCDyEAag0KwneY0
FMkEtOfwXIPlscBAFAuu+gmAJFE/fYBYVvxzp9h7bJinD9QmyAG6emiffBuRDoXZ
hFeBnVQ3Pa60UFLUQukycagt2yVEac7a85cQeT1F3/E0b7wkZPLQOqYRQ/F2tyFY
WtoFpilu+seFre5Y2iMl8Wa5coMX0D1C3AFK5GOZnEmg16F/XlTL+vgxFHnjXEK0
0wJegdxyQADDlnLADb3GOU7zErofMwO5dpW8P+7YI8dB0dcmCc0jP6fRmH09l2y5
t1sx9iro9vhKxNsgVYL/JRK6dkdWuIqzPeOT7Gqake2NSItUyJkqgAvHTd7Q7EB/
zI8o8HN7uemB2/J/7Pq/NsXQCnLHkf+qwPV8kaQBavbVOjSoMf4nPdLJE6V1Hqsy
JfutWffy087Xgr22q59PBUAVudhc/GkIJ4mnaITHyydbCvZMMB8YJPZy5kSnqVg4
p6htszTzeufrxknF5iEmTodbXIuYnDzxtk2m39i3OZuKySPf/aetLYWKYvEXohKP
98DQ5QARCk11IV4Z89q0loDnWv3/VqsP6dcxYn7vx51mQn97SGst6+1NUXa+A6Qx
W8BNRhtXIJbKBQq/EFIHJxnEc4G5rRtS0PdX7QHCTpfdKp2RbxuIdTcJ9vpaw9XK
qziv4XWeirBGBiEorWRGmGDmCrthVY8GZ9O6O+0i8FrLT9A+4DB2HNcOrmRq6VVH
nKv97xSk96RJ2nTBfTZRLuiOOUQzyMbgHF2u9iCooyszXBRjpC012FyyYwaaBiPs
QCLHltjPIrjiPwg7Ki2Wc8UlGVu3ULSu2PVM9HJR6nEPpoSDbcZCnlXIOaopaSTy
ORvFCN2GwapE1A9wNYSGTYdxZdIFrbLG060IkL5NdgTdlOzD/LPVf7iTtc4n7i2i
+7L3M9ftZu2lLdUNJ/Jt459V3VTPyD25dv8+zgJQLwVnae1AwasL6hupzypbwtc1
PTA1tD4JIuc8fo4MeQaIf69RoxZZf87NCdAFVjsIfNOWf48CtE8N0cLBOyKXZKSJ
JiKUt00mO0Fl4s2gpESABf+6s81s678tvPDL8oGpz9nZye/0wKnodK521detK8K6
qPyXQrO4sNtpoyF5M9j0B7Fhuz7WNCLIlGFLs+6Y0pA17m+BhXk6Dy8yITYpcniu
t9PLYf4IkMkUECN2kZM2cwHPD0U83zFxR1OVHhCIoifRAf0ZRO8B7d1eb/ByO5rw
j9YQiL3Elce9jDtvGOGrESakMEaX8RRpq530whb3qPbCFUDi+PsoCiDKkZzfeX0C
wwovAxn69qBgD+/T6oWhXjFy1L0nUEqacDrwqeKEaOjJ+U48CIZ0ecsEzxmFZHKw
C5zYtpZ4WY8FpBZ+vNYu2/x63uMqwNPLIyedLMwtpdO0joMxvrBeWO58jXQSmV6M
dhKzUwTdGqzCGzHLWcZIvYmZh32ZftoiEkmPO8obtUov3+zJNzUqLeYcfTwK9Y0G
m4TJC+CINRrFr7Otkyv+6eRsvvscw15IQV74XFU3TeiELyGiHZittI9TF/2OJcJo
VZvGwy8GW3gx1NmddG30EmQYHSj5IpBOW4T8SEHc035AGSwDFkUeA7yHN3pgH08y
3oUpd5uS+0X/0wmarwex8yC22WRYK1+5CMZFvnx/eGV75iYnZSVfijktdaCJ8PHG
93pujiVrak+VkRWeDbmqghgKAv4o5d+SukXSxbdTfSefCDLwhFZCPGCfIZTvF9mh
CNDn/GS8jvyUEUEjWHMH5ZGOSjKN3i7Sg04hqglz8FRAi+ucoAA/qIy2c1vaKrU9
KFfk07LZf8zGM+lv0mVNmmi2o/+BsceV/uHf7JTqVslvh7aNWN3Ik9KzFhogNJuD
Jj7vpx9Dl0KC3BZ6hpwAMs7wMB4QyEtPPaLcWbBxi35uM8RS+vSIBJqgPbybZIs1
SvdBtyCUj3LVcSZ6JbNgQFm18BSBkRG/1bntvo3x8fssNd8Z3l/bok1OMlXDwxbb
tCz20ANLwOgFtl438m2oucVZNAUT3Iu9EkUGkWXCKIaTMDg/i07U4XNu7MRQcKdb
mU6xXLbd6IkGwf6fFQCK4cDCKSekPzHGKF8W39qKdKARxhl5orCcNEQU3FLO9l6x
QzZomg4BLgmAUZLEOUL1cLCzao7ZcBtReMXofiPIR3YADJe3mOIOS8pt5docot3x
QQGLY84Y/xZrcemGTCSPB/ghaAgsLv9jyMkYsVUp3cTRnhjsejkBs62It2HT4FEF
pH/jB+ZgoDCTpy+mOY38PCdvMdxM5ZkoASSr/u5taREcjlbDlbOik22KZRmiGJ2j
xowML82IK8fmPeV/EW3wJnjh3HTjebq6dT0Rwb/z/g5laDYsSEPyoEthKAqFjNkC
rELNeLU6AgH9x3gIicfBsqFn4KvVjK4ETL/RMR/K35stLmZn7aJFljgwgFjISI52
Tvb3pym4grAB2EUPUZQNqRs55p1qYa4qABdGMgmiO7W2CDCvjhqtZk8BeZvszFVf
+M7xCESkpPutMk6+P2KbDc/rjs5QB0bmGveVkfJQSRZYECjui0bF7vx4VBX+C+qD
1JaSe46dTtJuAjVOaMwb9LHDwR7JY+d+Tnl9A2VBLo2/P+ZtZ6/iyUKTUcebplKH
Jo8zgDD9gZHz8JVSIcnT4o7tGyDInl+ll9y+Yr279pH2KAd9n+1+a7QXWlhzSh/A
iIrT2onIXt0kIRinsNUOJBD8ogZr5mJRRYlrpbehpFTjmrpf/gf/GhliHohghMIc
HAjYcjTuCkAbvXdgFVoL9dDGwM841peaZY3mvWl5eqfqtpwThvBYaf9vxcpRllBN
zNnqiq+ye+2OT9tWpo2rxsG5MIPb92qSVrCBsYFRqGJIxXTllvuL9jHwMekBpFks
osaRuTt7tU+P5Xa0Fa7wfbIXr+lxwJJrEURSt6+Tpi31BS7p9ze1dr7664IHQkkC
RQXh9wMMBU7QtwPUSoezb7qb5iBaGWd2aZ/e/ohw06XTyrdEfFjjapMrw/QVXuu8
4P7Q8G0QG8Qg6St7v5498ipVuDGaJyiLy56vHTOStdK4qT0QC3bR0Tkx3OcY/Ga8
Dp8AlJfUgxQHBpexaVpAY/LSUbPPkPvbH5/bmv4YA9ZrcY8Xbixs6/Jp8hM/tfr3
06Al9ukV57GH5673jtemqK233Mu3AJcvNdudDcqIk9MzR3+PXdKWv4cj0DiEPLMT
5hWPonR3PItHCOkIpaEUCiSpmdZFEpu3FlVRH3uEwW3slCpuz8Th+3kps0k/mnT8
wEkh0OECUO4jI56C8TBUd1I0JNHDaAvz5ETDkXor1ODkq+TNtAoRVvUU3r2m1FQ3
y00NDAlbt7jof/hwMVots70CMKNDhDgE6glG1VSGReQgoZqOnohNEtXIa+lwDhKr
ZVr6VAIIJdtVwyGNUsPFxsEdtttDYfstaYhVbG4Fjydhjin96LXtWiRg62x4wadX
9vbvUiMOcOTA0CxfO8U+6yS0w0ELKW4i+JBfDuWel42iwGo62NjXKEgMcaUpcWqW
Z4B2L/ZdEqF9OsOVEKWRfWd/Uwyy91c/37Saidb4OX72TjbHFU6sRwfQ1IgZRHdP
SibFmQ0oJVWzP9bq5xbRcvXlvTKCNnGWTLP1uAagzCzXzC62egpUDnOuDNmq7aLU
9YwCOIvexBdczW/iuT+V/rH0XQsdYOkt+n3S2Vzn7ctDlm9xbI7aCsWAn2Kv/NWn
u1iDGeOTa9bQD4SAL+ezJLeO844xOq5PCFyioNNqPQncu5NbIuXP69av2+CneEof
IkGTkG3QOxbThha4ZqYoi98zTGX8Et1NgTugf4fiPcup3fdADgMOX/93bSGKQHgh
clrA8gZ1hgb3R3AEGfBY2XMaVslvwr+jFlVOeqgVUQK5ApFBKdkNFbbrWw9AbbnO
5h9q5fCWmXyeBAxt2FA9kTTxXeAgxJzYpQROmZ2yU54RhuL42ARxyPF9oms27Sbm
3P2xr8NqwxxFTIttgrhcU7tCFvxpraFYaJeBjA+kzQzzV/ls/vYiWaa0tjKgMDHw
WgeGabgZhFN8P90/XynZsnhLYRn38Tu1D4t7hzePOaYdkWal2VZ9VFUoIw/MHNbo
O7SU+qb9fIQv7mbDAnl+TnLEIkgh8oitsqimLjzh7DpLu41Dm8Uog49sxyaXfyZb
4mmtSX0CWc+cA555LDtcIKvS0ZPBdswEqStgd3uj872GZ6yyJOdzfKNdI5mM98Ih
upR5Qf59usVT/Ia0X/gnu+3a5J3C7O22P17ypngG9ol+0WMvVAgrToXZ30kZnwc9
ji7izY7f43vfgtMRyQNWBJP9RtxY3IfiJ0VWMMcF/Bjmxpy6IjI7zhGt7VrsPe4V
NCX6ycb9GA6Jus4q2C5j/hvSpM+/4WmoUHrsD9pk3k7MOyQf41woEEYb8qik8waG
uriU2d1jvLpgWWMpkXLl3TNVZI0Ncqkf7oD0hZXse4zS35lHss9OBGNKaW1tPzFS
ppAc8hK3fbcBS28yZiHD/S3HJagk4hbecNrlV1FB09gv2RngaCCfII6IuAB+brlf
v6LLPB6WgJJItvvx7GAgWnE6v9Qr7N0hrxnP/zF0ocnvMO4HV/x7jdr7UUstyxs7
WSubQKdGs3QcET6zVL6mvO8Fsr8JazJb1rt+omBk3DxmhJvDGgM9h0tk8+1PJCwa
NutBdmtIVP98zzaGNTWsxVHQP7Zxcx/f4j0vjmkQ56bPv3oTR8hkxCCJx92tipfm
eaCQ2mVQtNVqgOzS7lhYekUHzhukl65NY31sQKycJ0X7+aIxWZJc4f14Tftz+9eQ
rhztKqSKjE9c1jrFM3esqvi9QUAyuT872F4+ueOalLutPxEsSA7QtayBCe6eiMYj
0Bx/V+xd7fL6/NgZmSf2wn5x96LxY/Q6xOVE7DVvpKktz7sICqWcAyVJO1ySbXDl
x1+RzdF2jUNTwJB4i6dnzGMrPSjEapCL0Nrcv9Ovm5eIpCPaPT4g5LuASCeP08tP
cSJkabgGgmrBXBI0NvA7Cfe2HtJfGIb6GoELqF2H0XuC36Q+/fgW10ycRuYvvrqR
ix5tQp2wqaYqhQnn1nvENdBdVzwbxrgTt0p5+y5mO5gjbC+PcTE1rFn2Z21UNeJu
n3CPtDYCijDltWxP5jfSrn6CcUNH2QVFQq+mrrvIrQChLRSZJDKf9ZeYkhEgeNEV
FxZSoBWNt3MtUTInH1v81q6cufztUl12ALbzT4g9PGETZ5zyTo1+oY91pEv2tM5/
INaIjJ6b0RbfN9Fe94UXJlCYin/TzzRVKX78GKQjhqrD02MmTM8zpM3PY/+sOJjn
zex1O3yIZwPvBVNz6wdYZua1Ypg+of+lY3V88Fy4IWK8N2f0ISbP74tMG1T3CiQE
QpLxzBEyK/m7T6OIubvT3mjHUVUNWPB9MEIUgBfOM0q5AGlGqqByMIm4D5Ejn9vs
2bApILMOtuil+PMVtZebnGkEHgMxIL3vEz7tjHb7hGvn3i3b99uNQSD1hAuPAbqM
Fwt8vtUSHR/juJIEA8Wams6yxiEBUmKuiU0nkBOpOorI+vtcwpkn75fW+Wmasctd
bHZc1mqcy+b5/i/7q37mKhThUuwdFewUkuYW0sTbWf2k8xZbwCDGQXf6DMJydw28
zspy0PtmFbeszXLwMNxAT5zQAz2FEeCsh8ytaneVn6ysD6ahmG1GvFFEKTXJnt2I
bHphENZ+fttD/FQ1blki2Ud4B6RPbNUSY8q+TEgD7uT+BvqMrEmGq/Z5hw9W60gR
4hYRStfizgNDfX/Tid2tHzfp0tm+aOLNqzctxgMJk/+qI6UqVuBGloywQOi5rKgw
QLj1FciTuJ0jSwst9YfRJXB/oChjnoMF2Y40SWyno88m03kiXgSYmxE7Hc6RtVy/
gCvBaCDDUwxg/IQSqzfQgtIjhYaoJX4WbAs4sR+cMNUwKh8lgfpwC56EDuY4k5ha
KhGQWGbvyjP7Mo0xvpKuM3CiYTrEhDF5nbuC3vhs8qh2aP7/SvHqHOGMzom2CUSH
LtTxLh9gQDbgZSM1lw3R5frqiPq+2DZXSmtLQcCzmtVZ5UkZEAcrqCKDy16WKcna
tchdximBbJRH3G2PpKcRcJja40ZJXiojjnQTiQvHXi9TWvTrYjvsAokYZzHBugWD
eFITnwOm1MFEQ48DLyUa0J237+MGoayy6RkZniEIjLb84We+hiEMAfUmYjdNZkTw
8+67lZ8YSHzjH2v+R1Vuoxz/cG9VPre8SuEuH9M+Cyj3nm65cIcgdUcKPLlPXqAW
/CZT5a5/b75suKSPC2jpXvWRPIJgtjRMZatrxL15T4ou+b6B8BThxDyyIQPymG95
LsbmIPfvop7xA6thXLAzwtchQnJzAuaXIPZSmWSmRV7M8yniaU8HRpLPKHQ7GrZV
ahmBkp4W3pVd1xts6f597DJXCezJOdPayG2wPWjlfrub4ANCKBSA/CyqtX+Ewu2O
4Dv+nZxqOD+bUjAzoXqwv4Y3qf1ZxsUNIiWDLbFFib6qPzvqaOiVhkMRJnkZKuDb
sHJGFYq7dR8LIzJ8Si4TFrsOzztxANicAIu28gK/oonNrJQZlkELGwWm6SFqKxAg
0sLsU4zEKtAoXLYMNzASqLfjwYx1idpMNJfTWkvc8TktO1QSGiDNA8VHSG81kiS4
WZi/aoQotv4BFTVeaQhTKyVHaEQd8rE92/Xc3vCCFxG+DLQhNUhkkmgpK40W0fU+
l6iW1CVHQr6lx8Oore99kHE7nf2cLiNVlPuoKYh6MevSCZjfW691XmYuVW/yXJEK
5qCGjbRjWhjelLJUS2xP5buy11odEt2TZ16bq49UJ6avyhOkOVSV2dWhPoX7vwpc
3X8lp4yfT86JsoPHmjkYwnjrj4I0bc66WRNVzULDYOfN5awX/V0G02C4VbLD1CHW
8GUeJqON3RCpQrrRvkTe5NLO9hLoe54DRUK/tv+mg/XHFKSCGV4/O8YNrsxmLdT0
lhnjg1xUe6dMG3IG03VjE4Lef7C+HshZeZZVhqB3M9DiGWQb7X9/k53rT+LCNST7
MhK1C2ozl3nSEkyLG51nZzdTcp3CNR/gv+N9xaUIM5nLc26HfAfojg8iu90MHBlX
6/Zj5FkDdrV38LXYN4EhzJveyLD0fApbpyOcoBuPmoZIImVPVvKybrC2dbli+4H+
yfji4+adAUa+GKaEWUU1AEVOUVQscu4QG2Oy5yCha+n7fkzJDNPqCQLc7BT3tqfW
seyw71qqk15oktWm2Hhhbdr/SSKfSlTypGaANYIX7yLzBvYf7rknawF7d5XfN7Wz
Jwey0M3UAajYT/lB8TQpkTHWhtZof3uEvvxZUwTUmEbZUzKCYrMjg7rhtjkAnHuk
azVeBS/zaz5SrQXbhfMvu67DmIYDi7/wHw28i8J2U7/5xtXGnzHXnXdQzZBd3Sqo
l1Wt1irOALnxc3vABPVhkrnYlUEEErhecqEwUlD0r4w75CNjx3myJPV5FXHLY5o6
LCJcaadfwTU5V56ptR/QyXIhUm96mrC5ivqwCY2zzaQ+WxEOtQlF1KCsCWw4j4/l
ARYRpWgxBtTEDTzduMK7Zz6Cbuf/RlmUpjavoO0U3mqOZb6fPpcD1WyEj0ujsUmA
7VYq5PgL8GZveFJ/nM4ddd+6yr+rOv9sZbuRNh0WEkhCJObvu9yYOIsaa50Ji2lJ
S2Tcx2SyDa11FBkMnHn1qXfcbuAAqdlmaMwsygJH/ZmQ6j+S9CT5qpUZvcgWiVsN
mzAXTYEdMslyNHvvzGF5gtk1HTJKiSy6kdOQ4GiITVU1kczfMgAPRceTGpPmCARB
Tude1tX3NDn2jgjGFSqJLt6gpGPgBSQyBFLlcyyMZi2yZOYorrCMnvW7rorBkwdE
HzlAhRAj7VflcCWNkRyCvvlVkC/wniYCWZRIjB6ByyUGZPcSrHgo2cywMP8hRSUf
+N7jPIoVr/7y0JSFMHh2qGJv8hRna8zs5+d+ZplsyTXA3vAzt+77PRg1GXLse7G/
TjLs0przp8mGReLBKF+tOsv0IQDPmAyk877EuUulZiPkec0LNG4YUcOizEcau4fF
paT8onzhMwRJOFR+UifPXbqTe/ql5FK+gIytbU3rsEG6Wh8uIQW+fkw/NGdAnplN
9C8eriMppbtshEu7IKb8zLNT3hta1z/nKVJlt/nKuma7qJGep2sQYTeMZ65vUvAD
iaZGC16OWEkmyWKtLl8KzI5aW+jipKwUZ+r6ZdiSK3SgulcAMRngYReq27XmQjRf
IPZ+mRWoUnuTvviAOpxHqLkl0kjo5vBeIuZqFz24iVYoiRnfvNuJ2G+4tgj/CekX
KicZg7Ea1JpcmReuAWkL6pTAG0Sv2duUv93hxBjJNZ6uPvJMp9oVcX4wH5gc09Wh
YFAsMKhli4AyFTXDJgu4We15xiB+ZPbxSuxYrDF/7X8/xBok+T3B7XzgQroHCHo5
BMOlurcHoQNZDKhmcWmWT/A0jvJIPNxTStIgg9oKAon/VVIbgwA8fYwfKzrF/MDK
C2113pfdD08+5o9fvpnBDfp2KKJz2wAgB9793bKRZW391IozRVLqiVKftHa5uoL1
iFxLrN0EmMapaPnzvWeqA8f4KHNKlKnWf3xlNwEiNIsrxymmcCpxJQP9FoVs39HR
7YifWmG928/kzu1rXtBIiR5wl4LH6GFRVEzkC+hSXDu1aUiPxFQD0GQi3dFd3Usl
mlpyyXOuRCYhHQm+8Hl3tEQGb2nw3I6WxCEyso4yP4u5u20ykxcaiXc/lDCzHR6s
fb3FExbhUgpdIgFXsADyhM58G5qkKur48ZeEoFqsi8owA9haMb86FF3SyYt47TnB
S8ZD+k6e4RVCjEaWuKxgRGFyA+lWeS3zuHXh24+M1BSUwVcPaqDAn1KqaPo+jCnu
a47oIbXVyhSdUhBDKUMpWOHKSQ96fpj0QLuJ8SRlyanb2VCL1309tWIrD9IAVdnY
29t6xkM7XikiPJeP3ZnjXaPUeC/GoWXVL26b+FX74FuiB/P+nBrTzk4P0KkzbUcY
8Y/oEkUjUmmYPtwny9bMqtKircnCEVjouLclKhYJ2r6XlAGUIyeDUxeb0ON4fhfz
+ZQhj3EFHfTdCA77rCBdgs7UlKLd+YPWU/RXZEw8xDfVEucPlL08+l8+RGea3stx
/dZNfXv/P5nD01/gwKwMN3NL0mZlg2BCFS6qHkI+h9XAvowryKk8AqowhbR2i9Kr
VSGNC/rDprn6j0Jn0je7p5zBFcPSab3eEKVwVXOg1R4Kah6xJEhglSGvhKZRr/+9
pkHVJ2hyz97sz2PNdfHrJi0uZXyEZXYJ0P96h5SjMLy1UHocInC3mJk/Y5h8wjm1
2rCtx7QgtSL/sCXap/btwTTiQL8geQlsF1yr/4eGiPWbynlyBeU+BAy9BXWctvgy
HSBV4Yr2z1yBjK9pA7lrX1fR+HVNayzJEXu5/EFSX09cyOWQ2MOn4A6lc3MW42Nf
V1+G0+GUw5M0Bza5paBtJsCd361pfI/IN6RwfgyEqqnNmjT/G5Lg9YJk1Ur6ioS3
wdpCt0wq6hKiqBCG2AeBOlCfF2LdowLNE2wCgOv/yb6JCdkSwcGKGEGmBFnx9sVm
01IUd2jEoTc7qj7q/2VL9a0QeGdzdkHZvOnJDmHwftwQBnydgO/opv7RlGRQkwbS
H9fno8zO5mb3ymnyfyKHTC4M9AvLOtBzLS4JVez55rD7avhu0HPPu/e9Bmrjwk6u
bcRNL9Rgd9jTo8xJ9BLbXQDgzj/eI0h13hwzGQ6JN6hv41qKaZBW8HXDGH9gVEmA
rWO741h5Nnh1Hz/CwCucAXXtUZ7V76Mpw4I+T0/dj9TO7pu8ydd3BJ57FDcU0X2F
Y3zLCuxphcj98dOYMwBWoBPQVUt9YjNbczCYVDF/Hr3IFdmLz2yGQVMTYa6EB9ZC
lefvUQ42mX/ixsv24BeeoCbPBhrLHo101W03lqhvF7Daubvbm8cHApLAqB71ItYh
fFhu0nXLV8oFt3GkKpiblnFaUYHwFYpaSove9VL9o57nqfOH7f5xh84mHSYumvSH
s1qL1ydhLAeREBCv9jL0d9a+6YZ2Y8YOwR9isnA9nJnfwQu93TvRV/W97MZeF5kG
c0NFNIeGTATzX/9Wjzrom0sKXU1SpNGHxi1xlhdAWk6zDvkm75csqOqGmWEC0hD5
5LrDdV9uRR2vuU3Pqt9QuUZ1ZhZtF/LubtuDIiHuUwuGhl1Clg3BhboVMUoBLN3W
Ojft7psgbk6G+2CmASEVuHn59a2f4TGOH6Q4DhTz29EcDhqDgOHmWmQ+fPWHGK3s
dH4yEp8Oh40GeIwNYiPSaIpZJ4+rk606S4oRPAcK5EiBHMF3d6NOYIW3eGdqrnyJ
GfRWgZm0k8P1tQ9ojbnpdyZpYwuAOL5ZEZ3qNNF5juPHAmGA4sYHKZpuOL8YZpfx
8SQ9pzPIcxWjLyMbHLCISIQiSSogxLWZ05xnpgYVG6MWFPsK+7OSK0IFr64EKOgI
Z2jhkdLywQKxKYkJrn+lbrj0YqEIRZ7lDapbr9cR79QFbsxJWiVJ+vh+MIWYxzpQ
eWKcHIV1asEQT9u4CERrPC9tuAk5vFyOGV1zDaP8aHZP+PGBXyFcE3+igoNmOgIR
cKQROS9yisZaU4poLef1UfIxgHiLNDfYyynIr8fiZpsFfwzRIGiYea747+joeoTq
4iIAc+EOR9iA4l/g15CCB1DtesxITMcIfbifpH34tedYS/t+CqIIE6WulICXj/b5
ZylcLAomlr8eRTZ/WYWIybXBQBTSmf7MHLrqMUd7V7EFbFEy2XMSx1Z9NSbvKzMy
z3qzPAZMc1GVla4/6FxF2U2iWI7H1E01C2pEf6IOsBgdPORyyJaz21JGFdDxNTtJ
wVyY5RI8tp8w2+Bd9vfU0Ao2YrlV9qr54oVLZIxRy3v0W8gWeA1QP9BuyezObYtZ
WWQ9+P5bvoI0vJKluNxkwoaM4VQRxo572GwYbYH95IqySQMVT9reCrroZ9mDZEDM
1cbKflcozc42lnvYOzfZx0K//YvBIs5axZjmzqDgf2xvnwgR1pX5Zd+4Cd1P9fnN
mbiAsIEiSxAcZmCnCs03piw60FlFBpuc6fzc+h9Fj3pAeTzUs6uUBInrNZZfFBZV
fjsTjehSIieikBPRPvq5stlxAMxpmVDb8ivA0dah22YRtkyM1OwxqXej2kdTOu0i
6wFapg8ExiryPgkse4qkJcURsPO34EwysuPP5kQJxXsvyGdNSHf1s5TxrBmOXi83
0ny/OkNHrlmNI/lKgjP1bm0L8xBeuocLDmAeo4M8JCrr+i+Uj7EiZbcO4elqdhWb
XYpVx5b9iFqtLuhSZFmAihaYXXe/OWKAdSfUfasmUGClrlbYKblEtCtEUQp3GzCG
H/G4FdGfn/hJMlCtoSMv0odRcglWdh5S+YyqO8ghdXGUnx2G9nhteQpumh7iApQ0
NVMvIvjTdT7Z0qXmA20jCxY4n56gefXvHKaEnKjwr7iSraFLzQKrU6eqshP+3bQc
uDR3GEIoAwDXsnRgDruaXViE7ykWyquPCT0o0807LxXm1eClwuJi9QcaAaJexeQr
4Y5rPjt5DZ23twdMbDNMelztvRt7H7pDyos96AQy/aTGbPTv82d/T6QxvnrYxxSk
lDDZ4ATlVI580J0a7x/SUac/D55bfLQBJOqcuJioGskQqluKxe8yPkQHx8thw4nF
TaF4vdH+U7h30Mfmnhbt+AmnHasq+ImHPOeA2GPNOaJdt4zUi2UuX6clieAzj67z
YBBOv7KjNQYFHiZRHkZeM6Ebl2rjShTLD+hs/9bEo6v5DFrbUjX5672C0BnixBuc
GBoDIzM2pL8zbbvhwFiLc4CIrVSUawzxuBOOgVRWTBPx5CCKziYA4f/bgRTrFign
yIqz8HR8cWe43OuADAwemwfLSozGvo1I8g+bPLEW1OiHG24o5JRioheW2nUn4v3F
gBayDY+xhL4KTRv6EBtPJAI+AyvUqzRm6v4jm7aprOfpbQo8Td74FDijZvIRVt3y
ZQoPArCYj+1mXWHiOz2G7VBKl6FsNg8ysdpmf0IGfPeULkg2AaMS0srXD5RupCON
wb0t9Pd/Ljj0b5zB6esC1tT+FMC/tVu5XwTk5XWSfns5+3PBoDZ7bwZ/9R9LtsW2
ZNniz31UrvpWWHeLeEk8a3dVhKUWDvoCo0cRfb/y2NQ+eVDvnp8jvEL9Kq7UsoLE
L9lfMGuXRJ2duzqRqSUDiTNIPp0z9KTyqksbnYpNIDwGH+5/JlUef0nbe7+WdH7Y
BQCZl+Kw3TrrXC0M1ywhoLhHkCJD/e8VqL6fnjeusuXGdmgoQGKgSr/coZTlqnUa
7wu3SuIzDNMtI7OGVXJefC+n5P+0g92WTabc9JdR9joJXmK3HR+yZOncme41ZnAd
wKRnysAcVLPPbXKwkk8EUqgqP5byCNi5zubvvSKC0DInDMCcBc0zzg4z3BaIH4jh
prP08tulXlCay/c27xoVyAVuDeczxxazaPlfo59Smr9smvC4SqDeK9oE/PkENy4V
zFOQ6pmltvfs2rOJbHU6tu/jd+V9GwO9cWVti0Q5uLEGtmxZ6yVp0oRSX0p14IEz
N7Dmi4hzTRZzQZALmlYB7+XLRiqucU95vepCFQKig40GIUT72KH0gOXDOmFYPJ9D
SQ++dCt0z16YWDUHURr97goRZXjeIlV/VZSxFirLYKI/mhvhhQu3DXDyz6GozPYr
pyg9ngha5OkpB4N5JyJeNr43EMcxCNBgL/KP6LZjxpZlcTbqJNJSqRafl//ptqE9
sNV34LTJAaldQsPUMonl0/VwtOis9XIA8mElgQGWJ0zpac/4W8Tv3cCpHOkUFFo6
thlfsFSrx1UxPf9i74d6ZJTENNCHEl8iO95LGUNqNT3s2XcEi4NYhBCQhRmAd8rw
v+bu6JQE5N/0v2ahMnz3P67LxFh4g0J/j00mRNGHo8ACAOajQ8K9RUfGrH0+OcKt
IgLylBdTC8NOVcH4mmGDRsZw6w/li/65vu/vtq0oYH+MCbb32YzbPAJAWMUMq98+
tEMu2WbieQQZ6jkQTX9BJYEI43s/PLsdLry5SNA4gWA6tErrzH7RDB0LR++FevwE
cR6yHTUgrHJgMxBpM3JzccKDCHiWcNAv04kN8NhBQzdObDWaXUdCJ99FnEnyWshS
zSA57NW3eRi3u4Z2K3s0Bdjs14cxpQ2n3SP6pQhWyaBAheqNxK3xy7s3xIYdbVe/
S+mrvsz1da1OvSb12rA0fymjoRkNAnTRwZk1C2wQMogFht57NYo1508EtcgFfC/Z
2uYenS+lu2o/Hap+ux9W8D6UhYuXj4kTJbKQR7/t60E4k7IwxxWgfQS1YWL82TI1
2MV1NVfrzG8OVjiii3XRLllGChST+Ht4Vw72zetcwlaBVMPvKSgKd4Q/iWxvKWzX
Zju93ba66nSSw1yJ/yDDqxx4BJdKtYU+s0KiY2Dm+HlpTG5gpN9lmtD6jrNQX1Rl
bTqMNdp1cXXFp51Arh2QIH6c04ruG0QqmTq+g02xFQTdHAhV5kUjbkWGRQj2bFlV
glevo4lcjivEKqsMBuQHQwo5R0+bF9+NEJLAxeBMmT/q8lH/zZj/fDIY6lrjAOho
tJxEckIvporm88UsoKLflPYjutrg19QnoogVfUi/DemOFIHVxWDdQTBwUNt41C+Y
tbukDsF7SG0st9yG70/AjToWP+6dcrMPbNVcFoX2jYWEIQAoeoMMXef4RqVaZeRU
CEXc4Ulluif3St8MlT5UlBtfjMpfHzkJPI5wdKEkJ+IZLWSfac9C4L1JLaf/jURB
JONmddElD75F08KBzhnKvKX+kt9Qr4c4pXuznsE2zTW1Bmmv+3txHyLJQpJCRU4a
eCqwl1TXJ5gDH3XYOQhLk9xfn9P/kDm19xELYwxT+Hw9rahU2iEhh1GNGF8yp0SP
IR6+rmBq2GMxVdEshWKJfgL2vp3FMIJn0sR0gkbJwBhxP2Dfm8mqIY0jcF5D3JBa
t2U1dgoKvAkEQoxNQO0HyHWULO5Ntt1IBEY+edcANdbxMikRH8Z8hLoWWHGxZuqN
drXBP2MESbIALR7WaIU8RIaV1w/DTKZMfq6wcnTOKKwI6T1HYM5FszQvsaheG/mi
ODhSw9aJr6RX+qJkFOAUB9v5zMdhPt4ZX/yHa1VUHIYutG0rtcsx+QVcJWqCoAGo
b2Hh2EEoAXtjHWG+u/QaN3Y28Jx9otxhzcMySipWNPpqGqtsHcUfSDzyp1L2jeNc
mNZy4GrbWYcTXl7F8UQzcWQlgu+g/zj2KesoaxZW2RkMMUrk7VBkdL4Zdw9iJRr9
7ZPApsD32pEuAjt6RCPNlNU8JTvhqYUbaisKM9VCszFT8y4/s3fQDS/1yTJBhmbT
WXNuHluKLQ4SFXo3C3xPNSRxCTHtMj2nSvn4yYJrbNw/ZfIzvM225W6Kp/gUSJwk
WHBEpB9fHMpVlUxKKJ8IBQ6gd1XEmmm7RnZpTbUaCNqBiGbvwVADr0VjdKqrWF7r
mHQCZAQw4t32CGcEqyF6977Vveer16fr6i2Gi9VWJ1st/m0v4Ec69AXRMCebtfMK
mLsR32nqelK0PgEcGVwPE5S7E3r79fT/AxdFX2scB3Txhu/ANvuO4XsIbeO/caYg
TDtdf8GKY31F5d4izB1jSoiCxkiefRnihEeoRg7+kps/SeMU3ZsgxyryP0C5+bpi
LCLgIcoG7iWevAmMwtBGmkrcTZb5dOVQi7eH0fK+DDh6QHSSW6cljiVZ3ucgw7Yz
+GO9fJ4/E0CecOCBn4/tc3xkb4bAJDvdscMHdD0jGDm1ewD2tzTpHxkIm5DsNljL
aZjmYLYRylaXy7PVCBOyqpqODWStKlT7ya7zmC5v5M+E97sgDUbCnfs3FTwRSLhv
8J4F7X5huhmhYGUQdNW0ycIj9vz3xYXP8lLTMkEkvlVY5s74H3W6iPG2cjA8O63t
o719aFjqDQQL8W9g5IDE8QWDOnz7pnbC65N4567AGpme818fUTiaSV6KSnIk2X+l
F2mVEzw6NhAiE+efBBo1G7ipt2NNXLa8Ddj1cKJzlR/bitf2Nzer07q7gSBI+ces
oZasSWamoNVq1fhhB+ppQuKguCNoK6FEuEA6/Qc662peIjI89FlEK6iDb8UjRoIU
SHHbKBBP36p3/XofzHSLsMPjfhv8EhPUmm5CUYo5twn7QbRgNlpfdTaJyw0i5cFl
cpDGB3+WE7wQ2X8gOZ5F4Iz/B5/+ozA93pIIq2ZAh59LYW9kK87prMS7NSU4s6Lu
r8VxmHxKDczRzlFXTM6qKUlIKS6uZmpB7k/h2X3euCEPSkLNbjL6hFVkIEaIJcyD
35TuT66ObyI3DSisers9wO4QzIpCXGuk3FKqvuHxpeAFLJEk5gLFDdBRk9AlQGSV
E0o5pEoVys0hbtd8IqJeE69kwuPeCU2mj5GNoK8F8igLyf72fyLtFzDS67QBH1n4
L0sdV6kA7vS+htEj94WnKd+WzE0FXmVszmCOyMtLYXStzrkdregT3xz5jAdcq73G
FM0nSZQU2crGG0trQOeNtowfBsQQlkPhXx0SkK5C1vIbqvI2lWE/vi681mq3wXL7
l/leE8Olqb7Czudk2F+BgaU0mUioPS/PuVl2aT7FC3KU5F8ZYW4fUzswY+poXWG/
UdbV/TiZUeTxAz75BMdfD+xrnSRwwv5cm1HVj3P+eW7lUbV/4AXP4DnzUKn34Keh
SJR/oOfg0NExXviTweEcZfaOgYdHkxyszPbMJDzZb7eayHq3WYAZkuI0DZ+spYYe
6yRxom5ycZNzIyvW2Tz2bXaYACN534EyN9VhXiGLdP0P5RwHbWZgvAfaw5V4Rmel
FoXA+jHeaJjGdNFfZjrnhW7AvwDBQXZo3YznollRhRWf1VSHy9Y7PNMjP3UhNmNk
qndiyszrvys5ebyIvGrKhOFH2bnUp4heRie2Mdp+jNrBS7EARD9540/fYJYh1WS+
WLeOXhheOpN4VbGDg448XzBbbohwhdbjS+RTwFOPp47TrJCBLzBbkq4i+sCVN+7a
USwSlCD/SnVqgdM2KA/bKUHFJx8oaesq+4YKfVfjahxhkVIPrkWsES2dwxMz4dn0
kZWIf5mNGmzgjhg4YPvNbCrHdSFt1+quivfHdI9AwxZwpddaPYoIux4NkBoQa40G
btR9RABAyv7UQZdsX5s1fmDbXEH/PbK635xl+unonzSxbNery+uA3WolnJ2zXtJV
o+yRHiUUg4zkPz6qpXNGsWlBFJlR08Bul/nOWRzjximygxBQdHH4mVmMdl/UfBgP
Yv3qAdwF3NXfIzu47eSuapQrCoIkTJ5GzMH+DGKQqiMuummu5gXImImLIVrKnmdy
MCz4iOqyjOmJ0Gy/Thx0oSMsLked2F5qGswdq2FIX8Rv4323rek6CkpvaKlDHBcQ
OJJHbJYatiZ9cELBRK6cTWHP0F13OzIcdrwp3fxltTUGXC0nKT9XXAKKqoxrSmYr
bgRuYb21boL5bR6UloRar7MYU0fEYNFLsWMpHMHKhxXFRhC6J+/mk0UzQqMK7JgC
/HGKYfCqijOdFGy+69beXaJmQUCnsB80kAJJGcG7/chKl7/IPwjl2t1FxSOvd/aj
f5w+h1pt7lQsit/hM5OJqPOGvzFq3D15Q1iU51lD5OBOnXD/3ZU0fnQrdpOeKjVZ
KJk4svhf5lVNd0WJun4U2v9mx/apBL7ok0EMhd7OiTi94AbAigABqwuBKUjwuAZ2
zcPi3o/qq5QLZU3D9VxagNXvBBcPdhx+u+Oi+kFVxbLU27/tubunWMLzWXcYAvCi
VrzP63Um1WAnytdi0plrOe0KUhFThZZOfwmpuge6zbQmOle2U7GsvPQO1gPjISCJ
Lv5z0Tx/SNFVHimimnLIpaUVX+O428hsciTgxmOh/VkGDMktarQQABL3TeecXwhb
0gnL9/tEAv5FeyYo5YayCfdTRwOxVmURfK/N6FIar75uGx1JnyhTQfleUAxyLZNB
Ho2DwNToydj51HOd4PC+poRl7+HljE1vJDF4AQ1wu6hLBGnIOrF143Uxlej5Wawc
0CGGsi16CTXLDECnfccqK1gVQPQ1xqH1ANKJobsaeM362eYJYnJcilzgZnOllwcN
PQX1Gc6QfF5xdLNWwHcoA+nTU7rl1oAyBAbBTLWabnJn0QcNz9ueNMtHzZJS111h
niwdKUAIO0Q16pFE6dLaVrbIzeLXV5DYWkU71DVZvzGufsC/zZvgVFP1g8pBUBNB
w8/axGGhtFaLWJLCLd93OBGmTMUP9v00WBDx4OWRhBVCuaDjNdyj4NYIj2iRLiXN
hia2Ug2te1MyE1Pt3Wxja7lHv6sbPvkdmyGufp+GPmpzpL0uKKSF/VpPccwgn1+W
HAGZ9e49ZRLoG4TqjpUgAk2pZ+/E/vFQzLEFivecFa4O4fB/ZEY97xRM/WUAcgeD
7BPnT8rBBx7CvPF7Od8jQLkfMybyxlo1mZi2JEhnJjxNqC2Cl7m0Q01hf1VfAooH
Nfba3X70p7Cxw4CQvd1GfY1yTAB0TAoDqJ0UPs6YWEzlGtM8KqA2eM2bofBx2znn
cIa630rbVNupyUyeDy+LNGFlOJ7+nshvz/6fPk+MdgKGLGwI5oo2Sb42cHYd6Q5I
zDnV3+NbahkVmVnWjeYq9UKIsXd0vuJCNbZY8j2e/S/AyhgYHUOc4fBEtipyzg3c
fHGOfYFU7anJ0uQVlSWGL1fB1Fp1V9GptFtnOKkj4pZ/j5ikpN4nADv5ytLrzGem
iEbG51gYSsHILL3LBxy9SgWoype5G9e/gm35+XyXQU+OLvmjctXv+SjnkmU9Pmof
UTVfRJ4oMefySZI0LctQ/nudxmSxOK3nAvLlLOXzcPYdn2fkwRt3VkopCiKjSvp3
SS44Jq7zXdHOyXPVcs3CR5At5AY9FataTYd/lOPUcKm35vMATjUmhWrvWMC2Ucpq
pYaSNJbbdIWhQpIzuyuUYkL0OPUn8gtxwXGudzQSOphbwRzSSQd11DFDVFNP26JV
s26BIthxOxyh0ZGFrvy4J/8rujWCsZ6yIZNxS+pQNton0JFGVaSNBbRCond7nOb3
Zk13J17mbMZ/5oFu646SYU8K0RN2fCCUxEapoQtW4tH9Z+QduF3yOov8LK5TkC4X
lgPIK6H9/KDjrw3op4QlmD0V0OnwOYpmAc0PzqaTi7qMITgKoQnAvP+EBHzqF5Zn
gvwSkWn6WrAlqOC1G7UTKHtY53XRGPK1O1zA51eNemI1ArNlcEarw2IgJiwg0GvQ
0Nk3T5vXHouy7ytjMkzGvNsuAkYfWdbt4vGoF0j2CsYcRyEfxnrooBio8hXcStAd
HAr5Y84wjQZ9x03XB9i/cVGmEviiDcjlPsYpkv9ZFXWfC6OAQ5fgDL7qzlxOYhB3
mijbwtKA/xf1LwThCcYejg8zGUManpEKKjOJ4kOypKzAAdb6O/RyJHxDL69nzWeN
fDfVNfWdtKUXFU+veAv1LPQRKJaDMr9QpSql0E0R1Kwsm4cCeVQRazKRJpz87AxH
lfarKcnPowMD3ES5zvfrVXXYpxjL1ZHw0YG483FdGkP4tJ6/Ua+E2NXu6VklEODB
ceSRLwXA+msBwrJuTGU1DJYvAz1EtJmX/Fyc3mynALIEduQEsZRGbU3B3/RhKoUb
XGjr5ZOyLyChEVsnlaSWRkfwnEvLL6RtjI80WlPyMynju5pxoEnNz1Hl9QkO3D6o
YVugE8wyMLe9kckbR47m51S4gRJiXlzl2QcwxBJS24On7Pekd+PuwvaZupvF1+SV
B84f4meZbqabAce7Oa1qdz7OZMmlJgy4JRWIe3SidamuretHS7lJhZOSUtSACKOS
XEk4ciE7y8j1yXVJ6mAe+XiK581c4dE3ZR7UCFqO/Uf7VC6afHktILSJws97mHA+
Z5bTB9/xLP0t25a7mtq4i+VQCa7vOBO3FMYxAg0qQk7QtBoWIjjVhfPxkS8LT9WR
WB7sNSQWchuBhYi9sUpN1VUuFyuKTTm7H5hb37NdMyHqmtMVCpO2Y3R+R3obOygJ
B4lAzTpwiGE8QjiPc36wz2WTiV/3rubSzA1C/yfbiKdAueD311SDeh1aKQuZ0Yvd
E5hs6cUgLk2iog1VciChb//N0EoYr1e6pcuWacsDYTEtoJ2VYJba+1zdBsg1AjGM
O2Tddb5ZZ2BFbVB8oRCOPe6s1eLZ1vWMeHOjI597pPg9fDrRr0ucGsmwc0cZDWnk
UveCLboYolDvvcRcUJyyGrlXzurstiokAGM1dppjQV9lQ0rBKcPR7Dsuxg4S9Tgb
t0bQbmabdkNHb4mQcXUIrqEaEI253a79CR3GxcZ+XigwyyPRUZnJSycxshvmCSBu
bsEyYNsnMdRKh5d98V/NkY42jf3WTxrq2EJxJOr20psauEvAfzbC2CnfmF9XsZJN
ShQ7RGfV+ZpvFxzcetv+DWtfZSDtexCHbeBkzaXtjujcZ6TsbdpRPGksBB3MOhko
HqvM6zvESaa6IKkzLenH9iIhB69U3JvGwtq88lolSwPA+v/3jtiHXEDBnZqahOjh
ky4+cyzvrS1cMfKuB7BkvpRLgBn7AdaaM41dhSuZjsZQnSajiIck2XaE0C6Q3mgZ
lm+TnxhoQdvL9bk9jWI2GTqgywVzNSbquOUI6YDok84yrVQCOCtwd7ZCtM7FZ5lS
mp7iVIxDj78bpIQml5tE+i1kii0UjME9p8JkDtYFSf0gSrgukFaZBmFX54JIUswO
yRH7A7J1yK815KI9NaXtiTOcu7xqtE+kXwQESA2jkI/pzuhZE05Ui8xm1huQgVEV
l7aJHJ4SCMZcn/G92oEUkCKeEAKFGb7DxjG+KK72iuoNAFInFAsX5uA4fM5udDrU
ADA8B7iEJxAjIeVKFFwkQ7RaY5dQDQf39a9BKQoHShMIs1W0n90A6MO7AJ+v9Yf6
w6yOB9vCeSCgFroP1GG0HPZ9Gc3+Dv57d3YsB97FCNV6F/DGeBWbDD1yqRl9nB/+
iaq2XXQyJCmBwpEe9Y3JRo2rB5TMzl5kxo0KveeeOJrhMGf70HoHfnyOYYmn+Sp8
dOoBGvnraY4dIZCnX4HierU23E36T/xQVKyBhTwYvgOJJSksvYXoK5AZ1hyW3juN
acUCdjL1DHWhdM3lPv35JkktsEu/NZk4+/wvyYQa4D3DjZ0rsqOBV9B4GIZZYh7n
RbZbgGTbnhX3DE1BF65o3UygStj8n4vRmkUXJbE43Nm8uLAbGDI4YB3tbU65KGgj
zaYm/7Ojg2PZ0Ay5ZQkGQ1cWcZ7pOGNLnUQNSXX50kR2/wKzCulJFzGoKss7/w9J
nRY72ALnlKl//DaYAYOmwbrPkiQGqezqstQrdOauDijrfU5GuGF3Z7cxZ4ShXM5C
2EjEMjfy/shO8JY48chmKEnQxAGVygB2m08po3pGnKBgMQXqJv0V5IhVN/8NM/QL
zucIBOdEpuHr5xbh6wErVARiNDD2y6i9+XHpXdVZ0gPSukbCujzjKOI0Uehq3Aun
wwe/NSzosAyxLRM66XiPBfo3tDT1cVdh84wDRF9dA4LxabYSVEiCpq7cQkduXL/E
vnWj2Zbfd+W1pnB8hfPjWpp375y6dp6XPuSIAtVO4USJOrVITh+PQH6bgJW8YFuc
7AfWuHyhGMXjfp1TAG4Vo4eyqJ7OKA+CjhtfMFJGsoYa5CQUx+dehFmr3ucVOWUz
wHUiSxB7IMIJhki7QrFFqs3ofea9uXoZkgM/h0/pfEZoxklp1S9eBmnBSSsfUZ4h
9sek3qFvBMajX0wKbFupdCcHWtVtfUYc3s9y13wu8Ad9MkL7mu7cDRvKT/Vxsp/7
1PH22n7Uqtfar/+W5UgNPpPmdelsmileqKDNMSJ1iocIfXDz8feSx7abN+jrBvAZ
4IZnMkdRMhhOPKzgCbSg7mqM37Kn+MtVwIju1qAIMwGHUBEHxktYsvUHG8YuAqRF
vNGabIkzMcUPa6m5RKwlFaZjnaXE5CwvPyaG2LU0APhLxcMIH3Q54+htltWgkU3o
WlqDHO5lLYE0y6GbEnt7AjqinPbUVKjP+uuDrblDH2smeijpfE+4sFgnb5+S9kat
m/Cb/us0DLTEhP2sIugc0c+kN82hAXmlsb4y66wQ08Br3sKSIWPeQbJKXEflUMiE
l46CImqMg9C39yuOV5Ie6mfYz6uvSzMag7/DqxJj4AY+HE+1ZYDqj4SoEF6iX+GX
rgLRF4+4n7xFoi7K3JiYYEl4D560O7/Tl15BRp2jLKsweVFnX6STFWSG4rn7gPB8
lv2tzwvsXk4xBxlWSi8awrwJnHtOQC4us+CMf4e2sa0Xk1PX9bp4l+SOlx8iqZis
NteiwF9Et8Nf0e9s70JccuXTJJJvgjCIS1Z59IKmRQtXap81H0UPJF02nvCkGa6C
EANeeHYuZ4+JdT7F0xHt4zrVx7PTtUe5/OaGN9fdnKFyJy8eu5v2t+mJvUVLkvBf
ogY2q5nEoROtF+r/JfvTAP9Zlwx3N0yW7HhiiFxAmlMjW7rZSXOdBBq7GDdhCVYN
9fayXSjCCSzbQ4yngq936GYqU5dJSIT4lMHo/jnqSYq4IuZI2gbDIM4Y0EQ2i67V
ePUaLNqfizONKduCl4lb1TJ9zIicVWEEiz5/HbY3TtQGfBVt1nEa6wB/4jauhhLW
lGEVcbJor3I3b6/oXAABbACQfxq+640zUYZW3rEfHEAHeUx1QMowvJppV/7F0B4M
GLK1ICnZxan2cyNVU2Q3W9bHiJiJfAnFFV5I8cFi8XiJ3nomgaGXUgGLpgT2i4Ff
jtRp/Gbur0LNwrOR0Q2uWpJZVrCi/urwFOHzbS/VPoYTcWjqsOC6W6mYAIPw4C/N
eCiYlQYt9V+khqxgHnc3/f9Dz1wkyBYViBGb5iik3xkM8JCCLpvMpHKfOCbKuVXo
cyfKeLskyRHPNaWkh0qVSR871ajiAbt2RnGfCSA43RvFTck+Ez354484GnhB58pM
mPFX29cM/fitQD7dVzPFIymgyL5FAEjT4EAp5brmtiFrygeXf4U0SESXQrsj0sFj
aygK+5E6gKSur5BZ9MhsFN1/kTpTXBHym5U5En1BuBBUwhGHCPP4IZmYpGGKoo6+
mqvqjlnFHJRDdUISHxfYmW7UHPOI4UUjkqL3Y0t213yXlsb89MREceAmjvdlSuxV
53ITZMAZ0mxkxQtp2nT1F2Ro3df07oK6IhE+3ySDpomK9Nseso4Ht+06R2TzYtVu
KLucFD1wn8AC6Fe3ADn5DLtFG4XP1LW6dSqUzFoZdZQ075BrkuG39SN50/ttuG8y
+m1YOuTmFmymVj8yxt/1te/qjzG0ydsuM+S+kzllQNC5R9R4VLkgj0P51CSdh6dZ
okT170s6q/87MZf9NGIXtUDtILB98p46308sqOnktG2Y5Jd+PmZpuo9yfPrDiUhq
2OoAvHZ+Tftra7o1oH3MeGLwAx/eP9A6SfmMbXW6itpqcZADIREk4+U93JvpUl5D
hRTbt09++E6Jwhct4Cmcgt5mBK5/7h2js+XBd4FcT6COFtEQcOn9Ae04LDWjg5nZ
DfGIUPAZ1HV8dXTzvYYCYs8EY6eyYJwa1NLxkfkQu46VReEtNU6JzF9GVTSnkI3c
XI6UHuTCeecqMlIlLeZM02rdDYnL2KfvSv3nMGtaymFhfJJv297kQ34vQKVm+uM5
ToBX726LZsuFOJJIa1qgEzxeozgqFe2++eTGs0FVlIvAwNkEDV+ApyP4yhr9p1h4
6XEk1b6nkqPumHaOXNCfpsNiJBkcVHPv6MylokxAeYxzwICFjpg9NdzQhK9L3i2t
PmTcIxHpmnKjdV2SOPXtU3YuQb4Lyt3rFUNd+SKjxPGe8PLx5XjBNPB+qFly3KCH
JLBJ8avHIGa6VU5Etko/RyCcc2s00rCObfAaZe5R2R+391EKuePZKeVwcYArUibO
om+bWTRNr+AXhd1tmIwK174g9vzmwVyp5bcjtHCBpWqCV1K4g5Gi55rhUGeRY4Cu
UZpsITNmX/kNLqY3xJMl+e/DfO+oESxW/7snxaQ2h5TLZqahhj3ZaaPpPqtN8Ucd
aIerJHnvLhWTpLlZccDpTeCugT73WszEeJEvV1a/Qso2xGhdJ6RDGfgWggyF/IxO
sRT1XiOOGZ+ZSO/wvjVAsNAQTQDiqpV4VTLpBOqAzhUNvhZjdwMCgw4ZT7IeAQXr
CNKFwQXfUDQ2aGawiPG0PNXdAfRHl9i86WR7LRz7oUeESgba/AWWXW/Pg+eyCoNw
jnHZ1AE32TIDTH8I31bKiKfRYDMJjAi5kJzffgGb/UplQzCS6Ydj0FO4ZTMyM8p4
qYkU/jHR9x8zdqK/LnMKd7aZ3A/MqmC5NqVSb2DRVxmze1j6E0tGA7PpByhTa/Ho
G8sEQCpqqaBF5uG3sN+eH6oU5iY6PYhqYMAXHP3rB4TjG4iN5GtRYgIdCSnMvNxC
p2yDoGcrE/clGNMY1gX1/I3sRDJjaoJ58BfbvZAC1uGTL0qIvPozoWtdKAgXSIw8
Rz0oUfeMa+u+siaH4EOsuTF+JZahYUAqu38RzQkZ7dqumC5jFnQcwM0IVXu0MJzY
RHVwuXLcUh/RrqV+Qdv+ktWGKzxIw8L0ZPenmFeLwW6fBZmWspxVC1sxaR4OEg8p
XCAvqC2WplXsc4WRjTBGl16YkEAcae23Ct8lll1nYfbMpRPU65r1esnVxPhmXd9Z
nRLfS5UGE82ETNDoGcAtJX7WxgzaQ98n52NNNSVxS0xHqVvi3ieos9Uhpr7uBunO
XgEXoZHYJM1uArzWwkpLBGqDIIFY4OWPNZnboimjmeUXaegvkaIZU/wHaPVQJxHw
+Mt5+KmTKQqTv8y8Hv/adNiMDYukv/XaLY7W0IU8V+Vj7HJt+ohNWJNQzE5r2KiA
ppMkQZ8A0+NOl8psyBi47yxTTi+17lAlRwVDezrPOTGPBgFog1DTX69PB7MGw32k
6kTWlSg5AekGBTr6xaVfLZ15GJKoNnPs5BnToBMQx+Fdn7BFWpUmn2lNE7FjfuQu
F0tl7ktWZk49dJ2UdK2v/cW+fmL+eAWmB60xSqfL6P63pTLzzM2Fayd1N1a2Mng5
nDogZNhbtGtVIINwVVhhtHlPoMCHxbHaG0QB+eHV+lEhYRFMo7jQ9ULbhKPXzjjj
87jbYcpQmJ8BBXXg1pE5Xjx4sR6LIgPzRUZKNJyx6oHRLSd7khctt+74eSTbiFeY
2mV/H+USWNf/M9XiHa2EDUgKYO8H4nXh8slMv2v0nM16/+ba6ACQT7aomSBOrxrg
j1jPrTAgkwQ3eFv58Eaz7j5MC56Meu4VVvv3r4f5JzR0taXGyZ7ZVZ76LNRyACzy
bUuCFB9r93q3mbzh4d7gf0o0FxpckllKHklV0NDCwn5fYAvZzhNEJZk6WiyHkxJG
ttqa2SEfrXaAejfrNa8gqi9yJGW8S0n/RTZp4mgg+iB1wGD+GNGstGxJpk1Fu8gz
0iUbjcgRx6hzzTx/Vs7BJxvqk6prJ/9j6cWSWGbtz9aF8auo4jeuKnlYu8VK6K22
g5KlWWfJ0RmqTszv0B81dQZzbumvBQxhSigZUiGYyb+VWREzSF7N1dDiB+lAvFzI
N8r/uZ/XwNQZWp4DwcCqBQlowpGReJCd36FGYB4iDAY/ENrQSLAkdbGJ8RMf7RuD
O1WAvS4eizRVLs43M7WrbH7Cm9f8mmUEjuEiSFmHIULMfFLDy5dmtyw7Y9AcaCOs
bANqSHJS8Ufc4lmBkowCDUqVYNwy//rr5jiW7JQs+XDWxbrDAfqYcBl7YUDSS3JA
Ezgka33Hg0zT4g3e7vJOGO1fql40AjCmWuXlJuAA0VTzl4skZUi2OitIJApSLT7u
KejoVu8y0GO5hK7QvjTIpgtYXnjRy+b30QkCc8x2fzhYgZgvMJTa5Gh8YAp43Y0i
drF5I/V3xPReQZQYilKX6CKS0paVVvKCZcDc054oYkESVOtxES/Bc3F2AFu9+Gfe
1FHJkP2g3We9E61XLe3OPd7KkwECkvMuiFrt2GWbeIgW3wrW84r6X8BrvPKr0sG1
obaF3NJDh7G34vdSsip3JwE4sSWotbL53AXqurUeqA8eaPMLRU/6UEwPhGupT39G
Ky+5k8iq0izhTeKskGXO1u4bBoUKj09aocutr8oAbonc0ELLrO8rp65MzQ+U4xeA
d3hkC0f9WsgRhk4T4B5rmHXB2P4ua7cEV1JCsDTRzp+rY6ajCF87J0nCj4yWFPsi
TerkV3ZdzClUbujusPR8OM9Du7jtbDd2s8EejBcxo/LMOdC5bNT8R2SP1rb7moIh
D4QV9ZyvbZ5Skvn5aU2YJn6y8GrnTVHJIDBnk0gzjxekEiIlhkU+iwjVNpEsnD8H
PBat0dJnWZFFlgTcce9hUyPk0KCucY3klUi2yYsIRi3I5of0Ec+saAY7EpSa4Inp
JqFFbJzvV8e0hzr9i3q//eXF5ZhFg7+Ni5/uAsllaCg3kLkvwsqLNVhrvf4DH7LL
1CIyRmY/15KMDBJgCy67CgCglmDxJWi6kOt0HK8dcNv51t8yup+jYwcg7lI73PxO
1BwfXl1GJMnYCiwApfDN0pqUF3uyXQuatPvmSNRkLl02s0mUGLeqwTJ7PSWqMEI4
0HU67o+FEPBpqsPMPvE6LDF5d6SjNzi0k8kYANMB0FhV49gAQNjz8tU2LYtRfVFp
giZzE24bEu+36ZVLMQn2mn8HYB6cq/yg4V4FHtyKAK9kiMuOZDI11pQI2Zp72wRq
Hy+9oPK0SJrnG3apQhukL6DdmmpFKPQu+iaMoWEzlOHFUucSOHY5eQm3WcPTzZvG
XO1OkrAd0W6UawJ0vcB3tMktOFaasdcTsXHTUnhM4jyZaXupoITg6R2kWfNGH1Wp
1kMokU2ffS1VmFeaPlTIX/yWMWD5+dN+RTO/Fk6VO9g7sF4AOd9xMWh0oV5bwL76
U7uf1nkniAw4HPGOZPjWxozMeiTxblJM5Bj1DeKdNgiH0E6EHrIHMyr16HhEoGXS
hs+XgFv+jn8XXab7sq7jORC8ECqwABpTFymfniv8abwElba8ajWYJNNsfypbLKsf
FP35D1tdDRAbJazDSVNKTX6pdlHmUQAtsvTxtmI/HXh7mMuFUNyxof0nBtGfznWr
fcTOQi0pZ5NlmG5d6TMpI6gMdzSqb9FeHYW5VCgbKrHtSvGkrM0uzC4cahJbK6pi
pWzuPwTUNCIHEkjtUmrvmSqc38pSpIvJB91Ned8DU4Bwm006s8MAtI5ci35J+rky
2qFU8TLKfiQ1D7KIKmOdbiaVL8F7Hooz0WhOeIbQ9sByTQKpWqlB2DRGSVQOekTj
8nC96oN/bhrn2MG2f7h6zVIENLb+6mZ2w0/dpup+acHhq4YtxzrAIYYjCTNHbi+5
wRNQ89hyTGLjygGttncZKKZW/hHUXYYNbvjc+WJ8+74x0l0BJ7TEvB3XKbglewSX
gFmabrHClsIuczWYKhE8pp2xJT+1dAWp3lmrdz2L0qUPDKwajCyJOvucE/3EdN+b
iKHM8K7InwJFcIfvgZy81KkBzg+cbO+rG9Wywi16enLfGwXipwzooqhB8HU0EghF
q7ec+tQiFzYbyfNzc0FKONXeCjlRlZAYagKngrNndzld8yCRUC7nU4v5LUuiXQH5
N3M2gudkMOdVAamlQrHf7wMMMC9oKkVvodo09hwPHjKH5DAEygAkAZngcR+QXLyJ
GE5W/ezlwNKHT7CM7qZxyvzX5nTa2weJ27rXrtVqqXwcQddXC4b2L8rodg5HkgqX
3st+vcTojyHTwHUF0gqApFtGfl/xYPENlo14FDT2JPRRYw3q6YCWtdF27ttFNMao
j5dK9TYIJ28oOUpE68PpUe8yBZonUtqeG2XBk2IrXMkZf/s2AKgNzRKBRyvSC8xE
fISX+9XvEDWZR0Khf600mZfE73WvsyFijgENUU6qB5y2yyN/71J22pkYkku3r/EX
Co7XLBmuxDgt5RH+q+pV/9kArObPTXi4lM7sEY4cB1hhiOO0l1trz5iVD2ocWnZz
98qCOX5mitWhBgUOHafXUjKQQ7W5umGOHISrtqR3bilyMqPXf4sk+N1Hp4MOqwwk
+HiCm7eWGT0zfD774e+39km9tMwCKDFsr/vqfnfHOUdvgOl08beii+83hlnqKZ/K
KXITsII43y1MRAZXp3yD+bjn/tVe7pUQbXyzDSkoTCs+5m96GjTke61MRZu1l/al
U6jdtumf/85O+z+FscpepuhciX1V5zAQPE1YWNdA/m29n2+VsdQy3sEHE7ZLgnUM
Zn6xe/MPU8xbBAaRE2tTKgZEN7N/HfM/rbStRqUXU1RLbALUbQtTe0LOTObJV3Vg
9IfLRL0v0u0iQ+HrLbZbzhvGWKkl1UwooLFhGoo4BQzFvkHOXn04ak3GS7abHGYp
7/C9+Axt7exuy5ct1dQOqu3RfpQXbteuhukUZ//kt85BqfvjDkD87VXWadMKAvtc
sooU3FuaV3Znjx1IHKvYk7baKQgnaVKkUK7EFYIUzHGmCbTxw8nuNxL5oCu3uaSk
7rwIkU/sOWH/NiGf8jiqNyVWsuC8RC3SX9Jmtlp1zweYKm6G4z3fBjzi6omfk+jS
o0WlFCQXotL8mg3GZ5DbNhtPFoUMX7az3ja4Pj1Hy05aVJ7hi0sZXv5lTz0Vf5km
Gp1UNLYvQXaLvyVIwCN5XxiZVbR9cFe2hrFnksXubvf4rgh4u+Hh5Rgh1FHST/Cc
7LlBSWx1HVLOR/khwqwyLwF4tUoi7zeA3kBoi0qIdV8pnFa7WFbi1SxZ0mGH2vEv
75YsR2c90auVFTKqSAweyCDvk50IlFh7xnrBIIh4GpGKdhh9MbGQaIIdvlvVEhgN
+ES0FjgaLG57rVkZXnhVgad3tYrsPIMk8xxonGREAEKKvr4cHyhNQvqhPir0s+C9
K0axJs6KTisGpQfEG+Bz4eIkkOH/cFjARv/IgBqnWN5zim6stET4SL2vz+c3XOzH
sZlxG8iwhxs/oC83vmyKni8QxLYZXkYeDgND0zzvMOqadUPEZQL1sF1OxDXasqgN
+O4zurpsDnWrZ5T8djmJKAVM9+mbAsE+rmBcUsCCG+mbLRcYBqEAaZb26xHxcuNm
hxc+6bhxY5xY5LWIptIf7m8+gBOkpWohTsVfyTgfXaMZ/wFTuJu2/XMFg5qjwiOk
Ftzs0b5UOZYwGik8kIUxpvVvRza206xF2nZtKOydL0sB5PVZJ24bpPBRDwqgvmYH
tM83PgpUurwHSNiMTOnGxpPY0+4hFGGm1aXsNQ++iVvcJPTQBHQ2dVM67/11vYwA
8Q0dHvVRfP1yld95RrEyyqO6ZMW5JCMtDIwhw/LXDdb4FtvS+sd9taZIzpTwH3zy
cTrLJEf+VbwABJNY61M4OWLrQSkWU4DVBGMOd3Lk17fxQiGxfQS4QhoWw+p+3ZMl
eSQSg4h71AKIG7+BnMrLZfVtoj6EtVb8C/ubdSbP/buFQQKlXp1aDVKFBJLdbxia
zAhN7IfNC/8VkAas8tS1g0a4hBIdgzyyJZth27eu9mWmLTxnanmGCdN6pfr65ypR
NRDsl2LEV03T/7Fs9bKWBcvc7NJItkTlAhxaUkEvCUXFIjQRmyklGrYkCkMNbj2I
WaNjSKRmJ9PDjT5iXG4uPF1IFkHCX0k2znxW8Ub37V3z+MJ+HxW9HReehVo9odOL
zreYkzUGnUoZJztVdpTLsn2VqiMlLyB6eT0vWi8vxZQgWGtz6D5MUGXUj01C3X1P
/LizYmpEpnPSPDLdfj12gBT0qUsGSCVICN50RONTPXAzKH4zbmaTbEbWGurRddhY
PFOlqJYJ5lo+M+DgTnb7EfDp8H0JmjwH17IjTklIl6WgEA0OTqITyHjHZD8te256
bvsitnePQ37OvcEckwKkb3Er2ULvkBp2e6VsmCT3yNaPAn7XV3sVw1Ff6y2Cujh1
EFwpJvbg3BL8A3DrcYuksVDfmR1sqfNxeOMhoX+F6im9ebVd4OMOuivrxin3IR+H
V+DW8ftsLZSUby75JDO30XHTw8AOhqgU1wFDAXiAFisEEr36Ff91RoamRye9tLyN
XsGnm3OOABJbxOWZ9vPi9kSM2UFsCzthvsswJEUgpd74OiHojxXZ9r8W5laUQV1I
zVJ7cwC1u6CFQF13EUJDc2AdsDTw+fONyR0Nm9H1QuGU2UXN6OgU31W2yNN+MXqv
HW1U22DaZYBs6eV8B8CF5j+H5wHQ9fspfpgC+WNynUR3/0q221MGhzg3HQdAxp6F
U/9I2zS3wLG87wih+kXdwMwQ6zTT+G8gCjNfITXCWkDop7jCoHNMlMkZyiC2XuR3
biltpPUgmKdQGy0cLVpu6hVCGdOaBt+N0J+NkHvJn2YVdEJmpSOfm+5Dy3q+vfJZ
0OUCxYKR9CKfam+nuZA41xJJWxlC3172dqRLXhWcQefjArz1DqRrURe9vagmNXMc
LFtpzBkhFG+rt4md66u+iffzrb9jx7dDF2sIXlW80zvATV5ytF4POt4TamZhwbSa
VDlvXtgiK+LAUi6fz389wkIIlYfS/rnD35S1RbppE4HWSF6M7mP0ckoz3itFz/ol
2SlFxWfqrTcOd4b0OANwzu1+iFwG0rdRXvwknjpOGRj77yfNHxWojecuscRh/ctp
b0BSECXMRKvh7BDS0GLFBJTcXr5D0u2grVWBuiiClQG/Xd6hQHklZA90u5bZaN33
EHMz1esSa44K7MZ/NRnmiQdo6+eFTfxNxT8/Scq0eSwqINn+EzMEIVOzm3DNInj4
I1VmTrwXYE2/2818xDMhNZetgJYDjBgNvc48RNcufz346PkEnCXDmbo4UMuE5LUB
AcL55WqqdXGnCilfSwequ/cZgfPamXid43M8XmtqmflBLShLWPNAJFtJk10CiObO
7eaamaJEKi4KArck2VFYENlqq2eJUxhZOwiSpyUuYDkSRLwtCRI0czbF7QxeZaKb
SCrmUQepbwIohcZ5wh9jN4OWx8SbnhUIzxY8LTUe+Q16QkMZWa/3NXkMzrhSnpsq
5Pt7xaTx88o9PLZsHKDnXUbNpi4s6osXgmt1fGRhTCBKKXhHAxli6/lcuXZ9vqgI
u3Qv467qVvDj1N79GRMTK6qk+Ov5vVrQYkdWQa34llNWXGzqFe4m2GWqe7mQoBn1
2T1E9iSbC80dEHJf4qf/KUtFpN6tHdrwAY1LVm6VyirZhkk13JCgo16bobjY0baw
bWjitJdogFwhkjCEwYFTDneP74+ztcvNq29HgN25FCDHub4WfUCIY2XeYCR24INT
fBg3HXi1Z2QtvaT5XojdT3hwhl9Z/Q8w/+pG5tnK/lWtB2zW0gkwnvBlnfM+Wvwr
VDTgyjCKPCeZTXCCHceMP42mBO8zB8ydZByAkCdd+1qhBYtq6uCPUKDwhB3teszl
1AqGnwNWhJYKIzRwyLtYi4oremqvip2dMIDOMZ04WaudtTv2NvVv1DNS0S75qu5z
7+5v5EKrvWrX6u+vOHBzMjziRN4Oj/X4nldeYQ33WZyL7CHq0cCz77uUYDuz404U
M8OeBUsYi6cbqbCuaaapQZCs2m3jJvN0U2X5W5Mf/ftJmwW6AJeheHwwPyWxtDVD
eeKwYkC428ME+MXWynC8O6CqTRVwMUHR7z2JPpTrIEg29rwC+i6stVMWT29RcUqa
/yAuQG4s9PRifGRAbmXJNMMBBqJlTAYSYbkK5PgmTJ4XyUtmTte2q19Bh8SmYjvD
eCsW8W+A2CCJKazgMjFM/vPkQ3DZqYUBcb/kTCaltoCkNtrzhrbCDI3NGkXKl86q
IjwaLNYLwS7wQCkFKabCjBU29YhuAAs/zP7q16nPBVP9eKlM3/aGun+ygidGhYnY
H3R5P7XfvSW+S36maD5NI2Khtdjkywswwpnfo/KtMSeHT48Q7lZejijc8a5Pv/L2
+Opr7zVNca8mvnkYTt1LF+TT6/2XL+5dl85VSQN1Ga+C7YS9gIO53Mau4hr80eHu
uAPvLjqmBKNGpPWQi2RCixItFS6r1UJ9hL+i1T9YDRx+tcaH5I9kobMlTdsUM3OY
86fMJN/eGeYkKo+C01sxsHQTdLcqD1FsrNXEFhZdWnLRMTOCUFnbx/M3AdpVoXaY
exgDHggoBEKM0W/n6TCIZawGDYY024hfHHkr1sHwAwVKFIHJRkDNSyuZ7MR5JmFV
N0KmxqkwfMEZyz+fjsZZQfY5Sha2qINfGe3vjECjOQx6m3rg3MYfPgd3frmvuBZ9
HxD+sIVTBlok3KmkaCE6szbA/MWVaVkc6Osc5iSmsSzVitPSxjPSA42f3E9UlO5E
qTK92VgvNY19p5Ek62kq0sV9u8BHNZdnloIbZVaORMWdgAuIcOZN4yvWE3+H2FSy
0McJ486Z3IW95BefYhzfIwB+YyqOm9+702B1j0M1RjtMZ/Dp+10PIafHiiRynnLa
3UvsbtwS579FB2l4syyB6UBfr6hLvsdqxbd+I0kD5iNgdMxB4Uh9m8JWvZjFEIGG
v2O78e+feFBUlI7Mh80zDq9eHsnwhMAFSFpDwEsI4DifGIX4s74hOyyiDcd8/GEg
zySArllvoR0MnKrRJFixayLw7rIvWmoFF03FkkxSHmmaZotu8AyCPNpckIrL4WOk
TnFERUkPJ+VshLRH/+V9/8UwuHo+BCPuN/ake3gGwMu7eXKBFNgEHpWYxd4wldhf
0Gcw0WSCJ5162IBn6yVKvdiwIr/Y6oCiuWu7LM8ScSVARQONUEeokDfKR7IrgBag
5q42rUPVY19BpECPaBLTKkeCasXtNY6RBX28tDor+1+TvquTCF6LYiU4rdpk+M+i
s1ol2Kvjw0aMymA6q0VL/cPibfWInuzOSyfTmH0sRKDfx1dSRMwmW0A+L/zi+fxi
G8j01TCeIOG0eQXa1KIFVpkK/XiO6P3Lw3+7zrfB0/XFL3DjtX26RKmWGtlwWOnr
tR0DgJR4tjKlEnuMnJBo74Tag1GJuHopxHWT7ItI8W5Gs/FPoTC9maj9cEPYVB2t
PFzdq0hrxYBlvjSvMV3irG8uHjqeCWgHlfTile1IwxWDGYihr2CEWkjDJWr1Fet5
pHMdBqZVhDsjBomZj/mSnA3JbXkcXbHd/O16jkDzWCozdAZKmMq6lBdL1ScJR7QF
TNgwxUH8I1FfOXrnVC6CpI8AiVEVh4bP+/9TAPT8Egep67fTiIykDlrGDfzww1Fb
i/S/yB0F1Vk9AxDphWa1FedNsd7sUw79vwZJ0kU+dXSsCMfbBa0/QGgc4I7yRHuH
2CdA2184g6um0/4GQ2ntCi8ZLdz8fnH12bUI64I0Ftr9CR2d0aUwRoZAtLgN0sti
Xek8kkUj14GUXlkwWAlUShJJPvJv3O2yQZGmwq2DeFtOltdVA5l4MTlWC6gdJNim
46ViepeYrAHHuR4A2+fXIgTrebTECv0tw5Aow7IyX7D2Mou8Qo+iRdfAOL8dOMlV
iTJ2I4l2mWhZLWy0HSIThop1GmWcMaGIrkrhh9/Qv1+uKKq3aK2xLJDN3x7Fq8bl
BnoVIjsrD1ikL3+UYWFI+SfjxUNRScS2NrqTrwx72/JSljJZsyqoOFBohDhelh5G
PBn5zfaY8fIbubmoXUOH/h6gqLvj9hggelYyMZjtWT9gna1/xbDinp7ox0w1rySc
JDvdJQbIQ+JK13x0RnpZgfNdpELHApZFQ955Z7I40D2CUJ+UXJfIuynOm7m14gFz
KciLQD569aGfUQwWKnKbiMU7jsdyCXhovlzyNZQqLAWYDSgK59lVUtFY2PXjK+tq
2MjQktcVIo+DwXSgQY5JbiCOwqyMHb3kNyyAVWKxGJHvWnjU/CNZUBNerl3q5Y2f
ypsfOYkwp6U9IT092uUu4DdTWeT2ebD8Rc3Znz7ubpemhJEEAyiGgHKdaspWv9X5
/YCgpaUwdmIVgRx22xcmIandalmDf6peI8ooaJ5vqw/yBGKvTNztJ1Xj1v07d7Zt
EiXNm/cGmTuHt/9RkbNzAYN6NHdy/CRtB3AOgeRtlBiofygGU1f+U+YuEw9Rhf5S
5Nuklul4ibsvHfYyHKQZ+Y4hFOpsRi8fY3wLglIrKLLaPbprIKcM+BkHJitFaQYQ
D3yawF6Mam5N7WYBKHawWdb5VOig3VC6zrhDBArXJ76B/WplaXBgb7EvH41MOQaU
kLjpcwobCV0p5h44nGF7R0OXapVeEtnsnpGGQYvMn5DLKdyHpia4h89jP5i062Mq
odqxth9+WvDNkakgZ1A8KNnCU6+ayHzbeOjRGHnx+Z0cyXFyP6EpqA5nOCRQdyxb
RsX9CcUL8RPo5HngD84Y2hQatjJn5/upLSuQGxGJswSWJFauUW2uMZ5vRWtEIzvq
ebZrfBFMoMYqtyKH5bmD5kAddiuIFKfKmkQFcHEXFO6/rQzePdVvbBbIup0kBzqr
h/rRuoquaBzTIzWvVF+aftY+4GLsuwBhmJ0WIZI24lszlHjubFYnuO8U+3ECcku1
MTwI/XcAJriUDWSl6r2htQ3dmO8u3BnGGtN71AsW5qMdgRyU+n11b9eIj9gMeDvL
pvUqWaWQciVgCj1voTPFwZ7X3KCFRImPm1nDAg6ef7iuoV+Q8og3G2/ia76mwjgy
bVW5YB17uI/gQcsB4sLcS0Umo78vvy/oHgx5kKQxN7jRd9rQXkBS3Qm1J4egt7+j
5Jfa+JuPGPjO1Wi5Jb/fXVWt36nWpI2+TeicXyVdBxU96DwTUmdG6mMnDVYbh/Bp
tYagmY9e4bevcXLXW5KgIyLIDRR6ikqQkepwCGRzBVUGw6HP3bWYVB8oNeLEAP8c
uOltZluGRQCmdpX1U3EEIiiiH9CeL8l9+azaAw4zpKX51rVG90lrXhr2g2n0pD59
EiKgqMCXbXSEVNAK5ouCSDBlKieDmKpdmiSCidlv7rPoghi/cQVZYShdkwy3Spox
urrV07JiiI7uDBOBZtzFEqy2EUzfYVIB5wnADCFVsD+7HO3NKXKyKjBTxcjN/xNI
qhdwlG8Xv4mac871khriXSXpQL6GE6R+dUm68LF2x438yY7KvFsspzASYHLzlQwy
hw7FS33nunF1xFz3HX6y76n+DPBG9ky/rAk4tgs71zGbQ2LvEHkoaYIkDmGE3VIx
iGPrhCaczbQ9Mh242P/9N3ZpVu0NEGq83caY2HLc6tXtFvnKoRaD1LFcJkRlbRvp
gyh4KJ73OJdOv3T7flLc57mDrO8HnFexQXN/Iw6jbSqn+me3//38dAE8VQ5VP0+k
X0eFwrm675ZsXcxaswLA76K8Rh7HpuKXpnDZP6RrMUSwxeW3XYEhcHhkBGZMZSqm
FNV04RSw+4jigL+8+gLXf0kk1wol+HjhY8m/gsqXCSPgJSKeJgUNlnq4ZgvMyxTJ
TbcxZ1rsCdcLJIMt7kGwu7vXnX6bU5QRGnRhauhnVRsfEWgpFCpWdC23eqSoEUVW
dZbTdB2Zc0XAnFdUhNflKhWz4GNyCuYiJ48bPmCdXPpxUF46a8oYEpRBPCqb6Bn/
iB9MQ88Bgn4J4+a+WK+LkfAYUypbsCcFIJstHnEJokixJ51JGQi80SY5PwMMh/8s
fDQVXc/ibF+vBXv1jIrYp9dwDOlgy37PvNyTW4z0klCKknarVGgBJbO1ft+t16F1
YISoHeloxTOpPjVc4Qd5xTxBxO+ybjyQKpNG+bg1sTfDZRwfZacg5gg7OMQyXe5R
DVki/wqc536tLz9c7MYrwbCak64/6GpT/wxbcVL4TyEg7AdbFXVzeWVQASWMSj1s
tEjbkQgdP+lhheRqFeYfSTMC2nPlCpBLEPZ/ZuYoYwegBO7tlPH3cbL7wN1VeAEb
VRO5slK5DZZsjyCnjTQ9kZRhAZh+Zuz9YDVprCXWDUvWj2F0Ww0HiGqeaE75CKeQ
ULPXA0eKEVM7+62gAG3a8hJQeeFnvmo5JytkngFoH+vP9EBXxIAmPqht3x3EAyAL
a63IaTy+J31g5yGzLRYJIaQlPrkqCjNzNbert2arK2ewnZJ+56yuHWPWRpGLn0YO
3+bNTLOyNaxP6bW7N5hRjjcomy1qQP4Vde/QCMnRQ0Gs99t8pssRbb9q+22M7rat
XafMFEafW0ObAdHJL+5gQRKda1mP3tKZW57BlXUTyCjgN3YCU2RNYzER1kq1LQd5
1+c9jpESKyWU8Fy8zY/0ilDPZJ2yHIXX3+PpmuUbtW487Lm+z354b1h7KCt4BdBZ
F/d0+O1K96X8h/hsS1rxTKlNhzbT988s42I1qIWL+dqyHJmqvYUT9ERw7RfUtUc/
tdTAwvO/9K/ME/4bB9QM8wRf4+Y2lImAmHGOEPto/Z9/Y1YRS/RxGwidaOcOnkJe
gr+yv0VeDAdBuj653MN21MDNIXCnQiAhcbpbICoMqx+czkzE3m90c6zr+zdmCuC7
BQri69WExltRoqUCv904d1t7EUyyzhoyVofLGvUtHycGHlYKSQWOPWEcRdAoTNhW
JWgNYh55jcDyeK/+8Lqxc6xXi6uhJxC+pY6G1ZYnJqQFr1x2wtGh0V1Ey7o42B1b
iKR7/5oWU6gNy2q2gSwiK7KqudMGlLKUCSvJG/uWeQ0rk56G/afKJH9r7NSefL09
PlbDzTKbq7JGTkWMhaSC4KXNM6R5dzDtZGq7439L/Enj85hp+oNMIRrJhy0eyX7x
ntad1dXQ51tC2qQ4TGAneUZOu98jmgp+fPODBi9AoSOogqmo+qL56LeNi8x6vIbu
ZN51EhD7xAWzVMVdxCwUWh4BNVQ+nwE/2n6g7jQSJWhQVByCbIKKfB2ZlbDOIp4t
cIuPfE1ZFA8YVRZd4P6KchDN1BLkHo3coLPSrVw1+D2Kh3MjGwDI3eeJKIfB+BJj
Rt9M+k0VwmhBcqA/Z8bzWI+8TQ8haTxJP7LNA2adJKnB+l9Y/RAgQe0FEDjLC2Fv
yzl0QJHj5dU4GnLsg3egMYx8n9DXDFq7nAHpdptvczURzOp7mJnT7dmvJMRgvAaN
p//UMI9v5tILAVKdKDROScTvakH9XFQdT312Gq3YfxAhkHGJEjVcngvJLANhqfha
ZRDzlUPXMDa+0lo2HT3mar0unrxPbYlgEBq2eIfnPScMd2GXZ6BE20Wb/r3X1i7M
pt+iPcl11PftaCRcfjgK58Vw1qmElM/Z586+tI27iO8rDX1ZHTDj8skM1hpnc6xt
i2siXSlAFYNFCYhXcQlvjg7ovMO2OA5yHbrd6sdaCSnQ9QwyZAhJnxUtTuJjq+ru
ri1E4A0T5usZW/2ofo4Hq6qqVi3aiLUzIW+/DKsF6ufIhpre4roHzHqJkTDvynW8
gMZmxwIjGsb+ak92OKsENiII0HE5yBCg0UEdyceXGg1cQVTgCvaOLZGJDsKKTWpR
SBdsSF6jFQQz6Ut1i/oIRHUgkbI0iOiNzyTwhmTKYt/tqPqu+L/gzxjI9GSACN44
DXUfeKcnAmm0BDVhmPLdPZidCzATVErwkubCSm/x8uvOQmTWTINI6bjPKr5WFt5/
bXd9KAX74XOkoZA8kPUAzMPGQcjyzYgikC/z7q/v6ayDl/HSv2p0Lgdm3Yz0eWax
CJ7xOXTNSgyEq2+iAbBn6rRf+FQPBI2ubdSgsQMEKmdQwLCjL2hu2I/+m7ia0Wkm
mF6hByexw47+7vx9pEYOtlSLJZAqeOSbO2LqrF4wToo6TzabQlrf+NCOhmLSaF7J
3KXejhKaJU08N17wK9pdCQ9eOFHuXen/eWIDg+yujTpAz74qyCqq2Z53LV9GywSh
RP+IFRQZC1RGr9C3TQHItDI03TdOwCXofxBW8xlqNGEv5gwZrZGB8ZZ874x54fRS
sTWHmOm5gWwZlX64kT4LHREapxD6yUCMHV8/11S/b7ZMQu5ku3BiGXg8VNdwk8WI
FAGJXgsi//RsU4NN0vY4KyVrCJJHXmCPvNqv+HZCTATtUqHnN0tKhd0LW9pehndm
q4ESoF1ESyajEmtdz8M9mo1NLuJ2uDTDl649JOl9Faig9aaWAP+wBdj6MjHAhzMY
5jUiB0FR4tY91Yqdp3YsYcDUNEMUfLg3NvfWGHhCOAEIZv8y4ZIXi3Dt5YqcdPBG
F/5jK5UKZBxeVoc1VKjcLvsXb8YyXr9HWhMxtzBqNI5MGNjLc13gsoHztY45TCZ+
+0Vyt5klv2Oi/01ibrkcUjd/mXwGCghIZkj1RBat5YMtAbtbDcGCXezLe86O83j8
NfB4hB77mjJ4oiFmBT7Lw4VsTQgY9egUPvcOqs6/a3tR4olFsy0tZ/kU9d80A/fd
//wBBzDBGApXEZncFN0MoZSn+p3e+1Q/NUMmGwpQ2cqRWwPpQk7bXYSDit0cms3b
bD9EoRDuZP6v/1M/di10NszLiFoBdMNeDrH5CB159ZRZizGk4QMbprXFABXTxki1
7DzoYfYPz0RCnIXjMJrGXi5FDZwkqnoFs8FCSbRERadnqTboWcQqwX3OwS2a2lRF
GdKiKH9rqpbcuGTqtb2KzWQPO5PzZ30AIhrYSBHCTb9mumeAzIcmBb3xe7jTdqNN
+de+g88A3UPUzcXnaCyAp3xYbPIeD+IYGUXAX9EMOqMfqyXBgw1FJkJGBimFMLLd
lRjKF5V/CdRp/vXNMxZeyxo0WgtoOvvTTzL46sF631lU/u0Ld3ujBK6qYq5JDTeZ
jwttFLaLiaHNL0Newmcr0lijx1Bg6JpTCzRmgL9VpqYzVh73hjBfjjTK6BfwZu3+
fieEEkvMagGt4fWZNxllnE0jUfFSfYG6S1b+6YEJiuhKkcT2ZL8M8Ez9A1ajegrZ
DzZQzq06D8SBHiZTvcJL6MUWjwHz0iZ7L8zGau6MYHsEFwrCz42n+nXiivSwpc4R
xw2nZYVs9j/mMv6slgEU6YO8R/r+cCKyEQ6KRmqws9v3FRk5B+fMfPkk9XmPzi4p
TlgQKjQFqZYWnrQ+/Uv/ijkOJHXFilAmyrESqKn05aLrwRETe4A07foL4zVXEsxY
0dnmmljaj/zqpZVwsZGa0ijMxMqDqGClsfy9thrB+nNGVX3rXG9Ybwh9/vnsR50C
q+BufZqqoQxHZ7hmsHmyFi4mi4PGHQXU2+1q1ex/Ys1Tf7B0VahL3joSnIt6x0pb
4mPhF4iz0pNlWZPfsyQ3g3NLFvqcmhL0B1rPQEHTDken8wuN956zYW4ANhn0qZIH
Oc/1u0AuDux1m6CExv4Lso3kt2V7s85gXVJEpCe4ear9h+e4T+QHV2dHGXwEkWQP
BBPhHBdCV3e8MdCr1kBMCm2dnLf0GSeg1sudT3Y/Qc91pkilcvUF/JpJta46+OLM
klo6Dzu7C3PhUvvM2Dd/DzpjiH/ZhXNP502tYVa+TCCpaivOVqbImSbk87Gzn/jJ
lK+Hb3jdoanaTajOCd0WPvg1sJYMkTdTSPRjJBTnCBbepwA4VWeiVb4jz4YFo0XI
62tDH996YU3MRwZjlWSvoeG13zTjt83jw+rTUfuCjBkoQs1JABe3tJqzPVePpLBJ
64S7AyiB7jQ9h48sSMlWXB8dXCDFiAv35MH0yizNfba+Hbo0bGC5lJny5YF7eHie
giI0/JTP0rN9hzpg/AyemUVp0rd77QuruO07m3ShdFR/A1LELgbbv+GhXbRlOPc0
1JvUBWMbhNyJ8+9Mvzhkr655pqvOAFthEZhALmJtez1SWxZ4rA1QW3307Ex7DiBi
32PNVFExncs6li55puoExwmZNsuAH+ReQGGTM8Qfx2iO5qD7xH5U2ZAFHnTzKlBk
a25t/tgWhNur9wLQyp5k/oFvjuNhAwb2xwjzW/77OpLxU+3WF/BFiDdshAmwLogt
0m2HRXHF04tTa+3tnwoiD4N/bY6o4k8j7/QeJaIpG3AIQxjaA+pX3vWjQu2Ghm2y
tQohVpKQeUXgxbYV0BHRvndMkAqwvnJyYcENpd4IzFnwkMRxr6Pl3UGdO2aR3hp0
HLVQtLTQNKT1UV5Bd4R/hCbOVq3+h5YdJu75wk4vaNtmnD9Ls+TZ+uz6CMCGvDx0
4i0UwH4jmmSleZDOmG+8Tx5WIxyjtaieYCEixzZNIJpIU3n/fvG8EspRn+W/VL6R
g0exLS4LDOnOwfjn92xVSUmjPCqN0pvp+7lSfsRJH1lzDMdWSjU9ovvF+DHIcbIB
jEOhSfbsreWQwFP11r5bOIUdKhc4dNDZzrW/PfA8VfeSZ30CqHPvA/lEpL/eJ8x1
tdM+Mg7KGbHI+TTo/1jyR1soyLnVCjyBfXeTccqyUyNI3DCTXdh9STVpmfNwgDTK
DKqUItTeYOa/0rFsuLHvEqeLsQkUcUXp3Gt2h1uBmeakGodWARxojcuKrD3VhI9C
fhz1TstGNnNCjxwA2lkacKnqMML4CBXJXSMJKbh/KciLLla69Uy21uVm5ldBrUzG
11R3wEKLzIEBFTqQN+tDlR3Lde8Rzs1nuWScg1mRTcFWUqU/PQucxoHUhszaBauQ
2BUAYRF1VxE/e+JHDQiHCMe8qdGYrF30Z/SaxjXU5pdwfpmeYrPWAHgWnMRd9i7D
oV/ZjS2M7G/qOjEr0wgOhNaChPsn5m4puln4ZpZNZkH6hQiplm00UBQ/3pBOXO1g
Mxmd9tUX5Q/QDYKPVnQi7WWYhePfW2Lqo9k7UAVy/LXj0B9BGeZQ+VNGAkRV+fSk
bI5mOTkJaRGo+ilNK0xiF4aFZzEP3Z+r9m5MbKYmHGBLvmX6FArLp/Jkn6zpO3Kp
2vqxwfXuyPiYYl5tIbZ4RANWmBlynkmzmDAK6TK2O7KkfUHAjnWew+yGvOtrU2/m
WiBMfqwSWJthBZDseR5NbA26KxvDwjYYVYd9+glHd4zrI8lNzrHkfL9bakh1g8IW
Z3WOJIn0OtLQ/21Sj9l4XAdx+WqBN/FrReISbLXNBeSOSvd2YcX7VhkFp2Slb5T+
UGM9xkJCBYXUhf67BqiUI92W83PTX5FlBWQNQWj8AOtDxtaHKIDJkbTvvcUk+tV6
QvzbkdnyyWNnhAxM68eBoCwb+t7FIvOwhMsh0WqwUm/mDuJxWh6WOWOTpU7UKSOb
p3qYw0eJxlypN9z74FTZCXraGWSA9fBwWLbDRZEQ+QQNt9/H3rcdYXPsURc0WhcL
i/bx6/PvnptJs8H9ICBTnT6I14il35YmBJCP++19nByq++I2rvewQJd+atDNii4h
XfN3bXMLaLatwgyAftUceATVPqtEFp+H0FZSDHiCj+EfDEi5+inogl/hHDGzF632
mnQWBaIYJOKkMFc27cLMpAjCUuel++FugB2y0AJ9oJSmAbSx7AaEHxiYn8nImJOF
TlEqlDIx4lmk36x6mxE672t2UZeKYhuOS5pwraKMK9yq6eNA1kWyyjJ+V4fFYYl6
XhM5PYt72Io3xDZot0ALsrgBuz2wlPjrJv5FAms0bqoU2JzEKkJT+qSZBCMBXVJH
VjOH/kVmRayUSnqOYW0nEZzzBhFKM+68s3MaMRQ+h9tHyf+Q0elDJUoUH8GHyYxJ
NxVg+PioVHHQiiBjUnDCcJdcSOZQygbJ7LOEr3jJeUA48DZMbLa1SwutF7MuUicO
5SghNoDVkw06J/OhaEAAAmP9kgLxrE4u/BbbfAS4S1lLH7MfFQxRaiz/2nD344Uc
/VrpXzIWAu8Q7u79iPHkO+vbHEyBcvji5NMOrI+63FL/VSOeBBSK2CHLFSdcCfEw
HTOO3BlgcyQf/VCLrwuuxyfKeSdngS2aKJXcnpbfTjxSgMjQy64Zn4+LAiBBWdRp
c5gmqgO0tLE+Hjae1lz1BiT0ZWq9NIRwjZZ4opKTQNxKpif1dKBGZZXNhESVJbSn
SUqaH/+8WO3QzerhxHu6CQ2J03BhLZ8yrra0dRJx5aQWcHjaPi83N7+EKl5zqX9H
q+zDypRR/IB2mZbdnIjy8Z3mR1rAWa6GIfX4nfVMDzq0r2sUZpN2sMcjz4D9oqW9
MTGE7SVY0wxCmSo1yqYX5Y3Yo+wVpRbbepUMarzpXujlYbiWUN7vVjStQ3Mj/uOf
le/G796s89faeY2uFv6KNfC226C7WxiefT+J7I/EmBLJmrRjfbUFYeU6uka3jscg
C88hk7j3eYzhu117ICK2/Jk8cZLUDLpw8TXtu2ORS8uu/yQ0Aq0ptMtouSLC6RS3
J+BnPFd6rtHQ5Z5CU7gv/JPW0iaDSOSeZZDZvNXCq+jHMDikojCyHjGvYv+O8Chx
pRLI3o0E5Q4/xiD/2srP7Kz7+2/ybpDOiI5Z5ZmafHe9TIya4dkB09gB5VSkRtk1
mP+rF2pTytqvrsYnauEn6gS069l+VAcMmah+OzhvxRROb2bjMlhCueykjOT5YQgr
slhwcLmWmMCoMD4DQrCbAS6NyE/VUdQh1czfH5NlYd5bd0tmx31Ob9MZKb+bZX2z
97isxShL/fQIWB2UgY87HcqQ3BrMc7/3APK1qCMF55Tq2zQ+vieCEZTU53FoSF3W
ZdqSe6Zx30EASII40+Ytway581T+c4nT4gbBIC6zhB7YFYdH0XkcO9RsNFYCChX8
Ueo/uaM/I/QOc2UXPzaE0rEI+22LT7lQe8zL+7vy/vaaRdr3qM0t+YM22TliaV2M
hyviVqYqxbpi+31eH+3fP8Xcj/cbyVKVFiB0EitfW6cTGM/5fvwAk1u7s2qpw8aI
If1EwDtzfb6qsn98BxqduTIZ2KuR4Yv8FVDHGqzamkIGNcOi4fAFvWEhFbbnvhyr
me+beF8CHLGzh0dqpjUl+SGrhRCNS2VJpPrW/T+BnkK4J9ng4gWZVNGi+R/BT3gy
Ij5jreqGWqTFQcaGFRXm2oszwYIHrtlRmdtDaUYdboDEn8EGWUELBsrs7l7XFOqQ
s8lGtBItSNhaPFJStIaTLaWt7hXVSMNiP0BeGqk/jQspdDE/nrAygGWzxlyPWrLA
xoBiXzqikaqSC7Q4rRU6rWk/kBXdhoO25dLnZGUcLgZ+1NmvWsyCldRbmKHWJB2a
STxJkl5gni7QbxJ81COYBOrK7RMYI3nQPu4DRVFEYMl0rwRL76bgR1aphj5Ez18g
NDOS7tjryhrdpJc0OLT3S0e91zQrxBsEpcq7IvoqIdCY/Y/F+vLkSQfLJ3FwL5Gc
l8LiB4LimeQwsVxegOFh/re3BHzLT8ixfm16uw8LRD3d2e+sZO0z11R3V3sDvG5z
XWaoM3+hTlth+zIk5mTQpDmxYN7/PjkwCCP4M44GfWSCYIDzqWa/86jbsV1gC9Hd
BxyqGLPfzO7tBWZgj7Y2S8Tk7tx82WzcGzLrgUIs4CH2JFD1xUXf9PMCmXR/+NI5
rIRrhpmGHAZzW5njzyawSC4S//Q2KQ63P6HkdkdHTQ9CGQAI1wQZ8wo9p9jik6zN
DkPHiFHQ9GHzdsnWOUHe/gPN3xty0Lp30FFOCy9nD24gUafWhYWZixF0APayFprS
+Qow0kfPR/n0Ruan7pGThSt1S+2XVYQHeHTda8CAPObrW03ujSzP/3vtJR6ydxkU
o1aI8Sbf8wUnKVfj8gEo6CuoOwl7zgMqUHprmrLUqvqoVhZGiT95SSSYaLqu2TxD
XrxnyIajgeYKsI7PHfWTSGbML4+S6P2m9gQqYRsDhVxNcMXEEtsbFMYiKu7cLkSB
5w4LveA8vm+G4uiOZereGm++Mt3ZbC4Ukc77ihqoo185IE434+fx8Uhn6jn7bW9b
j0hBpSmuwIBsDApVxAEpTujTz8BWygGFg/fxcssyo9rmTzV5kqpbTFjql2qFVOKH
ZhMksFi0sElXMjJ6Dx2en/n8H9YbL3DEqkShxeDU+Omr8mg6SVfIiHlUANHM4avs
xT3Tzw1QjQ2Sif5H56TrSIw0T6xg9O3Qz5SfgCQ8spe+Se7QyP4v+15Yjyb8R5sm
djBrly1uw4NLZZv2WPf8VeqBfHyJmR4wF5u7M3VK1Tzb6QZHbPFzUpFuRmB8Qi1N
gi4hbOXIFV/vy18LFiTvfsam81QdFPnba/6ZHQZhyEcMw5ifM/RIa1mVTqElJxWX
iq/7io3nSFgl5uHtXg58r3H1ty4bjJzvEJG7IFdxdadKd1L/DP4V3/4Mnx4cyS+9
NUJcnD6HOY5pS+o/MYwBMGnidayzO6I66dFduNM2BRvABRHfSAg/eN995KKd7iwZ
0dgvBs1b7m7t+Dd8D5m4W0kY5JzzRL3Bff/WKA1KRpAtcP9H1nfVMPmhO0ZmTkoB
a7Lysgdzo5qF3UVz7Q9VzLAcLxJLVti4/X8ft1T2aad/WdCGlMjat3HAKmQ40u14
tu5rwAIe1gV5KEGe+5ITccy0KeVZRvtGN40ByS5+lLerN7iFEsJPJH8BmBRyIjIY
Fy5jZrmRSVx2MOeZ6eidBxPG9CGW6vKnYL34O+PHidKqHUwcM0yz1nWpVphvalv6
m5y1acqR2eb5DgWtHLgwfqbJTLVtSx7Fma8dB93TUCG68PCLx+pFyKbDqov/reBJ
xYGtdqzxmNo/3uO3wlV7844LLgMEXDBCGOlaUqU8CbC5H0Bl65gfPJ637Bg+eAre
NedaTNQDIRUgsQNlc02aDe69rB4tPragaQzbW8R2D9/6pw+T+SKupYalCjd4YMgY
tNtoqNUt+FRlUHkRlAQaXS9HY61AcqLzPkPUd0UQZnv/Vw5thQYFwwk/0C7V1+pz
JWRY8uy6eISUrwwVVg2nhDtKAXlwZuWJwpC0Fhdu0STKXUa8ypH/DS0T0H5unaZ2
We/we4YCoTLn8SaVPID+Y4aq9BVxtkMuO/i82iVsRZ3FpOtF3SDdVEp8sb9nfYdX
+QhzTxdjgwFiZLuYYk7LCmJWfj88/dUdpkywmdsI/VIroWuoRg0KRVJIK1bKgOSp
AK5gDwKr4sETEbZFQIAsffYtnHOwDQv0goe+V26KWazToipU6N04CHfjBMPkbUJx
QJRgdm/Y1yZCrHDTayqhclsIVHyBV7iXdDaJo7nFk71npZAD88c/51Bv85VuRjQH
mQiKaadyq3Zcbn/SM4yHGFMoxwaN23UtHwt3owFttrn3QVrFSm9Kb9Rk21rAvJoP
9ec/6eaVTSGCi0cd8pDVaY0RgsOB5HPBYyHBA3AXO0kqCSzx7/EA9V59hPa/PzS3
+297ldaAn994JJvOuV+IEVG6u1xxFoO50cwM1KGXwHIJu0xP3/gWOSHdUXLKGvs6
0fKArmlPiF146tT6rExbNMZoH7Cp6dtSPAYncYgsBV4XFgPqVmtLyX4EDPWPb0ke
gba+wVCnvl1jih1IH1yEXvL/xyycHaXuUaKc1FFddMHo05Im4Pum6hb48K2sEaFr
GIU/D68urdpgOfa/qwQD6pVNvLv3s/YwSMuWKYTe6dow60dLHXFD9Eha3IGbeyRx
mfJOr7Zdk2HrJQHWEvrrcAIofBcmj8B06+KGy9HHNjvG0k13yt2LZU60JefUEIds
XLN+t6REEDYRNk8dW9lAOZyGOOhVOcHyw/zgt14wRkfR0DozrolN01AVYl2jIjMR
pUBYLvDl1kZxuWpr9PcHP/0UT8QDMqUvR9VAxJw0VS6UUy8X2FlAlAg3K+0bxI0+
1XayQV8wrwwMHjSxO8OYKZ+IW8XBJd/3SYUWJaZnhZy022PmPYWIN2m9EfVn8Y/O
CE0PhoZLaZOqeiyE1SubHvNqNVQgn9oprQPO67kWFe3uvm3nyeCFvUlyFR+Eh5/b
y4uNLtfU/5VWEx/XTPXi54yMv6W1MvIm5vKra7yaBwRDtZ3SUcWbKN9eLRz2AQEo
g8MztjD6HtPtNAJEHBnEMq9PJ484ZMeses4TTS0blOu6rmVpDWbaKkkMsFP2Qk1v
rSfGa26ARJQPRffCE8iapyCElUfnLEc/BTVJSLpW7tJeVUXzXzUKRjqoN8rKEPCE
dzQHP5KMTIOECkoryv0hMkK63v2zBYXYU224gXHWcqg87I5OxbM4uM3zoWbnbQHX
oRkS/La9ANxE42oSKBhamuLlcKw6usTdespQij+JSighSCsJfApm+HlCx2klglV3
xMNUD6gjXWmwzyklrwdnzYkLCJaExpnsAm1PeAFPJjv53zizkcdC1dt/yZsHPIbx
AU+DhL9GJScLTu+jqJl6tGITck3oi81xpSGLWqNoy+OvormiDQBlKNByARL7qWuB
YLVgFtXrqt5Jd11sCOjVequeGxjrliNWqvbw5i00XVpn+2njEpYL4v72CdMXCyzU
57TB56IcaaclbQ+K72QE5PxtOHPuFwAhkIQktP2E2D95Rb3QkKQ7WuamlQx/bG6o
/aCZ4rowUDczBrHeju86zzxxkQK8zJh1jDjxCHypMegKxvGhBTxF25Wmex769l/j
LMVIiIvVDBiv0ki2uVhZNB4x9bekSJvS/WzFk/N6qbuQtlCcWFWjlP+q3Q3d8Pc5
ycO5Qmq3UzSj2LjuqryuKKBafbJj92ny7nyujWAomDtvM7N/V/hBDjSQMa8+wyPK
XHOu2R8kkJ6OZYKNcdOC84psGWoMTpajD/Gz5rSRr65SR9HdJGjcbIZrcbgH/2mx
Wd86DSqnG5y1f5hW6Um6iGG/9TOi6SlS1o1JlQ5oTCDTBzFDzCp6VrocBqdcEALI
inaiTtKsFBicinlaQvB1N4KtKVBXuMPrMORYRb8QsGQL6XuzzutKvuNbrTnwkVC7
kP/udJHdtX9luztRMUq9yKUL/eRNApzv4tCwMzAVLN6BtfzXHszd4fckoomdGNvS
YpuiAJ4PWpJeoprSmjJn7lJTHKgPnrE0vIbLJun9fDEW+WeYqNdMiOm3KyMVPudy
pvQZO/G1HPXk2hRBZxk7ES31+KISFB/E7NxWpigi7BiNsXy+1IwQI5JCIbZpG1wj
LKiMwEDZdLLy+/meUOgyqmvtL/wjbFMvjCzEEtsBED3jSEvlKkGxsQpduPwO6h+p
T9jD4Enf/HQ638kgrnmXCz/0F9zt+8jaS56CD4epWFPCGBL02UiDbI5YmpvdqS5v
tPEPQNtb73yFIApAEUwNaof+BpjLefArNnZ1WCbe5Zgg1ymvLs3BzdsqIYoJUMEF
hoQ1YsaDD/gMd9qesIK2/SpTu3AaXxJlHalk0AZAEfkg6zUMBOuGGKGr6UD1KXS9
5cM6uhOjur5m26qDzEL3QlsUgyBhUHks1AGdtfifx1LlBCvBExQEhrXyqgiuVewi
UO8dvgu7xU5y1j6GeQ15WVAoa38sVbVWmcwmUeLP9fuByAb6+j2yRHO7ED11XPiI
yW9jLJ6lBvJHI/pNR7HnfQfoI3V4uCWLuTXaGDClfrRyZpg552O0P2hzTOfzj9YS
YrLu1TSr6UjkA4ffH2ElXT5lgtS0BVHnYoNRkNRWmhdMu6zhy9MgKhSyP0AbLo04
uhqGlwzfgBiUJa/8PsyqtBy04DOrmbZ+I6c1O2XhKf0LJD945bIwbaaXIv1NlHvI
Y7W9Z33l8/9vwRCAPxnmQmYeN3sglFrjowgNqByW6RUJG5CZie5oz4eh4i66PiDB
1Ln+YhE+h75MiZS+snZnZad7oED+gyZUvFc32epT9XN8VFverQx+2Z6jPTm+DDbo
4a3/ttsEM/TalgtQrLgGsauMM/G95LTGujRduvzppvyDoN84K/J2Cn+iq9RRtnA9
plynbckcs5MhJUmUr3ywrDiivup8GG6mwdczXfFthgDNGcYiPL7gP+vOUw6YjIK9
Zls2K7Fqpig0twFv8f9FqzesPp4+2c9HiI5vJWvwG+5bEcX0m9lAa9Qkjmvi7AQf
JJ+M620Vg1zWe9kcW1F0utuqLrhSxfyOrRFLZl/nRnVyO2urruMfmgDIuD+NVj1c
3E6kK3OFETI6ImHjaZ1glMzj2UHczsN0hWGLdwhskoMqE1yARt7HHcpiW+W1gYbR
FuMzlVcfqeGAUNZalp4xo6QduGQ3zuu/xObwo5d7XXRcIWAzi96uMrxeJ44GRecy
r3rqObFk08Z6FXbhtuOLyRmTibtt2iXT3Bo719mJgBs3WmAc6HZBIBBgExZY9ySU
vYZuAbvxa/bNKISe2XzlhfuuR211DXWXA4o1B6kA65+QbJ21uhv+cGFsutICgHYx
WajGyznXp5X2cvMr0WW0OVIu/CueLdfBEXDQIV2kw98OJNdbntp3bWSxUL8RWVNq
IegXRr6rAeprHRKtWSJ8RQ4VSiZivPXyzhvKAqcF8Yu4KoTrG5OPZmKoYqs+G+TM
FPyxtqzCqX6IpyU5caJgVGfRDzzD8y7RKNxE5tON2lA/9jVKBAk3CivV8Q9i3sFb
boxzuTy4XB0KqPGWe9/Y0CYkNIzqsAm1DfWFtdpmAv2aeeKDInB/sImdAUZX444I
tqMRqJ7ue+P9jMY68lcbSlYLuYoNinGS7trsP5dz8Lq3uW9mmZ2BuGpjFs1hfqd7
ACONgVvovTakpSafIXHg550N49TL1Yq2230B+OGdkftUYG0HzN1y6K3lRW8ADWRt
4/GeapwvVH5t5JJ1ZqCW8tyxUSAAPlQJr/Ut2sBfy9CHDGHVNC7vXYehIFGLZvQv
BbdRkfI3hQia3qou9UnVLBpcD2hSeh+oRleq8BMTILQ+nLsEYxRJFYkSojsQ2484
dXzUpMuJf8wapzk929Iv6PIXHII5UsdSG+M/WTusnNV6OJb+dmdtTdCKPUabJZrY
3jy3uJ86T8uaGXXQwYjL4hqmgqQArhY3Lv2Lr9ulz4MevPFJG70ntFzEvoGXEK3X
J1yFNxSUZqmuO7HMU5hXJSpaJGRNIMn738bdpYDAEHVhRrsrHVkIhmgod9ekTVPQ
kqoMSWl+Y42MvfUkZFeTxKDItv2ZPPipFS1FJcmoR3rcrwQkrKlYVM0Sq1XTPIRp
NJhdIw3Gh7A3ZcAUQ7hHI4JeJZ5REhvDNEzNfeu/sUa2s2DaZO0J8REfgzZUUQ1J
Nu6tVH594GAPcN4YjqXS20YyB6hUOfi80W7xtC9H480zwAm0qkpKMKvqa4wCqD5J
/N1hudQVpDTxTQ8TiR1vuIdk74e2SE3kB974fIIwuf7WLjPGxgqOsqLG3z//fboj
Kf7FZASprR74+SuPTQQ8cBMF97/dlF7BPXSalG9FeXca0ZNYeTDV8QDeP0tg/pJp
DeRWSFBlkWDMoAO54ftXoSahUagmblkTwFwmWZ3ZwFzlYydmalAyjLQdm8/xNYIA
GmNKAh9i0MNGN90psgpFWDmrIfGjd6hXxWohln0SkAQBebB42mOZlSYfx+fMvIa3
XXhIzRMzPXjLfaBpKzqp4n6EKr0regvR4ww0xNsDEedl9SaUbtZ7dDxxO8PMR6WK
j8F1y2tDDdEsA5QhOqihTDDy3SQfHEISRQ/TH4F8LWqGqpOexEPlXoQ0vnqKy3Dg
WaUZSbl0g6oO2LTt8r4VtbA+oU7yxKVbp/IvwQnNfzyCi5cuhO1H5FJrV1VO5rfG
VyyJk9DXWCdz0TxOoW+APIlkEPc8Mmr/FpOSPr07AFMuLa0lHsGwb+5JFUIYvdxT
ewcvXBnK2ipkeg3ontX/cN7bVPnKr7ZiUpFnQJEtnAbFvSxsi50t24C/bI9KVDwV
rfRMf2k+1gJ5s2vaDx8XUn4w8FAgn9xYRRKoZQZD+jBLnSqj7c/iIfqzKgxhIEM7
895XCXzhVC7C4WAdjuWGcObDkmoDw0Y9KmYtvlZDK377LT3uDWU2T4O0hfNX0DRT
4J0s7XkFTINEoWNcYKggkhQv/eIzBm7xjaifprrQXg7e7wR5pOcnnT/3/4jxD0tD
gMHfRv1/7Evd6nz63fIkN9aPWmFAclpgaHTk9JDASCxZaCxXRDL+FOnmfmeoERS1
2tS8HkAx6Z358lAiNFGfJga/rVe5Lu73husplBYGn8kgrR1+ZJv6MCoxv/otRvHy
041o9jxCWnhxDKv9JQvgDkYu8g+wGJ2k7Eybv37AFw6X5sDizpUwNfSAM+YWvG7v
x+7Q45GWQymot24KJSjAokNRYxtytDNZ6g6z0mw5q8GRT1MjiCR1FQtmpoqoPcNi
DkHDc7fGpbLXfb433X+RvNo73/twj1cwh/7vJXr9UExVHd/HYTHLH9QepnVbkvrs
mnHu+f8cNNm2lnXEVwjzMQn4Ivi8VclyhQzqD7hpFjsWt8ln/n3WB1sHqbOtva3i
m+8J+XyBlQOBw93rvmvgewPjYeG+l/bMKvU+Yxih4wOrzcu6hqLOb7j0seATg1da
BL1MQo+VfHpH48QKzabKpnViwAh6vK87B9qK7X98uD9tTDBCq5oX2RAG3+Pt+j6s
K8BlpqTI04/RptEh4N90R+PgMtXp/WjHppcAduKpkOBrs/nvXDfhgMCJU/EssEkJ
kIZH9rYUCg/u8VgIOKregiNRgee/L4HyRF9gwcGN95CH86nd/Ynk1ih8Mct7A5Zu
xluWFe9cfLgTf/60KANpGcJPirO68rWgW7EofCDHJaHibGn5/Fc6ity9SohYuStA
KTXXbDdGcwhQ4j+Jb48YRyqbRdKaZbuRkpWREgpBen7lfc+o4XWtLd2liyfpPa97
pUbMATZd877mSHifsNUrW05C/1h1Jb8YY6JF5fGppgGVUyQearIJ7N2X0ddYH1Dr
UAtaPCatiMwl6yoOXTqLoQbec3tqRRZEibzfJ++5JL550cqYsaDaMrMGap05RbRM
Q42a7JWoq5COijTw9CQw2YoZj0eU/c8ikaOlAEFxmcpvyCuMVTscus3djcSmZ9E2
I6WtHJyCxh9qOEk3K6cs40pNnpqljC490AcGofhiGlHr4leGiR3NTuLnSjK+FsYL
UdBoHROOxRmZ22IIK5LhBSdv0qInKHByGlnxexSBzyPC376mBW8jNp7DQl8grUPo
PhFiss064AKmOVm3MRimwQPpPyGliSUJVymoSToXpKvgdCYbIqQFKqFdoY7T0xI5
leWpB4IkS90SCZwwnqhie3sguSGoqb8vBRwso88dsLuXewXbbFUbmN/ocJGhfIGU
xjAsbbo0WHCSoAXe+heZ4mylb+QF7MM4r8FrENKYfr2EnD9PUjA463d1RU6jSpza
a3KSm/wT0umgBY36dsK9J/+23Gy49kCTZYhQmqsfo1Tnw26L39o7VL/idrzyTF/W
P4+SX7IfNRR7HIlqooL4XT72dNsI2j9xFHm1hDT11BxLrJqay/YyeYlH8EfiKmjt
vSgRZnUYENXDoaY5qfpjPs5B410gJ/3w9GecJoBo4IniqtHLcbfKlQc2nqQHk5Fv
t6Iy5wtyG4zcZ3nDSBBXQaDnNl0fHIAuE9znQw/3dW1pz1qnWLBGoLHqWOGPW2Dq
2MNubD7jbR0MroxOYhzMdZVa33rP142aLDO/rh+oxiSVArwTsOOmcZTzrn8W/Sp4
NRyo+UIgYfy0EVaMKNuvppAGTcyixqUlvG26PE9/oOOGd/gPm9c28WyzRxPIFCTl
lmM1g/qb1N0/48LEmFcslCuGZ1xnDj14ASAZMNNRa2pPcNKWE6SLi1kHs++clelG
xJwbcMR8QJkijpEwFYe6j2dxdrQq1glmZMW+IeleryoRxtbVoRaTjQee2jxTAS8Y
cE7gJ+j7IO4uh//ts+2udP48AcYEqqbxO/zS52mUJMX9Ycvh+iKCWN8lWIIZMxT7
/rJdZYYs4AXhFNKOJPI0QzoyR8yu7UVMZnL9OxkLdcUN6w5//1NGnhAaH8YC5L/X
V9UpPwB61DeYo1jyAU4BCyJC6R+7Q614vE04r2DHPgKlrvBXM4LAhTbsqHwdvw9r
bbTtMniQ0tAU8NHF5Ov8wm+QBmIcLfXw3dTFg17rVVRvnNpFbVGVtRMcvOg1D2bk
trZ7x96bviaH2SQgNZ1yEiujK3bRgqUVGerriFSNj23jRTjNs4OSWW9dLwCjf38B
uGwrylkE/EAicwitU1DEAzH0DCgCenvNr25Leq1bo0Sl8a1A+dtAV1G5omoEt5kj
Kx9R6NnZP/EFpgc+Lh8i2u1zyhbiF1KQEdBLfx/vXHRpcKhkDsKOQUSWH3tE74Qj
8Q+KCa/izcZ1EdlDwK7KI52f2KOnVQh4mZIWgc8GzKV+/dT+n8Q37jncmxxfXu/n
qQL2m+cfOELQ1Yr8/0sBMlyoXdUPLUzpmLmKh36K41CG/ytZRmuPRhTYzsBLKHzK
yBLgd8UfKR+o/HPK4d6G8ei5bxchKF7j42zat9R7KE/HIw28gMlwFvQDcKqpn4c9
0bOO4MHgGqKPjXnUQ2PLl7rEEoReiegsIw7BDvJSyPxQVMUDiwpGXfDb7GWwGmZT
BHsCvazb4p4fmmi83pQPitVWM9vNWBeadJHi+F7rTDS0V3rhVpMwz13eOPvufbGh
3OwvRtm/Iwfdl6QHT3mLexgE0uFc4WHQbUIH8aYIhtfu4a4mdNlt3jiAHJMGVeVF
CALegt59RVD7SuehEhFtQ5HSoMbfDJ4Du24KNguju3fBLAKPs6szDDac7Kwl7H4h
UD984BHk2UJkBMQUovRkZ4TnHrDxi8jw/DRWsQ7syP3M1foD7WdZsZjJtdstCXs3
qM1jKQGKakVlf8oeiHrYY6oHQ96NOXXDu5/dzF0ZXGjOoPeELnMyk/k1b3Fzo9VM
okUBu1IkYJsY9A0SXjKGgI820mFKO1qAntx652cgJGux3YwA2OlRhQuD6TDfCGkb
xTtyAaSiEAzam8d5fREZH/gFcqrbbQy0WoOXlHD6KmhoBrmPpQji5uvQe8UY4FSh
CuZOJ+mHJxDuo7zO0LpWcxO3Cy3TMHAsrURpfj5q87tFe1GWNoi/wBYLROUmLT6j
e3wB0s8akt3RSpzYtsYn9WNoYCTTIh8/O6mxN0oVNXker1BWO2lGPvj6qVN1GobJ
i/yYs5tCV69v8HHQYQg3CsHFYEQ+0BE8W6PDyLjBXKt0EsjJQHMy3S3mtDHFs76A
VcasN8OAKRtQyglKHZoEHOyRuwAeOQQySP/L338a9vb9Da60/IPTp50FU17mY55l
ijBQaBveP5179+iwFYYQajYFsY6LztjefE/nITxCmr/VpbmpI1ULF07I+MUlo1F9
Y/yedY5XaeMTQfaSKvhYeZMUgOguCMwkwzjHJzx+aOfCnyFaDEn8IGZjO4GwaULy
aR5JIHh7FTUVUlnncNHa3Ur5IIbW8enFt9TOBQKqGedJkVbDQn3GspjRagwVw1hi
/2lr0jI5AHbznLHm0c6k/1sMulwTFXKN/NsdW8/BtI30ux/ghJfThZDQ8XeAeRt7
JECxZdAoox0FBiudA4BD1VOeCkMgzSQp9ZY82u8aHAuABjUpN47rjYQ2fHDKomrX
66v9RN242kHAF80x7/fwluN5t+/Clwjq6pmYY6TmazLfYwVzY46XCG5j1b7NW90w
2pY5AqbdytypfvL9Y0fasubPsBn5vuvZdB4dEXuUyhUoKAwqlnpMe94wt5dOSNb8
bIOeOZic4+aogExyUpKPRg0vu+JzpBCLzmvSVMvzNgq1VbOuOf3jNh8+k5cqHaWP
zsx9LJOiQhS7GEQaDkfF/hB8v0J0TcCk1n5sWABDvYep8LSO4VxSFXiKOM/9ubIs
eMXiJ8AKYN6YQzF0c1Aqmom2S/fqlQutRBW7J0ez4iRi2UR0KYURR9NGWBofPS8o
QcFkiXyc+XtytRRvmrH6Z8TGEMs/77MPsaZpewuP52tmC5iiXncgkNhVWFIwGVMO
SMMUyiLAnYjQ8flVvx5ngouWCpOR5ThicvKcJ8M8GbtrdKGYTyUY6aIz8cpgi9OE
thN9gdmNhHC36BUEFLxRSSmdTytDiqPGq/ngBB8mTTnp56gKD6oe+5wjtwNf34Y0
dAdbKirZgeey/jXrzOjbjoNyICJebHQVy4JOo9p/ZM3Mne6zFE6TUaj7keuL3kFm
8bHm5XvFI+anFR3zCcgYwnRTBytwXnL6NkYHqveMfg478wiMocJy5GE1p+cE5e3Q
qFwBwV3HFwb12wGzdsVt+gAqnLUBjKp+GsY0dcRdUM7qi/7jMXBB5GvOD/Augne7
4kX3ibWZlCTUqozsoOXUU3w0n5YhnVMgBiy+Rt6WhyLN6CYYzE/r4ByI1Xy2TPmq
Emdh2UgMNEXSXd6wAqptCdLHz4bp/HLJgpc9RIQ1AYZBefamlpV+bctgM04t7TCI
soewVSIHGmRrHlixw96QNmkSTxuIsrJhBzZlo8tqB6xlEb1HXVnItgSWv/ZoWQM8
7q+iO1tmIVjzcczmhiQZMqsUQ9aO09Qc2ogI1FVmupodulYMbiEMHKByYvXD5boe
pZ2Ob9IqjMZqYCePdDNVn2+f6zZ8QViNhv+vmTwuaNf0SzUweI4bll86PlipUwFJ
ysGQMy+eHnBXgzpcMvYIkivgC4yrMy8/S7y/sEJStHQ2Tl4eSbPvj0ybhX9lefi5
TdKjdrdrT7FwLUIt7UngyyBS87otiM+/Rj9u2gKa2ZZJ1xefs6B5TJni23oBXM2Y
ZtdwEeTr28HwDA8sWcctmaJTAN3vxDJ1xEl0JDvPD6Hj9YCfzWCh1d9sDiF1Xkz0
74bKBO1NLpi3z8++PlC0axRwL45arspt+c5L/jwEtK1HOuDqv8sCQENljQ+7CCbL
Ha/hjfZ01B6ztKEc0ErrQappIQGEZRIWNdivDTmTPsf1KncQzyxHHd0FV9Egr6rh
oW05B4e3+91aztHmGPjb4fyWJmh0BVFS+F7Z05AIAL8/dDHM4edaoyXEN98huuRD
SS3XyEb4RVfKu904EhUDTHURb6rkx6l90JtZf/R4gH8qmUNeFOO2RaVMvHRty9k8
dHD1XzpfhCCOXsMX8KL/sOCUBTtEAG8cXL8M7pDF7l4RCMj8ReneD22RNRVFR6dl
o6cmCQjZX1FIJjyh2TRcykqqMC2+4XsUebuP0xEqzZMPDcP3EWVVOGQtTKiK0m0q
XU0FL8eVu2VSfxjiRSRNIcp4V719o1in3tn3YRlxEeS8Hy01qZMLUOmFqACFDgKh
K6qA311g7QAZZhYU8+8AlUcoXfxzQNn3FEMI2sebjHjygKtUcMJLAawhJ7SdVCsz
D9zfwDDdSY6fjzsYqOTLVqWCDBKXi3+29TnIPYoAVWiYh9gE+n1ucRQRWbxv18RD
UqWr3ySXaJNeYfSqSinpTN/1+0elV3YH+GM9LCXXWj3tNDrep/r8auACPG2P0Kg5
kB1mGsneA0Rly7hWOG6kyqSe+X1lfSeqxJlDbGWio1R5FJscEdxitfYw5BUVHzZh
31Y7cM5VrmDyTpxcwKsubOD9LbIJMUInRN86Y9ZgJeERZ52bt5K/wJf81UWYDlHW
TzVahkNTLqBS/0Uxhr4DOS1XMhXm/c/afCpZMzLPuxoMbdCbvm3uFtSwOT1jxLqi
MOqHpkk6sNZW0D2v0/ym5FesVq6ZimDQ8Cr7mA0KM0Nr9Q64C4UppUpIErAKkdNt
tflYbfi2t6x/M9LHIMAw9u3jT7FaRdOeSleS/jMLjHSSwvZdl4hvT/qYW2EnuHck
kdgNHNyLTMSf8Ds4MMZljP3yUf8anDT0gz/8mHMbzMWn0ck9QzG3cwAXEzXq+2bi
GPHQnvsj0efDLN3q/a5J2KFxTzFEyh7k3ydUpDD4Hhk0lcUgVJVd/oSRcYIzbZNo
XAp0BQhFLh1zexP1Ng+HMuN+q0HbtotaviPP4UOe6vWF7S3AcUrYdQyG32Wf1Cv0
4MILEQfOinSldEJBg2d08bgcbgS1HbDMSN1OdZoszwqYJEq0KvSfM6TPCRrgu4RI
KO3k9KF4Bk+e30gtTzunBp0sCYreSidj404/nmzvwWyMyqUz10Uc37q0dnD7Dx+F
hrMqAk23ynlDWJpo84SCPHk7WVGIPfcdRRzvTigSgA4Hg3HV1sfIfcQpNcQqULx2
+nyzuzx6X/+m0M9U5szCZhykJCrSTztX2+71o6MMUUcA/8JpxrxN2aD96Z+Dnjmv
6HhKSL/HeQ3sKdA8LNze5G9YC2fyepOc3bJIIWMLi0azgRZ+LiZJGZ+p/OAHPIhY
ujf9b3U9HndMk2c4QpjOLTq/Pf7rAKVXSVDpBRlv0xF3010+JCkaZDADLkWuWpiN
4heuAxo56HnBkC3sqnpzp6FMLLWEx5OL/7fQlzT0/J4Xfjh+xk9Dkej32wJNsTAs
8eYrjkfX97gaZw4wc9AD60qrmM36rqcyc8cLIbOMZhGcKB/VcdI3vKnViOsrHRqJ
vVcoHMFOnLQ/tqk54z//IVwT+R7vyLJ8DxhWGXK6LoRH9YFK4l2j0bsCFVz3BTNq
r5LFbzyWxMDW4HKAKon76oDfT3NQCgqqe3NHG2qKmKidowWr+mDd2msAMMmkq+yQ
MjMXPcZBhIhOMKr3Py0c2DpoQolfZH/zrJZZEJSBkppI2Bs1dg/0pENSQS4zWEwY
IwV5ZB+qJHzs6rHQlUxvsBc7AXYON/Tvh7SReAMBiSY/3/6/tDFcGbyP1W1RGBp5
CIWFiXPJolP94YWWSMhwRU3368asq8Tl96j13WMZ9/ffCl+RIr1zOxZ5Y/6Jom1P
wN2MyCC6lhLVAzYrA6dpAb01RlUe06+690V92FudffdF6iAZqGsMqNSWVyAwN6Fw
p1jsHhyaMuKjWOaZYoyS/m1gR9UgMhQFnTrfEz9j2AEHx7mmpqjAfG3YoqLH5D8G
2ZB8pR32LgAZpS2biH4QdKNicdWR1916atxMGFqV042R2rv8jTzs48HUu2DZ2aBM
xCTISc1C4bL5NsrZjL0bEraUf1B6Iit5r5Vb62T72LyDME6LaYrQR1KzkKpMGAV1
3fJTRWZejDqa+wOCzEsXjW9lhjzCSqh4S9ABmfbfB27GTyywoR5yGXSnzM8jCRmg
/ntrJiLqb2m9sa/hE2+TeigpwhZ+uAq4vtvibiKKDlfzQk23MX0I4oOraxuR/gAR
zkoy/h5T1D+B42hvCldrsdES2t8hqXt0BHGnFqUvxkcikD5avl6t4lJaDSBM7Ytr
qkCrum22KxOD5UdKEWy8CXVYn9YM3o1FVVnjiPmdbRWPDCFZFdhNK3wUZ7yXd6dE
YLuo8/tzMD9txGmEPm6rLFOv416ya6BZyZ4Q9Vi7sINeQYqPAYhU9cGff0RAOvUd
eJMForcMJi9mGs936r3BKIDRzvlNkZD/qJ6DdDPu7taao2F4Ew1Ilfxa+ZTSfDYW
etCQP1koRTojO6wQwbhC3TARLTGlK2+sjGsjEJ4P9wokwX2LL4PwS4BEpLeO2lvB
ewu3wtPKfv+fjVOhLTf1Lo6YcI60WAOWyAhbY82CVafvuqnzkfN1xl/V6q8yyOyq
rzTGX+raDLV/nboVI53wg0afRRRRxarAd29XOjvuX48FpgJKS/3BxZ484fnYB5MG
VeR8M5YZ26nUsPJMJIs36rmGepBgtaz4yfuQJMkGud4Jd8wlG0YQE5q4H+nugOqT
fJGrzqq32RiB/Ja8V0is06gfRSAv+E8VZt+liOjWH3acEJtX8J2UBIws5vqFYVRQ
5z5i3tKxBay/y+TNtFl+1QvYBCMyX9zyCCmElC/qfFv/2xgrNV+FBdV5xa3zKUrS
9SKNC65gWEdo/U7E4ycEi3SvjgCQjgdcvwzWo6UKA6UZdJkLvGvTYZaHKtjaTGsV
/KJ9jJ82x2diB+roGDOY6v25vU4R0weBlmGMGsWmilGBKJrPTHIbRWuRz8SeLri2
Si2KQ3Pdp/VDTMS4JU7bOT3ABOwkzbzGUcLsw1GUQC8CVm6TAdBA17i13jZyAWMU
yAK8C9TV/xfCfj7SggG8kLoR73qdvjJKksE5/MBkdjVh9/cnZ3dHlCD8atxIFSv2
pQI1ttAJZUJ0apGUQFB/4RFsOw0I2hJDuNdW3X5wQ0U85uaUYUIpDntjJ7K0KGu1
gIc4H8LIferx4ZVBXtwUmUBHDeh0r0JY2z5iTNLokjk8cPZTqXVuwV+dgNqjejRy
ek6vimZuXV0btqDLrcnSc70RbtaZLbvXitLbw063eth+3inbCmGzXwneVHeP7Giv
E5eiXE7/pGkDPMJrRWU/iHTvgTM1aOEtRWP+4u94oW3d4NSt+Km4aEYhPsxMk16R
Rt6dYeQg6V/C5WKlRrYzKkMPqFsMqURHFuDet9yflTh0QEPzsGk22JwbAd6eecZ3
zoAAukWyRJSzJj/L/LK1rsHUhxdJc5V17VwncA+URAklASl3yQR2Wq7Mlr1xRZ1z
IBTAyGLmcUyJQPLC/XsSWP+NX0OSVEEso45uN+IBPkh3NLEajqmoyw3bQysxQ8sG
9Gulj5r9N+9cHOYBPQzXXbs15BfCIZOnitPZ2jISMcMwXrv9zrQ5B6yl23Ll5GUc
WmwC7FGW/OkMpq2gfaMBCm6esOH2Bneiyvx41Bhxfg6J+YCiSmMtP+RJyIELxVDL
x8Sx3SynCwfaDEDGEB8boHXt3CqxlbC6fFHLl/JDE31Qc1XZSfVG8UPC5RPG1Fo9
tb58pRUD7b4ShUpxSZgVlIVUx6jt0o7V/TgJt/8YKhAEs+eFg67efQLXQ1gfkXcg
cmIXY48EqHOzzGJ/ImO3qXbTds8XUdalFTHw7tg9xlLY9uy3MyxR46zgxRIWdgSv
WgzBgArPOuu4U6Ch9xyyLTYgnvmYWuivnQWDAqmjPbgtUI/iGomUO0Dh0vUcdmVf
kZagqvj/KdWw/35lggb/d4K9AHBY3kxCTDbtz+Egco57Nd+6tb2vM1oy0yO2gkcn
/RmzQHPTESHCG7j9BjWAH46aH7MfaRal17l7nx2MwjelojQkwV4vIUbCDHB88Fgs
ZW5RJk9AZCUIUkoQ+QW4tnmhu0TLnRKqpPTcT1bfJiMICRnZF56sjT6lsmg0URmh
SwfOlDtiARN9aHYddH0WGSiy+ywLCZXurKmC2XxMGraxxv0vySG23Gvc0bxzG1r+
whEHv/xdD+ODMycBFGxDRNzAvimBXRCUZVJi6nqoBAd1nU8/8UkWvyFNW0BP+KQC
0RxTu7xQIRpYb8W1JG8VEduj2QKxM9W0ky9pDFoOUyxThKkWd3kwiOh6b22mw2cz
T6zVJLY6gSxF6O2UTkR/L6NXJVpA7HHx1TK7R9kNDjLVJNa8zuN+naRvOnN3XOdy
v0JNIcLfjlefgaB3qll5nQKOzihLVYAh59kmSPTmYc0G6tXd+B0kdrV4ssEbjOUX
waWoIZGDhAJzM6L1PkcUMD71n86bM5t7far0p8IK58p1b0LzTHibhl43C5myYCP2
U9tol9veYnwd8u/0gHyA4MZBXocYWRyC1IFvD1MiWkxN1hk7PfW57DaVp04dBtl5
S2bA87x2v11Jq+sji1961uFzr0XjDu3LwVKw7VQnXDwYVJSa5+VqW/P6jEQHXTx8
N2QlFPx6USIQQgM5Q447pdRkxloAFvTev/fK5URopyiKoQBc+nCVLBjMuoLtddle
XLWpvQAXzbUXzwQa/cdj9p1k3tB/vXmjvPnd5CfGoWdpqgRIEv3RsOuI9W7i5/gl
Kz/uwrvnnYYSSVVm8daMHCQXeOU8RV39SuaI0+skWOVcSPGZi8jb2B9GqEfsDvy8
JlRrQbRTv74NUSvQSXkSY+GDmHdeFJ4a6YVXnQFgtHAqzsZ6q0X5S3dmT0aote10
bIKCCH6YjeGmT4JDTChpz6GG4kTPAc3mUWUjh5IO/7lRS966IsyAC0eXf87wgMnU
IQNJ9g5HMpA5pOi0NdTnNQ92xFoQrqjmSYm1DvmxIEvEhZ3HI2j/3bko4I+Un8Sd
gepqbVj3nJEi3OYi0st8T3WfpjY0izLpB1oyIXheAe16FZ3wRT7hYJJcpztwsIIF
o7gBy8dfc7nnrfZU0/fYtqjt536qQLbSZGAyUonWeoLU4KJUx8ha18tdYQsqEeVT
n6A4SdrsfXlquHSKw4VuzwE+zaVtHjhVvoQJNS94OA1MPNu90STwMvylmOTKgu4B
TPk1m7qca66QK95EEH5fiLEpJKnePN7Qz1p8mv68VM+3zossm2KbV4HDU17NS7Aq
owgmSNFqwmc7ODq3iNjcS5m6ekEm2f/ZvSFyidUAjsvJq5K98STuD56/43ajTURE
nWyOLgadvahen45l7vAL66+rJnzLkSi6Hz+HSwiriLi90PrMQ+HHPmoY8SFo/igr
UY/EzlBqcfDXgfVR256z5wIWMjO4dCMWGv3NvOvV64IY9D4uyUeARL8UW3JGbDo0
EEDhnyVSO9+SDNyRdrfvduVpN7Nz0spa5XzuDscc0Os1CHDOBqxl4UNhLZXvLCRn
oFqU+FirqYHnDbNP4x2dMwjankxOXpUdxESx6UE4IkTyTDpwYU9mVzC1Na/PMD1v
XrL240/x3jdWMyyssS69FRH6rr1O+gSs51d9jWtvDvm3bfbe2fawLPNTUzDk5IfQ
3AWQ3AXb2Nnp7DQgDRY0QqxCTwPxYUdoJ/N2vj4e7QGQSp27eQ+n7Rw1Fxv7c9of
WI8Z8jMsUSMseL8Il4U7l8u/wBejNP8/By12Qky2m4rMg+ptmeI1n7gMxLeWd1r+
qMeCfhXl4DGj4F7AGdxX0dxr79RX6EeAaX6ff7bS6HqvfxP9ddG8/q6gSoWd+3zP
anOFxNING+zP0ezzD4nL349no8OcQQWcBiktf+zFu2RIFlvivm6e7DYqSaHNWmbb
J9VPpUMaZjp8bY5i8WzLplALFhjg4eRZqE58yTdR03/aFYGj3SJPoVqNpjQ5dPg7
HYVdgYtUVI+UEW0FYMEAUG6U2xRqSq8TrsoUD/XfmPgDwHD5rcN1nUeC9QEle1TB
2b3BPudB86KsIO6Y4mfYvcqoHdAOi3mXUVpKRuUTFKIiSJWpa9t4JCsu5orv7r5J
QtKerX+z3HOYBuEqH604LConHbF6CoECq5iyOhBILXWopKBOP16o6EHxz4BjO58l
U/YRXCQMRKNpnE4E2sWvLg3aKKbvHRSkVXmcDXztG7YrPjZxi/S54MQFCEeWRplT
ln92raTFWkFVBxMwmSDYrqqIq7Vvd/iRp5yIlaEPEKIrrjfy3RHXOovVR6f1p82m
Sj2g7Lq5GaXkZmDrVRWJSAsADeKWTD/niX6OscwnwVXkqDNJREqHvnTwY5+lG4UZ
0WGVv0YnBxy6nLehwP2DfJW9tG2KJMj4dZaF+btOFTACGCEopTM/5velivzhLu9D
Oo06EhVFFuntdGlxA6hDqHJF+c6n5PTokp/0G4AplNO1lRBEZ1b1uDpw+8khq7iO
SDT8i9e8Viues5VoqMnC0PAVbXo8J2UKWej5n8oNpkqRA6bpxPf/O01H4HV5n87J
lT2Wjpg98/snagp8K/ome1FOOSW50Sm/d0N53SzTNhoqBUzeqzpW+RHVA7PWpHpZ
yxKU925HW8EzIszUvjrEWhSjrXgzrNlH8Y1pWVz0XTG5vRw3qTuRXh5NqNH+odhp
z5dXXJjqF2TuLfLzecXwFquW81h5H3dSXG5e2AaHjCLd5Kw65vXdJUG9Ls8HWMV1
nYwn/qG7Rhuy8XuSOvq6JXketgFTCJn6u0X0ZYrTnUZNxKRr+Lkkf4LxmZowHQkw
SNpAsOb0qQTJDwCiWRXMs0qmoUDlBvVw3j8Vr2cRomTRxv9GsmBTIeVSyErNPOf7
DvEJcO4z5o/XCgjrMlu8PDTPBK0YX9lsjuBEFdw2K3kpJEEQNetOQOPJEoX7Bhaj
7UfOrd7U0AiYk2uNWqdMPQB4jjPOBcfXDTccxUEqGurbjj5dCF4Ik4t7q/ccIcOd
IsUKSY4XtYtwAfncWXaf8YawuNkaw03DU7lVZKoeYxpP68gdK96/zirXg2vIIwSM
uE7FkYYtYE1NgSApIg25W19mEk85IS4sKdWJK4zwsw3l/E5mdNG54WmT1SQCkE8/
SJMMHGsBS569ATPiI2BuhbrfmRJDbHiltaI0WbmhcpuLyoRXTWzWO/0y+ONGaLR6
TjhXLkpXhHc46JdQ4WQoi58k3PSBRPMX9SDJMW6a74LG6uZAHD7pGtMehuo7KKXG
Bw5YkXhDpUDsbhjbp871sk60PRLz2Qb+UwQE3MCjBB+rMp0cyd/T4Gb19iBnvKzv
G6PSOTXny521cCMHQ0xPxmvZz+q4/GsrNxjl9BCz6fDc9m2EmeWU4uQXG8CHuGIH
aKER+/hE4lL7eIV2lvtx+IFLrggTt045ONTWTl0jB6lf732GHbLxXCzYEcnpCxdW
iQk4YxhoRAj0tZPSTvmTE9ih/YON4HP5idIH6iknTiM/YWuhn5X8zbYXoAHz/H9/
fempdY6uEeEVH78xR1yrEGLA2+dojo7kdupiyllJMn2vIKc8tgiLoDGJNgnCzT8e
KRksYxTolEVxm9/gnfUF5YhXE4eN8yb8JJhI7E0DZ5cbRugxoPueHY+kK12ddkHt
4hX1GRxS5M2fDyOzyfR/vRjdLLWqqvzFV0cD7EoIXzgFEyFmA05Y8Zrb6iwrzHUy
ce8PfIdZnB8JzyZZbLZJ5EMHdGXs1VblAXCUKaytq0CV0ZUZ0E+yQlEaMGddStY+
Sq3qsGnbYYICsX7AnMW/u7tZbEqCC0SrBD/t3gbl118UdH0ZiKorFlj4AyjTIj9j
LEXHib26L+nY3cebCOV3chYKQWUhh0PW2ZtJBzCDuMkYHCnC84OgWi9Obt90QUKS
C0movE+xoOq+aJgi0tddoVjppcEwqE2L/v9C2O1KgU58vtQOGwFX6US9ASEni/sO
pU0OXfUQcP3E6Rr5k+g4hWtFYrTIvmwHPRve8ZNv/xnQ54HJtbIzSs2OC/5xNGdD
vpAbDoJyP90uLbQE6FGuUpAYfocpHyI2OtSz5nJde6V1sSNvbITe/w9DXCoIapPP
5zry+IuGFqzhxlgWFFu8L5WOzceZ6fNpCQbLqjSdUi+vSG25kEATncDQOGp8JylX
Mo+96yh6Y6YarVrs/s/f7ExPVama58yeCqbBYkmZfjB0TaFu2DROJXDk3OpOC+UI
T+tjUzjUs+0EbgSpev7DzWQXjdT4mHD0+1L7TT+y/ToIVBNKWA414uYRuuedl/9s
eFtF0v9UqZdxMNN8YdV+o6pObnn4xwZW6wmnvY67dKVaNcReXnHK+1vHmyM5uBXS
y7J4dcym0SNGNGBU8GvDQmg0kGEtMGZpwUxUNWIx+VLuhIuclbR5HaswMK2D7Yqv
3s8WCLu0TPHb/U2hRGIsLVymE/kZKN9oGd/JHGxCX+Vz+koH7u9MBJnUjLzstl9+
KE5PH7Zr81KnKTKyaqohBbxl5s/EOe+ttQM7A/aVga4WhExop2lYstWZlYWN2ASp
NkhOZPvxVNhDINXlfotnsnlLdng8qPIRF5TJIiPEei2ys1X7Gcml1Iotq2HRqOth
3fLtmkZLxmb1rLrbYqVG5GSgABhn3Gl9kvKlRawtc+fC3IJ3TdtLsWMz3w7lj5xr
l21zMJRO5OG6DUPVTQTuxLQE6ZLRMaREmtsw9u1nBzL2lz7KRrmccH7nSnWcAcQb
j48jk9oMgeLLp54tbQv4Kdk5y4knqmsrIdQnMwOEHWHO6l92m2uUiOksYFkXOdsX
bquRKB0eFSmtFjeqPCbDh0ad0aruzmwTClQBXhsa4amH3xIWd23ISpruZQk+pvHj
fIgzem4uNy3FebhGYwVXWGqoe20lX3Uw7zycJk/2rJryOudKcb2Em3DEuYYMnm7s
fl3O5R3AkZNYCIq0mvjxTgW9JSbSJGWy25aheOJlWBOuF+ZUPqok0UXvf6mOoqB7
RLbdW2V74Zu9nUeTfcpBtXTjWvnro2tgHrjR5ZZYfUeD5EYhxTAm74um2jsB1YbG
9di9gvF4cdUCR18DdMudx+gWay3Wbj5YdhYx0COoBwlF1YTYskCFrH3ikhz/UyqA
7bkeWmu4CPcAw26Udb0xPxfWLGleFniGHESJuKOuUduHO8aVIPJSBaubX8Bx1846
FBkijZxBZLtJrwnrjC1V3lLoAlQMVr2JnChKXz1EHmms6th50onoGm8TCX8kk7j1
Nec+wymZPN/8dGxJ8yBQV+8Vz6V8olgIR2qtj9DlrM7I9s/1PWT7sscsTJz6Q1Eo
ASoZUnKIKJusvaH3oAZeROjvx7WwA16rkPvWz5FYSzUldrRPrMLt79CBL25ZzdH6
9ilkYY5qFwUJbjITOGdB4rNHt6tPrwAEYmTOfYcxBmP2DPmPlhVNmM0vDZV3KRO1
g30WHpZ2HkKt8Y0Uuk/HiksJ2F9N9mzSYmAhWjYgz3KerLikJj33oFb3+MbHHz9b
VvJzh3hOGvlDm72QB75qRW5TIHt7s6ShRLpf1sed0RatPk/hqNmWerC2sY35i5Wo
qO/26t9T/irSCSsPA3e1n8hr/4gxbugmgDYoKjCxSSfA5aOaJr87lxnwZiKFdyEk
eWNMcglPfPTfKRh+SH0JG/FU95HEfMhYwF9PyuWaPv5SWp4zY8WcxWNW246uQr15
pwDd91JesYfgH5kXpGpRdwJQZ+nsnBcwTMSukFViJKpmZXnUrntuQxBnTvObcqca
jT/fNvcF+jlZSb0XHhHBMoTa6yVRVieyp32mzXd5sCWC4UiHML/AFm/rV/+HqiJg
+jkzbTCrzOt48zJulesNsNlwLboZ2309Gr9rOt4kS/KMorRTNT2qwxVj6F69RMs5
qZByxkBZYL4Cch6qleyXxvjkFxfiJ5rcUTL6mEVLWhKAuqiJJ6iPEqjrk++iFbgj
BUfVHxQwtZsTg69MQSvpZoboSjtCb+BDRaRd30VyAv8eORdYem0HUcR7N7RClw/V
bcAJ4BLCddu2ooYsKNfCWAnGuLg3DSuboFuLNvOhMvCWQIibhdNGFY6cfzQZoBSF
zsy75AeqWXQ2ZwWIhXdembgykLbwBwjPGa3ooo4L/zOSO2lEY43tikA8zVy8w0Dw
vIv+KGUvV7cFYD7LYVqm0cy+rIgWtfWCCUQxsVBtISYjXDESXSCXILYBR0OYXjFG
HX2W9WM0lcMh/C8BairS57j18ZxcKyr9ckrE/wHXMbTjDoDqlAIqnbcESgGckd4N
zUmqgX94NTcdvzGFhV0oa2uHmisHBG2+Qk1LSVKH46uOjnYqhLGjDh3Hel/PfR3f
D4ujwWKsWC47VbVaXO7CUV1RU9xDeQuwryo5bR7qdCPUlcJxq4HQF8fZvUVOhNOn
3wvWVxUS+tmd1JE9pssnKcyqSmqelj7LxgP9ULNa9aUmDnoukJlgIjh5rHGVRY3y
1r1fG0HLbOZ88+rTZ9RApY8qeYirGbx1u8LNk8uUpWLf/nb+RpLBqdIYT8EKdcWu
/i4YRnHkrg46GitA4GSUnpTKvhuxOar0XgmanB+pZLBRPDOZpuP+FdXRkjA8Y9aT
lrD9gJmECQ0WLnPAaeVfhmuinA1h36QNL49o7GbAFxpkH/j9PECz/ruXgSaAud0Z
TRsHCyD0LevxIv5u82lDz75YCmMnpZIw3pjSxkkCG9UpygdMoB7o+fHyeYH1C1rc
y1rf7vCnlal6q7yXKdcAl/ucpZNbFsqN7PrxHtNozvaVUhF7uqyllUXNMpRdx2ab
w6R3yHkvpVvanSXebuBn4IM1dZIevGmTIwVdb0QJoj18jAHqldhllAuYm2LyGXlH
zahoGbRro+8tUvZ78sSwzhp12Gl/8I9tkpr0oiqQIlbwfJ1Gd5EVhemuJDO+GDWI
0TxSqVJd/61y8JgP8yH2MvBH5qIWv4dtuM/ABtQrFP9Feiu8h2PXnHwpD05kulx1
S3JQhDwWXU27iycBylaSh5L26mov+Vk80bdV3CgiU6z/meZShxdL776DGdhu44Xp
HlPxagQAAM5DWdl/KK3APxfQbLdXAxmHRXK4EI2UajIthRsqH5m8FOk2kP3r6IRQ
3iyianyMyJFtIEggH2OkyoM1d74jqLVgtYSjCE6oUqR+UuU5FHNTm6kik3Dds2Ke
X2J+kFh33dW53CVhe/XtpQSonKZ4Elq+Kx7XfqIOrOaMnYHdXv9xmBtIcsCfuOVK
kWwUIj/XrOMlnFjZf5CgxR+FFasLC5iGAPVEuvGuDV0DSEaZuKyrz8Jrr+4fbLDV
MnxTfd9O5CSicderZNKkNv7Hy5cjmBy0bQSWdgi1tgKutA273McArWDjtzO9//CD
wbZKcqpxxz/Zrs4hgSG6kwEyIYEwG7R2fDTJhx2k37OXYqjna8TRF7kh7TBDIRf2
dQ9nU+XTtuV0R5RQ2Gog5mKR6MAO1Ink+Ys25HPtp4LIiZAQLNky3HGvaHmLW52U
57jmifcybkb6Nkv7glm1I79lEn0qBs+B13ibE0Vmec6G6aFfA+/qy0AkYiQT8Ubn
yvtTmS5NHK3LbajP4Yep3PQJyE3mN1DkzOsb5749KWX8/RFx1HNGs4M5PchsD8yN
5IaSc74o2xDXLtTweR70+KftLi4ZZ1p96y0SMktKtkf2pMa6j+RxaCeZ2VPGqAYr
h5fjGqLvHYTNylw4PYWDt0J01xGjHEfwXaf0cwQpeHdppkiMJ2slEAEIkVZH4Moc
8muJmX670MxQzmwcm1e4Fz9VR9jhVyWQe874j9GqG1GpEJn1PYbcslmRcKZ3670D
c1V8EjqfMo2xFdhTKP51F0AGlSrw6eJdF0uXqsH2pQa8+9RBgK9YKLVxBWWQsCMN
fZ0Da4eNyJOHU9yEyNNRC02oFZdlMgGHHpfJ9DqNJ6NyUhnID/Or83J35IyTB6lQ
0IN05TDx+yNmGPjcC2ICX9GL9nMCVIP+4h+49PMAjEAHRYPxlomnqy0gx7zZOmdV
tx/k8f6AMuxcCVrdGOEJ/caNMjeTk4oxoQmfJGqGcd56S8tdPJyQi/PR3HHVs/wc
9Wq3vnWcpJRMD63bNEyemSsGZUazD3RjruJxEXoss+wSMzo704/N9N3edUbMk8tP
40Gv0JMdwhDCdNKY8u7l5CBHlQKGVaiBlsmQSeYya454YTx4VXmr5HV+umtcOBq9
9uvW1+QTFWvOomhkNroWffsxk8Gx41CRgrX79lEjb8ASOqKVzuvbAOFZMYJjkq9z
hqyzxazd2wKrhSTBj4b29RR2Wva4S079EdYxResTO1agpUFLvBuNEfcIahNt6f4h
uPEsntlowxlUqKklzBUiZ/4olm7omCj2nZBzi4pMXkGLtmZ86XLijU2854olO2FM
+FCRBm1G8cELMZrwFffBa2s2oibWnskzXIQHNnlR6B4B+lGfzBvDof4YnyU96qCJ
6fw+lkC60AXorCfWZle8WGfIKDYxKdSJsOi1m/UcQcbAFKpqXpblWeoFY5an9VuZ
9Y7J8VYaLpgmgnak4qvy99OK3Tg9z6hmDe1OhygQWjBmYhOUJKxa5VpuHb20Pu67
ZAqYSWBT7UwEtmj+VbAKSvFbt+cvbhDrBoWkj5jKVkGuanTGv5rYpPkP4WwM76a0
eAzCPQ5BRZ2lMAXGPynN69JdlObve6f831kU2pR8E1vmKphSAKMnecIdovb949vC
QGieZ+Z/MVA1F0OBRE+HTlNX6jyQzBZEJfWkywW82k6VLQHzfV2SXAMj3YGPKfsW
+9kjjtcaN7MxnuMh2lG4oDZHUSgUJDiFE5MEXTniT7KaEgZCdnF8NXB4HPief/+a
F6O0sdtFUp98cSJ2aHQmBmqnpPI16TyuGM0KnRKnCSkkd5B8za7weGkXCpRXiNd6
NvCSe4b05tELZj/Q/ZsQvcZe+TMD4F/+rqFCNac7yDirD2rFY6eVukOMOT1MEJN2
57gIQb116NGLj0T5rl/uLXTQU/NgfzsdWOGON6ErvgG2IMH902klhfMkvl2mB+YG
KR72bpJin4HJdbaXbk9nSgkd+1M5Q2H0VA7q/g1tBBRww6loRTzRV22HDLAkmxQO
9MVTy9GWXcBViFRpE7U/OTyNGq1WgDGqpMFTpr8KNcpUc8Ut6pIiZ1cumszH78+Z
44Z8gGYBqT5ap7iAkSQTICPdWoW95RmAr5RaQ7lweFjvh5O3uittUG0ra5RYO2OV
2lDXweJLcu22Xf8m2ESC/vAWKQaJJrjr4f43yLa0xwbnkHrvw3McSlHo4ScdDoTv
StNmlAZNVwfQHfjiNWzwZsUP7uCYoPUdz3fK56PuZ9XVe+aYaombEWLghGhRUp88
w6bLS3xW2hV7VP0DPs87DFCaYfuP+g4dr7e6DExI7l/53SkZqQbYpa8kFusG6jIc
4rNtMjOEVnKTnIxI9+2hQcLAhPdmKlQnDA/Rn3BUHeRpecbWQl8ZZEnXBeZjOaxo
gqN/YH6rq4n6l16gA3qgLfWrRKWm+RWN25pcCwpeG7tTRjsfbO5J2vNY73NExWVU
lpPaUOJlVKckUHxgGPkL0E0BP9U/X2IisIHNDcqgGkrWvz7h7H08keuSdqFcdYAh
BMtCGZ2lZ7cMRhk+M1q470X4soMiu9JTzSAeMtCTVcN2gJEkCmZjTwA57JogtafL
g7D2jcavJb3bYEawPzd7QWKTUlQDOLU3P5rzEsgPzklDrbUhaw4s4cfQz4TSY0J2
1yfmEL2X01tHFaDPAytwg4f5CPopgFxvYH2BLJXM8CgOqYC1gtBJJ0HrZUgcNrNi
FEHJEM5x/XrKcP3MaL89bEctN85VDmFCu1YY0Z42xazEJ+1cR0r0ZTp6gm5wIyS+
nu8oW+Ee+7vY5ju5EXgGrX1PU1llYLGrog5S5uCNLajbgnNLsRAnQ79S/Jq9HYaX
w6DgU2lpLFgeDmhFKJwrQbjtFv2yNr8EbRckqxFQIPo/YokmLNm3veuPipZpFPyL
kpgpKbVld1Mr3NqnP1sBcd/7neC4Z92RpVobxYvRGROLTg7Yj74U+bJFAGdtMw1j
rkdEsJDE2hYhOBb740/y0ga4+N76wzjWyZ5BWE50/K9RhA31UV/0vIAXK3vB+8w6
g3q5XlCLSTVBBSZrWtDkLzToZ8duXQn9VIISULsLMI+pURC6B8HI99uFyNxM01SK
EJMQT/lzzvCB1YQsZ99vsGxaA2yfeUN1xxYqw8WqewjEfr/8nLEUfDvpKyEsBgNA
GAgjF8W16+2tQluNPX6EIn8hNrQMYuUElolHJqVRjvdVTmIa1FqPfUHO2scj9LO8
gnZCrlebqLgI2RLV1fYeRGALq0JvPrtFIQaLXjj1E9xVepqQfrcGcG6URzEFm0jT
ju8Vji3U9+IL1MfdoVHJI6A+lvKPQyIXPyeqgBzEFxHk8ksz1giLzfFPtibTqAoL
Wo4NZsbku4Fjkgf6xK+rxXYs7+u4K4MXU3m9etflGJn/nhtTjN1IV46JRjhi4IC+
q2MnuWfEIku3hsqIvd9JhMQmIJoFbKrkjkzIYzSqcRZWFFJsUVWX543I6x1eAy/q
cqXC07oGmgwtvz2SgUno9+nzrkiH7TKcZ4xaGPAbiqJVpx6mIHYJaTfUksbGFBrC
IPkRJPjrxlfIO+qa9TK+A6RsXkpo7KnOcixqWgwahXrdXqFfKF1z7DDBtu936sUC
jkn8PkVGN6NJmOmy+UNjRRvQzY4p8XtKfkYDENSfPuFnZ8ctBPjfEG+Rok8SSVhD
tRpyIRCJIbAaeflmL4+hL8lcHubf0CwrJOtXbY0pui++YCMWqhTbkK6YjtW/fcEq
BVQ+bd+FHoMsuA+KFXdnAnsiofvTmH+PS0fzZl/P/EuYvzoAJ9cBSbFL2X58wpHl
hyvkfmJyZJn6DFX6vneOvviSp8P4auPArfEUpRyxnrM5U8mOcbZ0CEu7GyGD2Oce
Zj0Ki1IAczgGJYrkbSZASmKMAdYPWxHUpZ1O6jM0HZwDg6kJv3Lme+wvROlWerkL
t4VVr7Vs72ccb0Qt2rnA2CoGUCk+rvA5kzcyaJED4M5efsL7tZVCZqRPvCE83Svi
az0cN19VmbbzMFZsyKwSx9YP946EyB3yn8i7cR2P6sEguJBpD16Jx0KFKEUABZYC
bWrJ/85HUlyVoNcmJgmG6GEQ0UdsJa/TIT91liqpNaowwTJPK9ajej+QbaVy6ztF
MIYhGFT/GHwLloN1eBWpDwQWpKL6xBPeWLdQMLPH01+Dsw/aWrs657POgh1JC3yZ
TijBO1w44TGh7QYBIYPez11ii9/k+j5eeScldi0i0vji8kXJpKXp3FMONoZHwUyJ
XHsBONOA9RqWuWbXIYYTKqvhSv9yuBfAKojUgAarVUSdSjxyZYxKraYBfsg7lsx/
k5HhPxwdIdz3erD8dSBiSLpvEGv+9G4vlXek8zc8O8+EFskNTJNpGd/jayfBq/oz
s6w0QkWBTpd042f5rsq/3XOoGe7Jdf8NevsxLrmp9HH1uL8+rANNQ/wj05fFRDqE
db0Z1vjZ3Bt+cOj2HfK/6QQSexsf/iBdjROW2l9xLaQ5r5b4REYKSla9MCXDwly4
iZTDXtp28VL7Z7AFAF4VUgTXRx1B86tat7pelrZMqEQM9CIB6YLM0r5aZib5XAWg
3oZk32qXvOTtODtgEcVF/+0XWOcGCORHs179STCAUt04Q2m44lnP8gEPKkv/qh7L
0IQyAknvLPICJLor0a29K7Cl5Bl2t6qSgyxpYd/gTfKluth7Z1a2U8e+hxGTcMOm
AgXqsgOla+Gk7ndpO++jiA/bIQ2/q+B59fmc9SbCC7f3YTxcgOKwcOTyo/OxbH7P
mRuGcaaUFsbABZs5unIf+rJUy3QhvooekZs2rrNX6Z+jLm3eob8JqfEmcOuTBpZl
WFYKS+X2AQ1rlh1A6FlF7fQV+d9pZJH+R3tpY7fhcpCJeSvWEd3kMrqeEjUZH6+Q
jK8qvlvexWfTU4tfTg5muBpZsanPz/5Ue/Qde+9ULA9ffmihQKGlVUD9loZ+PtXA
hY+cTACcJley7HhJ2LaSuSTV9QDTs56z86Fs/1TW/fiGNHC1i9wLDwykMDys6U7P
1nE9nPj4V7L+xvqbwNx5CjDcKL4lBqgi8kj+XPDrmVVRaq8xpZgiBvLm0qP4lwqX
ZPwlcTirs8Du8t6O1HkYQXZMhnjqzC4AkmwhBvoEdxq19ykkaybq5oIQqz3JZmPg
FBGG5txT5NAxxuWOzaIHyYNxveXsINfXozlpuRd3EtSWkCiVGBkKP1Vab7//8x/f
KxYGOlWfMH8AxZ9uVyTLVBK6j7/HZQEpwMVUxag7zRuJcCsoBQcYQmxTOBT5eGPv
5AM0G4WkLpvysVUSyFyf/pBRpHkDnUQKrGCs7hiaXmlCeRS5hWc7+0MDTq9ffp56
wuI4q9lXjLGOWfp/wuMwzOG8nnm2guBu+Z+2gXHCap7ME/a4RgItAc6qPRtV+9AA
4vlMuLui3BeE4QltR3/G6aCtt+Q5YV4Csx9mkAdTFs3fglyb8WwGoeKPpFTbK0vc
akOULKgeJSZzcZsZPlCH1YdY9WZx/IZE6mzxbt2hruItsUJajvFiquAVD21ZiUgb
1ED+O4H1t1gMUeqfpZ0ylVDyauBOsiTLg8KMRDhDvnIQuVdvlEzuHKhy8D1oPDFI
XmIelWGIvNRjT+0rw7AOgoUQIk/87yxfg4bK5/Ueep3TMDcgo6Y6iQp2AJaA8FQK
qxci/Hb/OZCReGIumeBoXpRg7gPxE9tfK6NhhRNsEdcBXVa/v7jrxDZ+lkJ3+FeN
CceyCEaVPI34uUvo04aURbUqU9IS3R/ZZdxMCsUz7Clmmjq2OaKAPTdDO3HsPPPM
3sjIZHkXx2Uf+J1XqhbK3ZNTr1P0syKwgkM53nsfPl+K4KaH4ZAQtZmzSDfkMWVC
kk7VWY2BivfyQaXFafoGjOLyxGZauOfKnSo2Sv3NN9nR2VCPzvEo62MGjo4IUnAU
M5gL+/vgWzXCRHEOO10kvZUJxH2xKe3VKwedvyF071QvVike4DouHajnkEPCdoHH
BX3o6wn4g4QbRPunqxe7egz7VwaViD25nC58Zpr4hFA2zXmD2vnsDkOmkDMF1Er5
xRrajNh/5cCpTP9dcdqMZLyjRAIUK8kKonN1HmqLPoxGqHMAdEHR4BkJSWdZ+A9C
/mQ6jY7CEB3mRBgbUkapyTWigDwC8cIfbRXXNfdjiqsykVAgVyWm3McwrMyy76JE
6WOmDEIyWeCQabbR2ufBILkTmzuqgPeFX3gv87/ZhcOqkXJyYM4gKo9FyC48vfCp
aesEGoA+SDV7tdvkUGZTI+1w8k15dfNhDUELY95eklrJq2jbG6obCEqVpjqbxqL2
cGFBVw+aD7q5qhGQVYi1+oD45Ueei7lyt4F1ThScwJTocUfy3tGSITDpSSRikZtD
e0TApJ+u1LNq9aTotUw/S8sIcI5/ue+WzR/i9kFBghSUXaj1gQXyvJahbBQmjDbQ
2wBH81rLDrW5nAtsKhm1nqau1SLQWqP4KYByrjp8J6vZqErlatlQYnUpjYVrLC/D
zmetXyEavk6+hEHkgw5kEjec5gjL6xOhskY/xgVNw2KDjHwi1S6uM524BJvUItdy
JpXSO9gid3dyeDgN/KFM0ynYDMonydpXbVt60KrWFzxvHfdcnY074RzMGHbqn5Ae
MXQ6w6i2t5BKlER53hGkT/ksbJXneBHf5m00SrSuyK5sUBvllWX7/lfuDjjwBo2t
PCwZtbFxX5VbRSPTW5FrE3r+X1kegsWUxDzASnofnTnKv1aJrP6l77bHXC+JiEYP
drlRHxKrC1VrSQip4W5WdS/kJuw6jRBEh6up9o8JfXVL6IkNNtFvxi4z8h67UYsY
MRjTwdQp90Ea+t08jPpplXw8ubw3o1BqJi86ndfNPJwgeVfeLcODGMVjSktBqKFl
snbdCyLJswNEe6uDqKyJ6vYbh1AR+miJ3OBq6nhc1X6RPuzTnox8O8xJKPEfyCNp
O68qC3pfnXYCM3n2fGFNlkowX5E96jwTZzaGj1In0vh1Ix5wK5JOEabxoeSlKVNl
8gulcbI7xlf9Dh2JzuYz6Xe4PLsrSNmmZ12P5J73JJePlT7wVRqJLiZpu9CxWjcI
PjUzhmUR980ejNS44egFI5k+zTgtWK7sBn2F4cUdiyX2wuu71etzSdOlqyAF9e+A
CeL4+I38cyP8g6NT6uxXmqltro5zHS6EHLZzrukdlO6iEZ/wWjied34VAY/0eKpT
vQghfBQyO6qE5RPX0/ywPc22YgupT0vStnIYVdV35A/1kXxWg5M2z2zKmPL0E7gJ
8WQXJW+p+KJDkr1uxU7yKjBtmnxS9ErLLTV59AR2i98pLzzPF8Wb+ZKM9Pob5waI
4AScRzGdN/uiiMOvN8KZQ+q2f/K7aiL7Fe3qIkMM8WiDHhB4yxsMuhP7nR05ILFi
x6PPiPtBOa5Zri6qX9Au7kofgE5Zl0BQL/XgGBTyGpVCnhl/1mYAPzGSdEhbJsbc
RAtA1WTG2Xvv69bL/k1K1zWW0zHCiBnws1UihXBl3HHrKTiZwezL6EeM1ZkuvuGX
ozpY1NW92uYX7oJy/r+Zdzk4oWHM2YDrDQ1NOjPFTRlHRBOL/uxCMXrwfxaL+bQ7
ueMruHJ6/DR0HBxwKyDHouRDGNzB0+hES0To9SXRo7LdxwKPYomQTdLRi/ifIKzR
AMg+ngowYuIILut2CkE1abKE1qih6osatdVN2ES+XshMTICGVclHauig3vc2+wwF
whIg+AFEPY1/WNlHq1hbQ/m1rybSQZveLxxVGfSD7zDzRQwo5OXPfLr0fwnN5I7t
3radrwy7mfxZkclBpq5Otxuv/ePudyOFOubW395MF+rya2FAdRmj7jJtHpQqcE7X
3SNOcyF+nxwPfKQmTCPDFQfUqrnEoWwwLyxxyl/kcwidqUubOAfGciOD1HkSBqNa
Mj9EbQ0wnwNLyw4bVLB6xbIiIOOz5KF/MtEIU8/M/JegjYWKEIH7XVTzEZTDbLH1
bKsIdI9I6wBxLOts3VrtJIS2Uzk/USylTc7+aY5Lk8hNs6S15FkX+342pR+Lc16T
LeU0BQIGbjl0/n/admrpnZRntZyEVRNv08BK64bvRg4peAUz5zE1GILl0v6cV6Oj
FFTTassmhqHRbu8SL5w66bBkHCyLbIh9hwGxFR0Zf3IqhYlbkyU/ckwYQqRNZ/Rn
BBvS7L0KBFif8VH6Ww02U/YKe7J5ryd2IycFcwiBhwIlsTgwXI7AZS63bB1YgN4a
E0oqMI20Qg3U3uea+zIPbV02K2loIyJchj56JlFNdOjoRRJ+oUmzvIbdB9Px3Kwx
a+QypIEyP1rqgMFERWx/8Q73PcxDipc1CxgJEQvbEgCuOiYyZ66s3DCGNWsc9xOm
0amvy01nTOReqCYl6m1J3WplOgJNfxORR3O+mEMPEbTsSaK+xFzBGIO43bD1jtLx
zSj3WxVmCk4+2xbOrDO7eKdAGFeS6jgZCttQ1KFrxmGQx1s9ROBozmPtm4igjxsk
W7SJDFVsAeHUQp9uKyXDNu2Y/AhbibZX09o0Y2h7pv4rMabfMqwym008rUYdy1UF
ezN31SeGJHmmXAzDKxcjz+N4FlYmZHfEn8FuyjC7Gcj06HFX6HDQZap21ocm5Q5r
scOZzRuWr4o5KCymE9odK0Cc7RYMNhkhQ8f0/RaCZdTRNXrpblL49AfJue3rtq47
uptSO3rechq2h/eABZYKz9IMGk8U40HYkLHE0DUq89QkjZXVqBwwxWhObb7nPe2t
8ldpZSyXSHQqI36PE9lH92tgJt7t6lfFw7+qSP5q0sBwuLNiwj7VoTo0e4jajeqC
PR2MZeZ0+RShqXz7BEFj7vHjs2OuyO0W/thWtPr67X11ebb1fU1zqoY91xy70AXs
9Odmw/hhCHceUF5hK5LiP8AJRZq/gg7O+crDw79fCUds4Z2CDVE6eHlDNaV1fIsS
bz/n9PGiH4Js6Vi9NSpNmQCRt/cdq2Uci/vkIcyOUqWqovZvRwxbDG1No1qsnYaL
scf2GLQ/ybblDOSAA8PezwydrBwEmxjS6/bfqeicju7dSWRdx6Xd+7a31W/488dm
oYiuXjH3ykhp8GC2tU1Pjm6oB0lG48uhKWX4/QKnpfD+Na7dbBqTD3tvD8IZkFfK
MS6OZJ5HfjeafvPq6eGAXm4Zqial9mquqEoqPzcw6uuT+Mv57tvdCTtR5CCHqi9e
dZ6G1dLX+5vnlyVdQlYrGNYkUJklYGpxfrJsqwaMpCavMkiQXr7627m/8AyV8YBP
U/zy/HPu8FrLRjMFAhfScHNYm0qm/F1gi7rA2vPaSWB7ArMzzEvAzM+A8XNkUGEf
ICrw/Mfc0LACWr2mrwRmvx9lVJVvdMT7ZXWafnvsYtawF5MXVhFOfZbxLm5Miu2X
WRXyXRE+FDcR+pYkGXCdYsmKtQTqIKk3wWDU1B+LgT/SdOrXzMpufh6BZgnV6SNl
eThRzoWvNKdFBg2be6T1LxelZ/Z2bQGp/bU836Lx0gWOD47QBMtfqTw1wfESlATj
fpIgH5YprS7Wo0/G6CPmnHwTgFYK1qe5oYyrRIzI2iog9hv+ICnglMwxQXQ5KR11
y4g6B2kXDXjMafU7UWWLO0Z8Mp/XgU8mlHIqO3HK2fbAYXgM+bv9S45Vg8aaEeCT
tDdqnHDIh9DGMXQsE/qnIWl1CBTiiYfgU6k1yrJX5Vxmdf4VRtHUMl7R408NDksh
RshVDF2yvMtfvRHsVBmv0FQSMD4u0TAnFS4yhAJ9vBEcnAqdNcsipOE1J1zD07pl
/9dypbr4G5/kiZUFYghKntQWzGZ7TYDiFPjY4jDI11x3p/sdoZ8ZbnzlEQuCnbFM
6hkb/mBiQFq4AL9t98oqjHoBVeieeYiemKeV0PP9oHvoms9UsMuHOVqRmDDb1yrP
9/dnAV6xMaxmYOvdvPnC61dYUFYI/tgyDgbT11EaWWNPMSBqVyy9+BnC3avR0t/J
fc3qDXNU9CSrqdNnLR/0WRiv2RRvUMinGtN5LCR/N0guJp3xLY9XljXJq4rG5ZsI
eiL5LtMApItyXugTEcG9uz9qFwo5VRGpEeMNLxMt3nmavxHK/2VgBd0jDD+/4Xoj
eOmEuWKVth7pArlUxFhBTQcyVGsZFVYxpmulx7Ps4ILGG7yiDPySTs1u44xmb8uj
poyJK48AKoXQqTY3Y9W59C5rKOy2B8X9oeBe51sLqj6S/69VS/8ihG1sNANxVFpX
cYA5H9c4wBNgHEXRrn+ZbsGChrXjdSmNRbn5UJVuz+EUm2Ugwy8JvWgH/wLc+hMZ
VhohoepIKFVMbVpy+IRuQfslOyJ1XT6jHEtwQUH6PDq/K4PJyOD7bYvKTc4VcTTB
V38m8T+oC/fTJj9PZ8utFmmKsBBILmIqXMapHNhU5PfuN5Pe5OtXAl+9bRFYGLQD
Jj/nkedBxI7OzK/bMNzw4zvGt5+l9329qsWHY5dd+pL5lK/H0p2pcEFZGPXkC/H8
9OioRH5Mi4K3ZcXRZGKemHPHHVM23DRW/S4YfGRJeJv985juzvfKB9QKA04LirXw
tOTgutLKhgWSqXyDIY4BFZVSbQKRhXxN1DarFEI1SkAMimDsuDSCcuKAFpJUOpYQ
8szvoKLmVcPLezjAmONKBJ9UaYoJTpUws6AlECKLJnA823pYOjFEmMM9lnpGK0+o
GSxV0Ay0owTXOl1aDe5Aham3JmglF8K2moJ9N2DugxsCKNHDwo9V/GuEIPHEMQlb
eqSLy9102tc5HBOCknqLcMioriDQAetT15GDZ0u8q8o2bNSARj18qeJD2s68/1mI
gLcQrdSbhv6w9xYDarQBzQWiaVc0fhhnaDQl+c+A4VTr+cT+tK+4IllOCkz/Fquo
l+yxblfFGCIQYpetzRoCdXg2rVQcWTpVpbk+qsjPPwiZ8o8kRVt6kzL2gn7XzNZy
FxhfqTi6zV1oq4EHZRrgzBaFCTPu0MyyZD/ey296gVZ6NuQugP+j0dfnT1S+C+ke
IKQOg23TDy25VCIBXzkSgNWL0DPiMiymoX8yiatsqp92fge9ILCkdwU4jRwlDTTu
hTvllisfUFzSShmeotF8+eeSSyo0V7K6fsNxKA7PHNQvifBjqVK9KxnxE6ftCMLv
R2Br8n1//nHLy6+tlJCYmAqORQuXExC8caQRPJx9Ei4tDLNZbwr8NoPaeyscIkPr
XHmMv8hJjfW+s0Q812dJDPKYlWR1vQCOG8CcXSbmKOBiRet0+GFUeizkS8oQL8Tt
RhuoaoRCMvV51+y1fkj0JT3VVhIvZEzRJBuzaBbCht4CxEbWSKLLMt4o384t40tP
5ZqntS0JBVAwowUU3o5w8UdCQd3MyL4596woelhF+W5rKGPZyGw22Mlfc6VJPvi4
qTNAb3fD82XuAdGHNAYslelSscMqwzUOr5XKvUNkQZbf39z6Gavdj4SU8vOfiQkv
fxdfDIA9S0WQFLi0GD+Uv7dptvCwDjKDl/8LTXX5vfDXbOYuA0rQOgQTxRHwOWRK
8apOazKoiGXgvGof74WdRKSkXzpm8FKnu1R8L50jKEfEfNh7FFhqrx8k3tRXZeVZ
0VYTwKv1lG36v7QF0pcNKu/MMl5XWRdayatwQVxfK44QlORF1gxoseHRlDtoZaq9
30HGbsaTMBqppKMHs24WJ+tEwU/wLX9TjaZSTDLeZz8inPrz+BCxh2EF7roRa1p3
m5YJPQKAA2CekkYZmqhfgBsHTJ1sl5aMVdmaLSZM7D6BX1ch0EpKbUpE1mNo1hXb
e77UVA6wf/sJE36HP4OWB6WCsuVYTNdi4kMp+ER9hAc+iDMsQhvOm5IZvCT6FR8f
UKyCJORTSvNgNxyGV02c4nDjRoSHOKIltMKHZYFtReG31K04bQl20+wlV9c6S929
Ai+XJxI3C8XE5v2tI5fUxySa9zL4FOVv2bNIy/O4Tk2E1yPidKptjmqiZ6wnievY
LPVR/tYQCoGWR6Fg/T8cgXmFo2vR/FP9ZmdQynf1zqxukXv7SOFME2haRU64ze/W
fWxoOIAfg6RFpXMMAf9imYQ4XjgEdJ7CPHszsgnY7ScKW2tMZHpMw8kC4U9E9IGn
I2m12Cb/xqgbV26KTqor0Y3NJWEQmYdTKc0QmRopdfFw9qON73mhlmnPGFG/jOcp
IuPWrLHvjli2snEK3jYXmhDbrk0pDKJRvSO+gQuqHFOi4ph/KXmbk0gHYCQWreAj
gHus2pCvFK3mwLzFBJiNcd+sw6p5VGAp72n7Buyr0EQ5Hm/0IFKg61djNx5In3vE
ffqu+tYd1eTcYXj2sArwbwZUgZ42EvYqQqRfdlW7g3baQU2SEEo7QrSoPIlaRswR
vK9QcL9gt+ZjT4ElxHJZSvXhv8/G7pCSYhaUr+4iW/1XDfXqz4NV2IZVZM7N5rpY
eG3/ECSb45b2RuZ8ryljPlZV9R7cVnwWo15gPLs8+NAFBjckyJyWqa36ZwPquEnj
HnIAmlyXpzqVaeWxjw/zP1N+3HdgIJr/AZO9epgMa9jP3Wvvaj/S8rSOf3r4dCLu
QVX10DkgPfviQpG7tyEawcjv7x5S0EK0TVqkwJdGJSuI+yJ6TKRuWuvgLjD7srfU
ak6CGEL/fSboqYw8mgN2ksrRVOkmQF7Avlmbi//vWAPdyvBPN6ea8n1IurxjhDSk
d/Y84en8w3gu3sELcfiZOMh6M7fIY0igOjuA7DGl2o4O8kOrskBA+gjvCJJ7GXeO
OvB4KTwExFoB5pck1Qa9go08NU5XO553WecW8jRNfI+0Y5Ngf5wu9gWlcLgycm8U
JSx/hlR2/SuQcmktEi6le4LjsYGdcHf55JHwDO5uh9j9U8lVgJBvRUb9F9ZOnyws
M5FYH0PwRsyldV2s3I+ZJoHRJqrZkh0YZBaSWXws4w36kgp2tZDE1p3TLYSqr59X
NB/1L5X3RM0y6VhlQRpfOl1roMgiMdG2cGoW8VdaZDHsjBy9JfIBjBZXkIW0yMBE
+ZnKhYzIaAXW10J8JEeDaAU1hZxnNiKEpeHeX5uhldqt8DzThqQQtfckbypTdB4s
47eDnZEgHv99I1LQ4NtLehy31cvJvt7JAwxNLw5hcCVVwS0W3jnMlGoogszMhjzK
zW050UUfZlTLdu11ySM6kB44nRTonxd+SvSAOZst5Kzxfos8mePCCoMhLavsfN0U
m5D23Yv9Ad17ZTV8RzrXKeZHN3fmmTmDFsU3SVELmrr4MI5WKQyQKp0gmLZV9GnQ
G9R4YHZi4Yj3wk3tGLmKmyxX3wDhAqWz+PONs3+It2izb6FiMUd+QKFNmdsgjPiG
dvRfSP6SPfsnqfwNqjhFo6Pgm2ukDMH9nH2VknRmBhhaNcNPXi6HicDBYKA3nfo5
PUiJcJpvxQJD8faf8ThRXbo5flWHICN73q3vq9ktwnwUoPDWXsQ3HwKQrcbugyDG
Q2+fLqU8DVBp88Dkr5yabu09YxPbtf+yQHcV/NxZgQeS3UqA/st1WfOP3VKZXuVk
OSAQ+Z69p7DrCOu7KiwbFgOO0FxAaegO1zV0A1juwtEUmOkeFMy4a7d9g+7/93uw
CQEo3DHdyECvUkJnBrWx9LrcndqWuukQOT5VTsiW3vW5THCado4Y9mQ1K2fP8K1c
ftTvVE1EsvyR4fW6mnyzCEa8mLgNLgXDb3LWO1fFbTLVUu3muHXFvS4AAqm2vYRu
CK04Rbb9R5wValN6KguSVfqfawtWk6mgSjj61XJJBV7mu9FzoHSW1rWzhaCfzZpE
XhyBr6puCcyC04pmqnZl5DCTk1YjfUHdyIb8cDqNXD0oKrhfjK+J/VX4Sat5rJqb
jL1bpwGP/hpxtEX1xH0XZhDzOiTHc3XyEQjjfy80miqKI1jUSLrLYG3ADa3yq2Hq
9/GqMUeGWZCX3HCwVHSqPSo5OyqTlOYiANbvwOXIx85BqaSIzLn4BGdBgr2OLlr2
1h17LHK1OyaCeS0y7kZZ98dgx58lmsPBCa81KePOGYiAgrwPgLoH1Zscd3Fch7P2
mOW0a+Io85MCX0kiUSFODciyVNfxVEckoL3ymwJTeg8yzgwoHRoCOsMXjGLhQlKu
Svji9arZikxCvDb4j0HDjmp7ysAVf4L74R6yVdP0M2gw7dQT7W9GGkhWhnhvDvqB
nztfdorOos7RFVu9nLcQXphAuVcGLfMIayMrjAZCWq/2ZAJYmJobzZ/oy7/1Peh+
JCJun6O3xlpzC7bXa6qr21cEwW44QzlC0BNErGlMGdNDm2qMYbD2eg1Gw8J6nPLS
DTzdly9TdKt7ruifaDQgg7HsOWKGTjKnGhyKaaMtub0uyctv7nzbGcnt2wHwZxVv
xlDgHbyhBS4F8v2NFpcBRHr13M0+a16lFb0sNOrzPnwY4tJNP3tn3BDn+u+EcB9N
ym7yW5Q3MWekZJ55zgXkwgwfMe6ZsDXvUoxoClCbe5FketVOhnUgfL1yGPa1I2Li
lrrrj/9X/d2FlAprGXc45FHiqJiWl9eC2567KE8BG3aTgY62vKHDafRkRYDZKD3m
QLroLAoHKrxYoEkUnfg7UjpVfWPG0TCjlAZHO3d6Kx0sukLtiNI4ud0lxA+fx56M
rUhIAxjwHcXQ9CQlUhiI4LGL8pd8hsXxWSvyO0L4Sf4/FJqhC2o7t0LkB+Cxv765
g2JkraEegT+WP+5k0VUHTfzROr19FDQDw8LotvR78pUYdPi/mf96H5v6Zzxu4Q67
8g1p4UXkQXFyVsK18Fx+weGwNMSLD/NXRHRbyKoDF9p2OD6nM8vZJZJ6bmBsgPCA
wiF/FV52B1O7ZdFZ4PfrdT15eMEF/95JPYxw9TB3CpGr36MehEbCYBe/MrPIrmy1
IAvrS1hC1PNsV4DwSehcNkBcgcOLEnUFVy53aAWdYl7QK01eCryiUKQoM0YRUbLr
IdICn7kCKtFT0+yqfNn0zdN2zWs5PFHbQqAW0GnPkMs3ta0Pd/r8C5qC4yHJCcIp
pqpTqxVi8l45CKMeyK3e8cXroqyXnmZKBRLWKEVpEVmnRztu0Dth1QTU7Tn4Gung
y3ddGnGFogU6USXozJIPtSH9IS5a5YNeUiP5dfv7MlXjYGCiIqC0Ua2woqO3r2H5
GrEtmCYBzl9Td7w6AYy1zgaFlFcKXMlyL2bSu58Xv3Is03xUw7ByeKP/62I4RsTh
LfoNhN1Tugse6VOg+y0Bxfk9QYGV0V4N/S1iAIzMsEAxWuYWTlYZdIIESUWLgFkJ
5EjJXslcLZJGsH0pRk4NgsaYXBDywfzGnVZ8Fg8ipt28KSrJqGvCLSg8zdXnoZgx
vWo88JChMSq5NKYNwoVf5JI6Jcw1qvZrPgQL+VnAHy4RhpThvzXVrWNxENnHduzD
4YQ3srv69poUICMV4fmaj3x9vFI5yIQgcX7v55u1fKXBqxYBergPf2ChAbbhVIrE
Pcat2ukVjQX4g2nxD73EIonSEMb7AkRe8L0ZTUPz3D0HBoUb8N82HkjAGbYCT0DZ
hJjY7Cj318lJVqvtuJ2xJcYexLi75IbUiETd9vOGVic9f0MBgTBlVVOmhR3qcek3
B1rg2DR/inosVt1ie9/m5rRZ+B4l0VIhZMAyMirVwKcN6EYeeJZyzpmGzJiY2Ij7
E9MYSSeRg8JJqAS98OcbuDoERTljPNhL89aUA96GfmiuSRSvtu1coGpPhb1feEA1
Iesk6UxupHMzfg+SmTN7a5MfCmjJOLu4AMltKnV7qnaxUkyRCkqedpqbFscoqxub
LYj9xzZRS1Wqcn12OfXtmTXMGR44aHgB8v5rGeoLrZdLyE2u193j+/OpNLo/8GOR
K27E8SqPCBkDzcJaBWaslXL5ivcyFgCyHc8bL0cUc7NSk1coq3ahqgcUhDjlJT2m
tWztfjIQQzqLwj8QRUXgtgMAydFUCD/04mf4t+DgygzTSOfqS2WLSDTOlPU2zpaw
SjwfVKOki6wCCRagbUG4jdOwvhS1xo26R6ZUXWk1dxehZTGx04m5LC0l/m0Zdczr
C5pOtS4hAJ51phpqfgOyTKSjW5Sk058jROd8PYxFmAIAtjBRrTTAIX5MLzeMV04W
f1rm8KhqASkiIPvLhz0AP+KWTQHf2Gm6NqdQzsJxl3RaQ930C58rv1VZ20rHDZzw
qUL8ZAq1DJuWbnxSyea1LpyjvcEvmafH6jnpp+hgBKMwoLet7q3c+JsOXhgs0QV/
KsSwynzhTS+dVRrf7h67JKrhe86YESxVY2ZQIt1eIlPLBitlkx9sPjsTutLz2Okn
ipQzWzOptUN+fQekqw/M2aV44Lcf8/X82XCaDuGHV3AR85lWdsKnI8hiE1YeDvvo
v+uDHb8xIgp/QuWN8guoxrTWQKrs+SiosXSeNms3VF4pAuoK9roHVrGvtXeXLvBt
Z2qYpPFzPiX1gkbrI1sk3FkWypGBEKKdJF6e7yY73YyZ4zXwU4byFDvU13BJcmED
fzaGOkW4dzq27lZwnEGY/E1P3GDHlm23s1YyUppejpda+7cNZ248kIG7tv/YwPcN
ctwWddeyVRqvm7WxuT/FvfS6DzXcYQnf5TZXuth34SfER+jIHkEzq4q5bw4ySEnK
ZQ3VZR6P2MMGVIYdNgl4vwbE83WgzlC5MBGycQIwsPhOTWN4QOHN2ENZrun2Pcy0
p9xJjy0ffr2gYliBOodkQq6poZL9/zs49kVcPI9/Lx/mk3Fmvq80fn77DboY+cEf
/cEGjeuqXEtW1VrJTYfy7NdICOydQnsCaFJO1Ps2/X8iUw2WjeIgYccjhWk7hSKT
8nkc1o0V9N9yG7BRUK/ysnOaZpn/ewAecc/OG6kdVZahjNc+EfBjfred5DIGQZow
tecQ+jItPpYM/ynK9Ix2HKbgrpOvSk/ey+A5DCHVUvufX0HL5JXGO3ecOeXqySvU
k8tEd9kIUbft5hBCDpqOx8W+qzI6B4Up3+nJzM3rcYQ+dSYOXwcz6Jp7Je4vjUh4
ldooNqMTffikiI1GkUwKrPVRHR7Rqn0H7ALmOhu1Y7Y1BPrRArOZTLYqjFU1GDh8
zt5a6qGaN0MReog+rBdk9zF3dfWQno3htrKa0HfeXaXWDXrB4b+0ewoEMH0DbGsS
iGSraZpfiiaeItznHqB6s8w6YUEVweLwOcAHP+5GVCRKhU0vyGopp0zhm9CXh+CD
Zm4J2U92bkeWFUIKeHe5ojmVHE9+h+Qj8s82zfwinqwLwX30EMGvina3k3a3EzTr
md2P7bPCd0eZchlqxlCAI0xzdFZnNMvYe9fHFHU39zGBoIF8MXJ1PZsw+cyPHKHj
MwQ4H6H0OQ5vW3Slkphqw4yQxWBuk7PiPyn71D3ltlbBFQUPmHKtufQ6CWfPSaO3
hTFiAdLOnhWAMzUwtssMhfCkANR9RYQwimeKzilk1aUTVEAbLgHidC+fNfqsOZtN
7zyenWxBHkDNq2rDviBO1e7iuvMvkJhxcCpwfgt58E5jueBJWq7NceK7wFgJKDJ4
SEIExOkUatAXpKgB/snBCWcrzHIJWMAmzXYZAk8BCp/deckDCRP+7l7dXlMS79UL
Fd5p+jexcELNpEALiWjZmFLauwHggjORBGWuQY/zj4cRDxApiXwIfaZY5VItNEhY
xHUnY7HOpvJ7kH8RwADQ7OqdBJV63szpvGIjAVQYKzeVi9SJ+8Sw9K7nO0bpyg0O
E5zOtAEgrTy5QpNL5WWsOgpCXRD7vKUBeWHtakMBFoh7MGz1pBQfVDelCskNoWMM
ZeZsg5iBjpYWVVMmOjo0rC8VYHOBCH+MwNT/SwEvphjlVACKxUD7QiMiJdaUcVam
KQ7W4Y/EtLwsPHLmZH1CRguQkKWX3wVSI8It65cH3WzkebU83XUWN2Jp7MtoO7I1
06roYg0zgqNKLBz0CLWLp4pUAAzQ4qqNh4OMdmjUyt+14PmMzSli41mP2CbIHOBZ
NogfFLeYi12LXqoH0L+T/CqlDQ84ynSL2N75s9zEu2xgg4LSlr3+ZhHSXfxgh8HZ
/WdrMZqc9nTL3wNe7Z5fgBL1e6SaT6oRCx0DuXWEKm3H79GDwVu8jZLZ3ldrrcpk
KDy4cwpuRuGh4aXZIsIk1uMIJjjokmJgh4kdKInlEV+t4g0pbzIUXEuy/0gZlwhG
QvKE7Be9PBRr06k41ocRsIVxtdSwG0wxwCgEQyA0GF0SEqFa5hcCZitcTq5EKer1
jiT0lYmhH/xGlaRDKbmHctwjPoBuWiM5rP+qI+l72ZTWA8ijHzzKMJnd6Dd8shoT
fWS4cz5I9b1C7WkSNjOzMdjagzuU2dvY+7oJ/ja8Pk/HCCijjEo2hZRe0at8wlc1
DA8dfb37T/3A1bO4peuZ1nAVeO37AbKLR2M5Tzf4By7c96/rEOaCaxVnk4wVObvr
GXVZ2y7yqYK1oyTVtpF9saWyL6gmxko3JS84A+qgAF0vfcisSh5QC/wt22DxYUr9
s9uw6TWsocGPD4aEGffY8dYPCNgQpIj+4Z8K8cc+wgdXYaHLdmJjRpbnwoZYEsDj
DHt+vs/XqnIJ+LYXjD5n7SQZALyTDLmJKE5pvJewNNVz1Sfu6Bl2itBzUEiGHbCG
fkPUGzpS2WTXsNM+I5p2Lc4PVBplRf4iadSntiiQCJdp/tqFGf9IWLbw6jT27Bg3
B6+xXIx1+jQ3ZITpUgCW4nnpoeIsARXCa9cqo2wyNxynKjEVCN4I+cTreuNkOtPJ
8HWutLLkTvEfCFxOLZ7vX2u9i+uZGxrEUNb0G2YBUw3Fel+n5lIidLrgsCDTwklS
ywWG2I64NaQysfidcaXtSszDRKbTLzjVOdh5drNTD5J8J5BpKvXEEPSV74GXcQhd
z78nygqtama68xr5vA+jJpUzl98lYPpA7guWx25wGNUW7Wnwty0vAlsI936lBFot
P9DlLIYHJBUR5+12UjRRmlYUzRAi5DSBHH0w2LDr0cWhl6mjYXz1mMWDY3SYXeWw
yJvM80hzwBcgoPhBuzWpuhu5X3TGxOsFL9NOhuUwcDnKSLpAF4rMewAarI6P+lbI
A9SQbUHjhvHQ/n7JFEXOJj42uAVPFAIetpGZQ69z9FX3NbB7S0nD3ra58e71MGO5
IFdLY22v1V47EF5TuI+/PhzUdEnoTs0j3tofKtopQrwNivk/TaQKVrmiVp6smp/R
V3U7GniSpR1sXecQVrkAwiCJWtPK9YSmUh1MlxtP6pA3Jawo+VUg9oVNY0l0gOnZ
8RdctGlnopi1oJ7vwM9b2M98pOIka9f8NR+Yrq+E1JSttMuK8JELw4TGJP7kpoWw
gdtDP4SO+0S35dQjE+WgaG9THWppaj0Ip4cnRorVw/jp8rzNtOprsho5Oxu8yHgS
FkufHjr0ZbyugGu0l5mSKC8juBhAArOSwRCu8LbYJcqH+152CZCEzwHtVX7j0RDx
KlTBuYFDmAibBNWAxMBH1WyRX+Cr10jsjoZ1m8r+dpw3udDZaGk6C+w15mvJL4tz
mJ41QrhBhQc1fVA4GQht/zUmCUl0VFxBLVetdtw8FPVHaFlJGN3oEXXwsyZvHSUf
VQKO/FSeaRkLWwdYRU8fb2g9C0EeP+w9gtJKUWdxkJ/0G5tYNBYwCvS8eZwlLiKf
eIZ8dmbMhhAAlc9eqWztDNk5ECj5T/W8tsl4sYzimZX6dLUj+HbMEoUOXpItR8kt
nK/C91PN0DP3nB1PXB3JL62V7XBnMdjiXlioNbUhr+MggHd4nKoCWPjCdxUSiZBG
C6EvrQxvZ0Our6EnSvUgilfEvcrWlnOWONejus5wqexn/Ev9/9krnjRW5v3+NdC+
b2T/kiZSJC6bVhcCnbVElQzjTP399+C5OJ9hRPpphRUknahCs8ZRBnWHrdLRuNn5
9PVMqXX0BtvgP43DTqKcpekgNR+ckyMnYvfpTkXxyVF/vMj2MzHC8Sbvku8iD3Eh
+8r5Sdqfdm+9wInhUzw090a9wEbE4eo34QwnkiqMNd/yfFIURXGR+2ixMQ+YNtfp
WI0UqGBKEP+yuicqJLcNAXikyYYM2RK1L+h03aJ2RXRqfoVdwlMuwvR60m5Nj33H
SuFzEeVtek1BFL2qRGaBhiRSwZFVjGie5K0jwnl/bACzvyY9W/2PxERft6lT7JUi
0Cwz5qIxpI98y/5Pn7S+OzVN87tnULdckg/J+rK1r4+lh5m27EU6L7v8+bFoKShI
aDyJeEU1zZncFv1YJ+1tKW7jfYZsYHN7DvdTuYC0+LKyOfOYNcu/SI1BeEmV6jDZ
I/fj1htf3XaQu1qg/S5K1w//OGZ5UzWV2i3VBAKvkYmDVhOSk0qRAZHIiff3QpJv
I/lFteMB28zdo5G6lPkID0p5szgY6SG+ix1yVIBVegiq8NfPoCV6Z8RCyTyZyxC9
/h3NgqSfgADMrSwcRZ5ZMH5C+LmUUt/1IAtKrETWM712SDRvnp0TWGFipi86g3RN
wylRTqCMg+v2Zm22JmoG9D2C3h0S0vUNwy/F3A50kcvl9NGEwiE4UkndMfElQhKI
CYv1ppXfeBTZBgwXg/pveYrDL5GCb5+BWGzT7b5ZC43nLGIUxma4N6+yDeArcGza
SvJaGT4o7zq2NHaZK7N+wfT1NYAR+cfM6S4VA09ZRb35+nkU0MtqFUntAJFetfKR
hrY/osv5t4e6FVlZwOA4Rn5UE8dkqSypRVpls9C+QhUTdo6iLX6/xT84ofj6Ll84
BtunYQhuJleOKENtXImDny8+iqu7plFg02pKbLmv2glcJewtANBkT/fboo7Hv9Oo
J1UnNVIK/sLQukPsrqXyVamGQKJyQRNMXeOhnxh0+aK+CzcJI6AGeenh8iolF51x
B4p2cC6QwcppqcPvaNee/N8MCoquWYXhYuMkPWJULRib7c3/JXf+g+1MIg9ClHze
ld0KJgu338+x7eXaGTER7X1MMrusPYpOMBCfLYBsWQYeY/XNrmGdJWY1BnN/qCbC
9DhgKkCRGrpuV+DvbtT6xNGu0WOyKb88F8NiU6z4T9yGxGMFqwbYHUiySCm605/A
onFcKaf2yLBlheHmyWObtFY4hESUWA2VhMJSfy+fy2LtbkhOL9JbNhkkA6+Baa0O
MpPjFulbTVkN8hbRRximfFptyJZX99ReZNMUJ71xaTfKA2DkoOwYJdZqUG/hL5Ff
nuMQ15Vhj3tnteEdd+0J/ECEaZCkWrd9rsLtpMcFMDMLyBzbdjYh5NHL1XK4p2AX
9CrPIJYeviEAjELD+AdswmQghyRDc2/CvPrbbX3CNTKSWGcQdfjj3iBhhYk70CCy
Xzj9sSq7Y77kKYW46mn6LfrzIRDvLBKGtjCUosXu3qOIybrKe6GlsPqbJAbtJ8hm
lZLjLLnJW8SZsS/C0C5GhXnx0LimFnKlj2B7x5ul3jyRLB+wQlLUaJ85pmZX2sCJ
iNYbWfojVcB7inLpimc7Gxz80IpEtkT7wFExuZ4KKhyTewDkkImLap3rdGCqBbts
32ZHchmEdBAbNwj8gM7xbot2eBaAx0ZFHdvC8FG42+2TPyQ185lAR5H+UhEoVyuf
kMzokVm0gQOl2Qk7utpBhWhnNaY97xX6tGEsVYXJDdal+RTkRmUwX5+LKvm3op9+
aX5FtxyrXTOb06BhD2ErBcR3wmgS3eZBxryJaL+kb6Va0W0XuEfPImCutPXym1sg
Ue7lrwWDcLP2wFqxfW9H9wzuQq8X2VU6kSinhBa69tGQJbKNA0QAXYeZhnNFcdKV
Bvigi2s6jld5o/D+8XnAzZwajRaR9/+fhqEj2wdnAO2aU4bxKnFO6kucVW3mcRTx
cuoXAJ6gq+uR11oVbVM6R6lKYohomGbX7UaoCH3nPwwZJWK4GJBqeP1VRLMKi45d
LtZIYV+o2yLgEdv2ZZHn2KC5zhQ/5rdTKnS4r5RpRB21s04ijRsOiK4GlV4RB4M6
v/dBj1fZbldEcYmXqoJMG7SxgTezjAb2WLfvFfLexS+W0S+Pja4z6frEyu0ZXHGC
t4ptkzqFSHTJnIl8F6tx8I2PuRL+4oel6mCjD5/sV+EsYwpWQ7KqZIIvqI+0eJuQ
8kiLwMIcPXcSTPcYTVKaQ24H5exqH2QQ1Cp4RiRRHCDd72UMqYMzySUszHA3g3BT
Et8gzoIA4ViOhEsaQHb+mIfwtj6P/w/xqsivc+ktcdq6xe47VqCOahgAPaDAN/jK
4OFx5aCS5eDgILe4EQfd0IJKTJwP16uZYWnlbf/VqKyFk++8Yz8oamiN6NeR2wXP
Uyt1XnZgSiRedsFXGmF0ewzl05+Y/Ab4Q9wEhgaEyATfYisDjFyXWxjrnUBwaTFj
wQVwdJacCs/j/W+lDCedxhX2J7xulsw6C5gqa5XFico/XAFrWw1E4bVU+cq/Zjgi
dRrJYQvFMULI1aPdRt45Lq90Qhc65VjwPYWKVNDom+3RpCUBCTYiuEl/xhF5T8kj
8tUEYYF9q5JApXXlRU4Le0TKBfyFlJjzxxRTRsTj7hF6cstA3BEhrdYAJngXGsMC
i0rUcjCR1FzTukbGYIvcg/j0Y3N/p3+0MNaCWQOlxvcBXf5esYSLKYFL5pYUH6XK
TdbUBHYQjdKvDEFQnNHPjflv++bB8Am7ttzHEZNxuPowDSOW0WSBO9UDr8GLVQia
R3Ywig2OeW/Kl4rzGxi4gKqyRBMWvin0vr0Y1fHnKvCMIEHYn6g59N2SsJ+qjdoh
2TsS3PNl65895nFkVI1L8wGnm3rr4H3swbOejPwKGyMDwxlLTJnX7w7xcySIdaLs
IhAUXXEtNWhenghl7m4cTrCHTgQOr2ZeZ/tVmeU3AI2I3c0gjieG+WZhQiKZ2WYp
NkUWTtTAdZkLhUXwFe6Ae39IQrIA5r97cBd+qk2/Tet8uPUWN7bKZrYEoCtt7BCn
5BN8M0O6iSuyJ++LUnpK2yEVXOJ2TjxQS8ndmDjyLpzExyeuzw/SrHHx956NZD08
jFPisGjDsJq43pkd4tSlrlvhZr/Wly4A61Dx4zMxxSUGEROkIF8/PGTgXTOD3NM2
sUHirWDvesS+Z80d4dLDWBoJC9T6MeQs3bNDD8C+813FTwk+TRnfyBoVvwwZXbCZ
JtxhJ60Eda2b3SoLwcDcE/lFuWWprpapvFS5tOruMoPp9sjm5ESe2xsdiKnotbYq
pdZg1GuHj2IUs4Ik8PNnJ7N3NItCIQbgK+N7KieZzrf0UbhDD9odxT2T70c3k7qC
iZVbIwqtwivguL4N/2yYC6gFURMId/B2nuS6VS8afszuns3NNOlhkl8hxk/LxcQ9
YtG4fIkcox4Q3R0yGe2JFB8z3UOQ9Fav+CyepBCh9gD2u7JwjzeSQnmO7El2qTsT
wpVTaZ5+1V1ZEJNd2paGQXYEHspaTsdhNqQxP+jFh5e6wLKQepCmb+BSX2YOfwW3
u3RzCnCqSCNpn1fjcYE5esUKbkZZc8iCJ5/5QNBrCwkiQbZezCdCyYz+a8BRLUs6
TcbvrvLWmg3egyIWM4XYzqGk21G9fFhvcqECrSxQEnwpEXRnoHKpo1rKxlvIOsEA
NXQ2xDvbV82r3W039xXQgcq1z9G2wWiq1/ELJP6++7J8B86j6VfaxvVHmtzHyDw3
McA+SndQ+IRc177k0R1YTj+WUJn/+3Ujb77EonOLcxCL+f/20yLQznVRiA+QczO4
cm5jAVnrWOS+AdpR9jBj5nV+a7ULnjEy/s89JGIqVf3yPhfZfGL0JVyj8IDnxPle
hcWH720ZgY20oskAOZBBwdWHjmbnfUwkOoOkvc44G/lXIxF6UIPQTK+KwPxXFTwE
/CMozcEF5KvOwWbKUWVYDaRDZEI6sKGtXPRdJoyc/hon/LM2tpkE7vLJX9WH2nna
Cyfo7tf9q2tB0yHj5wHFyxcNJxRlGzqgJMg3fRD2uyQVtznGqmkt+Ex+dvoW6TZ3
AF7Ac33pc/hBnkSNaxAmJ+CjNBgcrnpAI46tMccyBS5Xafwqd9vkpxt9run9lqAX
zwYCmWnCXc0++7jMQOSKtpGdXKnPrWv4wAPC7ADbjpkUZe94HLT4hVzE4RSyImkK
28BCrzxuXnvEZzOBYoE/reJhpQQVV9Ip17zY51tlQFEqc+Ro8k0ly0oKQBlk/Krc
eryShQt/bUHr5Ekaf0Wd3BmBSxWx4mfET7xB7q+1UPDcxjpmoHAatnhZjYqL7hNZ
JRMN5e6JCndP1spmtawWTrOnAzb1H6xIWpamEzMNnCWFtjaAcq2X6BOXZXDanjB8
+98yGE/STKD64y6/YBDgQDqUKy4BqBut10oZdjXpTfbjib6wivEDB5PBPEzOizrj
Z9MFmsVtCIUMGfvBow1gB8rHYULXf27tIXaf61lFAYsfBemFXL3z/0+kSKsgFk22
BNAWhgKN30nPFKltiT4g5cZLkK2jMx613+FOK5ZNm8Vj2Pk431nryLq9l8EsAdaP
pu+PhIGQbAaWyq35GZB+S9EKmvXW65Kw8pyF0yKyd7i8rqqQJ5sYlG5+yQz2LrbS
iilQ4n2tgIC1DLb5LGY1q/hdNj/P9bXt5NkSal1qKPE2ko+OcIq+vognc3yIGXDd
2SaFqSd4fTk4VQymT+b4YH8RyG3i/XVlg5UYmAmpGjc5cvTyqXQ+WLq2+YAzi46D
HexTxRqJyvQ6ZNcrO1DCNPwDUxD1SYVCd0WLV5yl0ekoKnk9plp9af9EpE+J6gvZ
Kz82/evrBZH5AE2aRWvIgsALI04K0+CVunc+asXLtMBQdxZoUgTmXNoakBHJFivD
Dyqt5KNxlUxZ4MXSEB57PxkDl8uvVf956MOc5Wkit0IsS7sg4750E3eetKWTx23k
ZuUfSpVYKCysd8YoIB5WK96GwOgf9KzGx32iiwSC6cdMh8OzIq/VG/kwPMOPxR37
+/+wSWN+B4NAr+d3uKkN7Ui2+ReUvIQEypqC0GqcbDfNZHg5sy4BLrgyC4TYQXwc
GwgSOHuW7ZGAuqwM15cAuukbANB4N9i564Bhh7Oa/BU3Y/s6KuxsGMJRpI3kSOpm
5lA8m5RlSeU7aNbrslW2UP0PPSab8bANEnHvoo5DgM7Qkcjuke7xM+ffVmWpL2IC
1RlrMWTmaZMT4B2P2K+ZQArfEEQjAFKvmllzdx7Kmcyas+o6mktxSUdFj5RV3HMC
NAMys1vPGt5NfOe/u8S0KtmYp9UGwt5qs0eSBT4HZPaWwKmlI2gEZ76MYoJ91RSu
hbFZT4V83c4Gu0vOA6Zsx9cGG1I4sNRYnktUAAwoFNTvNo9Roo0MpUvbw+Xrl7zg
01b+imO0IX9AEGnB6Za59d59K9rYuA6lMXRkd7jYv2zsZiV63qGLWgalesx0A/6b
nFCV2qd2CYoqFaqK9VyOHowZvNon67FLZawdborKA79PEebS24hoMZvA5TTtBoty
7dr1nYROusv+/PRxMWFAWVJxIvNuZuHgPFlGjpVdafmnqhRd5/IP+avPcaPdseO6
gGv68Z8lELCkU35t8m17+DzjkW8YO6Ozw+S/1FIPlIO1HKzkp/zH49L5K1xH8MX2
rbYpmfZEivaD0Vk51zxPcD2s3ufgbCRzh8Y32zzyCnG0gzXwbN61w7pdv7KSnpLZ
w1Mmo2/OQiKYPTMwaDhE/U+RhsDFiidNy/MtahW1bcRufk+JvMTcPLKB7Epgdwjo
TfKvZhnEhEKf+hIVZYGh7OVp2SvLUx31Y5hd+9xpOChfPqJli6F6Z7wCmUj+LyMI
ccftj+J3D2Mf9LHGm5LKOV4Fc2m7UcqnoqdeYewSR/p8AeixCZep+jCfjEObKCEK
HxlcmepjpimgE7/F0A6TDFSGCpHymXGvsb2Aq71WvFJQ2YB+NiTjs8Hd1vTV0Xcv
79yufmm2UUt5BVzXK8bNb/mnKD4ibqNOfYnOsTTPJcDvL4jzLgK8z+CHuggDbj6Q
tVVLOehlj4hGB3Iv242bUTILTd/F5K9Ru9MseD16+xJKmekFFz629vS7nyWp/goa
sfaGIssp/VTpjejzmONz2AblXM+0TSeuOUreFO9O5gL1PWagNZPhQaunlV3Q0MRG
lsGRFugLybgFDoGuK6aMsH3pzsNXNDVaXyww1/ri4AggfK+pdb1yvsPJUIG9Zd3w
g6rS+FuqvewSq4zAaFXAkpqMxH1JNgdxr2qTLXqaZMA5TW2EATJAIpD+5A1S+vT8
oVEhfcAyNp+VWGldUASLpkRORZfyHatS5yj+wE5qihO39hM/FJAVf0pVyDctI7dV
8rZoD0ymlfvzEuFRfcwwDiurL5Lh7AnjZzgX3NSHB8mQO6MM7wd4+scyZEmnMZeD
rnxakXlnRKpN7fInvN2Y5P0avik+LXw+wYMHm6xZ05Gr0QARy/7f0OPcvDVYkYud
tkQO4vvXTXaACfTMOblaPh0y036Upmt0PphdxngwXtmWGYjOf/F3qz7sfOskstG0
kQ6UVSXxyiMz2p8Gm8fKMx6QG9vhkDEMAuxvJazRbA1M/lL1xMfM7pQQaz2pliZQ
Z5vdCZuf2+mzUJiBQuWUi8NEMwCeOA+I8OSMmACMkHlm+wQZqcIbN57XJXwuCDZp
xSFnibLuUefRq5ZTFPAjtZlThkLhWq2lzWZ6Un8fd41ldftR73ZU1y0975u23WwR
/5pIqj3LtM2ZCHgf1X5pEw86NmxPJITUFCFBE/ZWnhHMVqvu4BAfdn4EiwSxUvv3
amjnnIsAZ/94mWQ4379qSK71kA7UmD1tiw5cLa1DnqiRphDmQPce8RGgOQXbvxQj
d5AUMp/Xk2FTKkq1UM1jzbKYs+WYLeM5FFuUa8NSFCWlM0V19Ua7fRNqMbHzRJVl
rPZV0nlQvwkt1/bXzCXYUw8pz5D/L0WZfxkuVqgYzRB+F9cGGRqpnWlJR/XftMYs
q5WuQz9tgWkr88rCleVJ5o7cXFZB6DAKNpXFmfmnVXQoZmbmmNGjqIi1RwcbciLr
R+Ftr/p8JkVkmHqqmmTJZ8IHl5DQ4vq2pIR9UyqCSLTY5gZl26/rc2xxPGqsZRLp
HzTInLpsyvquJhjMMWIjGT2m5BjVRX/tPS7xjF+Trv1M484tLqvJCuRZx56zICwq
D3t36ZEorLIRbWlIM3PmGD+dCBmEFNMIDc+S8tL1Ue0GzkC/PRvmAfcfu7BwGnwX
9I5weR62y5oQ6ZNiz8n+I5nbsk5VnbEdrUWSZxBFhePI5FV9hAskJPUVcguqXLAo
P31h/UAa+qjqoZXVVF9hit2nR5LFkQDTLguMkYn4obZ4NttNa1FUk/Q8C+gMadiH
D9Ee0tFaZqR/8dWGFfL1r6Q0B36iH3emtnAmdikFaCDkXgDB0l+oOjj7/8doBH+5
aUdHit/ty9QAuXs6uIXFP4kBomT33Eudgqmygvl9vhJDB10hfyUCU/xC+7dvZnHw
kEdcLudhuNGNaYpRAtBdyHnMoXlH6keWe2M4d0IPXxODuEqrI+na1MSDzSQdBkVu
c3kMBZbdA/eE6p/75AyeuBp8cN+WqLoaOuCJo42XO10crxxiMhPhGd9zmC11Fami
x/0dK1xVdamog9u7u2J3/lh85kHJepY+TCPdETMhngnJKqZ6kTWu6O+Q5gYe/Bwi
+1sLtmUxWE4zn5PncX8DTggwNJ58lL21Mh1of/xxOmOrD6cfCKiFcSncWUvGP7Wo
V2Ctwsi/0tc8t/Qx2HpyD8pC3Q7ijhLvQV8vTRTau9+TOGz4EgYcG7+l1Knd55qE
Dnx0Gx1zuHKoUoWZoXMPH2Rr/b1w+RcUOXvryDt4xX/8/WOokfgNqqyi4g66MFTk
BdY+gHT9P6jpQmiS1H+rVhuh9ja6ISiyX/dx4WyUELELu1xAboXrvaRG0hxwzkde
+zjQDR+eRrsKDhGilDTUmU3bVoP3I5LbCWjfGsExTjxew86uMJhMnt9/ZT420pR5
nkrmURlYbcBUaLnopdLbSYOlRVa96X6Q6po8vfcBqRqJSPAbtvFdcF2cyGzWFzcB
wxy0h3IO3MdLLeHeSk4a6MejfCSKhAZ7QmJjyODAg6AoOWDJ9q22Jw9c6/2LJPz4
4puACnken1cAfyT/eOvrwSSTjZl+uMAUnSQQY/56TBEw8rT08vv4kYgMFObddgdk
fbCr09wxBE0Fn2Lf2TYlC8mM1Pq5j+Nx2L8sDnBaHLlsATEiGZUilITaAtzyLvCT
CbCmjVhedHwHucZyXxXFmtWjDMaAS4VQ6WiwmQ/siQk+OmQNrhQ+NEi/80kNz9wU
Xm7FlTo0mhe9tP+9a4OAZEENN8Szu2vHpZxk3jd6cDPCgwq8dLobo2jNtBPsl9LD
fqe2p5Xz5lzA18/P6XtusUQJ82Zao3fWvkPPlRSpgF2Zsgsb/aF6vd8rtRNO6uDL
I6MRzimy1lWbLvw5RSweJMnakojFFgqfCjyo1I+NbDqCjAOWHrfq9XiBvDW8j5gx
eaf/VLMJ5/02zfhWlZEBhXVVDl+T6YfiiMpCQ83ROLz1rsWhyfB/dEqUnssQ2icd
eCVATRMBVVG6KSForZ8KnYME1wIJPjLEsQ2cjlfc8LtuR1ywguCso1Z1QUZk9/+1
qSfujlB6rBuxPyf7YMjsNc9/JH5s/Z0ZyhwdYBmmeEAJ4LhdMVuoTfKbIHFicCVC
cPz6/e+nFZs5xcqJ3EabaG6zanycj6VSpbjd+46A2WIL2oe8ElwG047c6YMNTYE7
wZ286k3OBUuRa2DjYM12r0E0M4ARUxoKs5WpZ/A2NMGKf7VFuaosQHYazseVThzM
iKpnJpjUvcXEqUFBYx8LfZ5gqTOjo0qjhFPf3ICLSXGzkmu4lBxiopXNOxYkH9/c
bey2hH3ZWftsNyFpkNkHVEY6QkHtgq4WB9qI8PcCq81/NZ3mJCciKZuOPEDRs+pE
aeghTfi5v/BuaJ+aj7MrltKTscy7WlJGsJh7hVS+0Gg/6Ffr5k8sYuwBmDmIdwrW
5Y+kijRp6pXk5rEnWGBE4F+afUd5YOO3mAhgWn3wIgeZL1L0u344pQsiFI6v/Bbi
sRVcnekvOIJM3NwRXIyPlis/q/4YTHylcSExHio7WiINW0rnuZtBOjF6J6Wuzumg
WFO8WAkwiT1e6LL1Z00k87hL0vEu4T86+515DyYXQ1AVmGDt+WRGJuTLr16hLvOe
LAHKnRSz2MsMAOHKGUwVfhzjjZwgjmyRUl0zTLFs1SBx7iDAVTki9qGBJGrTTkB+
6HXK7MsAI5+Hq5qLaLlJ34OUFJfJgN4X4o4IbUg6YX9CPxPXDvS0cT0ATWdP4Ps/
iAaaA+qhSZp3loQw0q666IxBK45LPHydQ68clTGbrHxLBndvbwVw3T5kcWdqicPe
zyzyJsIdc97IL8zK93sromLHILFdlMJIDpmB1sFTauLkTkr87LFDcJQODAp0Y3Y2
u5H2saZzRvWZxiEAS0MlAcO5BbuOzaCR49NtK6srdQrLc1JnXp2yf7EwejcZTsIz
t8SlMIU4q57IO6RxwFyNFiOy3hPOBDLCJUbXDQZ0nS9GHh1zgpkq+IoxkDG5V4WO
sMX+Emh7v99j4HYNUkdd22HCALqTJm2VQ0gWsb7Fpx5XdhwJIpwi24xvM2sXLO9T
SP1kcNzZrdXpi0f6maIAyZy7monEod31tPLwU0i1qDUWuz0ng81OYnKUOZod2ocL
7mIyehUDXxuFquUTlyMKP0wrpICrc7U7SAt5jYt9LQL/SOHHm94Bopejfr1bz2vF
DHUgqu8YkQBQqI4OCaJAD2GVnPXNWASQV7KAcBSyjO2JbA7eXmThP1ZfYQRtMHds
41v3JRMwRc/3rM46C5M4Vm14ZiVZu1Md3jSpG9XDxUemzk/p9mgyuoS0nEzBv1Rl
ToCjLzdAeUjpOYumaa/ZAen+XGl+u0pB3dzu8qnf1hNxJvs67Nlp/Ebde1UGoAod
oEM4ncycu+mV5wSbUAfabEbYy84GbHNOxaWIibQDQ06BzcqaokFRhX1zuXUoh1IJ
hTSr6gyUwIsyLXj/+K1lC1bwrBcOQqVx+PyBR1EbeylcPutw/LHLJ4hY9DwUkDhE
0MupOzLFUZQivmR2nCVNd/3/+FvmGGw2OJVCcA3RXodFXUCZ1hkEnj6+Ybdeph30
4wLI5nK9J7ZF2JOwpwT6L9UeXWQeKkOzOfcyqFzkAGzv4hYuW+5V0nzlL3Z7VXHt
RzZIJurHrI10S3twwhz/5nyMYawfpX3Wzza5N5P9++0EAogHOFLgR+pMqfo6Z+9u
+j/qAojCQMaKgL83eVEknPn5eEbwG24BonnnUCnQLaVIw9Gmy1ERPGlbO3VcyFAe
SjQo5jvRVwBZCzc0jM3sWw4RR2xrpw5AMEmberTkrTzmy7vT+Ny79/GYicwz9ftt
dFeORrS68UY5m9RL+bOZ0RoT85DNLMBzbwTcqyivi8mwrvF9qgp6wPpkwQlTot+k
ThOWqnka+v0u7bDQsSy8nj51A7rLHAxfzBE7CdCbRNZYDAG9Wjk1YWmC5ZqQrxYp
dcp+9iWCrvyX0oLva2MJUAlUjnryji3PQtfBrOkXG4vmismqseQ9cMJESEaIWBQ7
PPiNhkHNfheld5be6PNO+7P3QQczJUs7dNuD85KA5Ehag08nZtfeiJ16bu+Icj7R
pkwdTX5BRMBZoNyHpasz9AgdOTUvWSZMZxdK94QIRkVyZaSNHHH3jPSpa4DXLY4b
o0jP9eSu7qPZO5e+Yuzeo+gSmc7K3ltYVOs94Z4f+X4CBeNdxRbAciQquSP3KyFF
/hgBFBEY2PvyzdsEDN9XVGQ4WyHhKsekcdMqv7e+8SNHhG7UvGftbT95t12JiLzg
n8e0ajIUPtSY0m54y1phOKVouI+2JK5nbHFvLneoCUpy5RZGsZPxBsjtnrGzcfT3
UetlBD0sOJ+ekiSxmvcxtC0zVmeSP6Nyh05zAgp01t5cFfF36k56J8yBOqZHUlxg
SFkXnUYrM/VM+KrDesS+VBDcPXS6fMRsaod2vHSaCyzafMETvQaeH0uAHuE3HWn/
c3EPqNsO/EwSJmXpWRBSrrjTEmxL1MEk/hyqRGCg9T3OPjIeefUgLpqOIoWo9Zu3
mCliejRCw1UD2tZcvmgUCecGjHz/Zm7rZ8kJo/0jSk0RyqPNYpASEdU0jAyGHxn6
yOqnyzM0F5QmboMzJc8aDkO1Z7F/LN7cBxp6tF7yljAvwqex/4vKFOmcPBr0LH/7
PsakjpK/cv3FKGDKXwwKCKyieEuJqpUIyI6w8xFsebf4tCxtUv+4Jo12lRbmYDgW
e+mL+y/EtRZnW4d8ibOexxv5w3lFTP8idiQHZFbJnFIQK77UahjpJLi70th7AiEv
+yGmjsuw6pMZXXzMQK1TjefT2G/+idWfFCURrla0QCuuWqRKVxqkbbS1rzKWZGoO
F3UoBGvdMGXPnTBp8sxZk9Fs0z+yOAIbADf82EYx7Ehc2i6nADPD1HDXqbRfDx1+
iWjmHA3Z5+Oczl+fJQZH4Ywa0+MtK/dBdK+KVDIrpBKdrV92uh35y4Eq3+R3fQax
EVb97r7HSYkG8JscmXdhEAe7vTwxvAn4kDE1uPO/89g2ejCxd5vpkX9NXJ+vd1Pt
pLdRZaamCRfI5OGGopMB1YyF1O22saGIJ0m1zyb36GTTX9RNeLfsFCX8xdI4cX3I
7MleJTDEoyLNW+KdM+fmcOX/rNzoJGURdW972rG7GJf5O0hlHrMho76Ey1c1Ne2t
t9k0Wbj9dHT1CFzNxhtFJHN4oeoLyKGOOHKS12TWvRXN2X8HTTcHzOMK0RSGIFa2
TC0hbn728i41d9swM/rgGGpaqhk75hLTKTZXdBYIC1K4sZOqBBdxyjWGgas0Oc6r
5cnXaxOodZcLJPWS9IZC+9lNctyH24yHA7DPc6m0qltkKhHjb6I6LxXREYN2bKxP
b+1MyTfMg5ulWkgfEWj3RWoehnIRaP0+RyOZ2tReWQS86VszKAzXdhuWb5A965lh
gDZ5mO8QPp6JZn+zQea15of/Fg40uj4jMH6hf5yne6RZPE/btKXhB4E1FuBV0tLa
lQq8TgCBoQ8tRMzw01jkbNRhbqj7K03M14b2GduTIx1j1PHjm4QLugg9moovpt+h
oBaIuqGiP7tPs619Iw82vFdJD+pIdsnGJXWDejAprwWhWkMRsVmp9YAIumFvRKOZ
57W4GNupc+pWy4v+0BlOhm/HI/bRY2c4vOTzl9ONuIkZ/41eeEk5562dfXDcp0mk
JaHtfbMQ92nl6ImXdZZdb+7ErhZQv8hHj+RJ8HqxfQzMqye7uSjaV8kYK943Sjex
nO0sHYFVxAMoGGRZfpzMA+KrcXkwzBIRgXw/nDeGx0lrDTx1Ggy+W7PYcRlItV+r
nqDZwRK5SvF31tWxq4Y/ncC9IVMz/pjOxt9cgWrTcA0hXX/F2cxD1TYla5WBNMvE
p1HDiGflFwGyjDp6CMeEUjvhOmgWPoIXcgjm8kGusP84byWBMEcX9vtl6zDIzslr
e0JW81+qnOWBEch6sXDou7IipT/6g6iOgVHKeeaXZnY9mbxkCTYEzExZ0VsohwVX
TqxDoz3ZaqGKyqKwVOflqPQqH+ofd+EfklB5mhKQY6JniVtt5CF1ZjzS892gj4WJ
Ig3whQZCq1osR8Dz1P4OtUMc6E451nvxnT95de+CUDZKUWYqyzAFJzyhv0dG6gV7
Jv0RANTWJmSeQe/D8QwnKAzzZAnqMsK0cm4WAkb64qbUyHzTOHfeVmNKT0DFDl3n
PWJNOEGqmb5/jfNxiT9DVQcz+kX8hWKySOocarbe9kAI1v+FG/3lbGdP2EwP2/cM
ffPGX9xev7OeTsW7JE9zcgeL02v51YuDCl63CCz2izVBJrAn0ghWaAdDVOC5Ckz+
H2VF4q9mnykahs/r8L0afBFKKpP940yirG2fuJlU/CFUABvqNdmVgLt8vPPtgaOQ
E9msOk+opC5+zcpp0SHON3mgOSYY3tzfhhcoF2QcylE8vk3O+LL0Uv8MNkrueHL1
C/kfb1HCy+EM1bdV6ZPYjgK/WAlir0rON2UszZJiYv4ZQz/0lqfPoLqplTJmnI9K
LLdEaq4CP5dKC+UPA/kim0hLaX2p2pdPw7yEpOfpCaOv/R5++bAzisKjmAoEfV5L
FZ8xa/oH4Yvib2Gkca1k9kis2Tv3brYcJmiJ8uZAuRRuKd9H/PzK9zgdThzPoCnJ
gdchQs9ac8vxaw0f77cSb2z/vOp1U/m+U+9vc1QgAj0ew/5OwW1lwVX2jcm4oWlj
WW+AWp8hoXQExm5HTtzZjPkKKwb38oMO97YAEl8UZRLL0zjwo740X/OyzAvrkWMI
gm9MmCuj4GUdAXV66g0KFapTmUCc+TmmsM8TlU/uoL5/dXn/DrcssEkmwd/hh6Hd
hjxwf6DNzWcRmn9AoGvoNXGx9GtF44FDs4v5PQb8Bj0LdJeQwb/YseLC2x/v2O/D
pGWbhROHTyYP+NqgNI2H5LyNtUdUih1D1YyWN3ugLbmMMoUM6BmhDASdtYBn+UwS
ElRORu0RrDhLSKHRBT3EbRSr8eGa/IHjdVuWhk9xnChZxG3ckUYYnJ04IHxL0a/6
QPVm1FE+eCWhJaG/0t9pW//qZqSzRtOGGsFiRlSG7ynaR8xq/o+zUIIAYxlEBqzb
/d0QRUelAbQvqQP4I9FckeSqdSl1mESp3LT8/BGDV4/sOeLdiqU11YR/miq4SK+k
F9nsUtYk/NzvQBYnlB8lvnCpdNHpOEtUvRg4IZ88iXbOcvjsBfu+qINhfQod6glS
sdDoL+J28lPYOTFmOENS3qR8EWIS7oKC4w1PLDSqrAVCQbkNxw1W5vIqTyglwJVk
XAIrIkicmnuAd636XoCrBuQtV5XH3dRaC8wQ8mGB0nyzhvZBUwKA/+5yvwRxSAEO
Kj2X5iuhjCllLgcaWZha9+NSvY41pPwVcErnwBo+o0cyxeibdJGxx6dzo6wBOMug
o72XfkqMMhY2yMYO8IBQCoetSZUqJDeLDHweBDXg0MvCtBiYEBxtPLLXcuRRWz0z
aosBSZKbmRaHwBMoRJM2oW8nIF1Vt8uQAPcczO0jggUHIqOkKAEJBvO76pt5bJCS
7eSb/bYoO/zCgQWT+leak+25Vy74j5dg67FezcUNY1LumOju7BKTBCGW6Lb0EPDv
zEuD2GyRcYlbHN+i4B/15G2OPAUgmQ9kjBbOa81TxzF9YZgXscOLG8rqchhK883t
Eg0ii3fDZgErb4T0EwbSiaTJcI1rD28yO7be8XVIRFey/bClZGwsNSUJk1yC5eXl
IdF5aaZItsk9zQM9K3z5+kGn860tdu20NowgQ0dQfzf3J4NuOIi7TWEbvERbJCuV
vs/Yd8HOjZTuHkNy8X/ri5C1ipDvqRDKNXTmI8BruQXKByhGKnkZYd7SxuYcHu8H
4zTpDquY2CXB/uc27GHZhFvbBDD/M3FocnVN/EmrX/ti3OrxC8/EktOkgPSv5Ny0
dAdtC6B01rQ43rjn7kBVOg3OPYcWZO1SbOW8WsfYg/eCGTPeLy1z4JfEigZSYi+5
48WIadrpox72PZAbRdpOxvcU4IqEi2RIniFBQAujvJ5Wd3ovyGUT05ojXJHs3B0a
Z6u5jLjytKot6q6/zX9AEDEoEo+97NR/h9uAQD1CApS2K5VQbt5S50jY5F0CILfc
KuuhQnDMqS3nOgCPM1daPSxJ+fm6ZTpxBAY3lRWvs70e8y7O+4Tx6umwm489M8L5
zzEYSvr+JM5lapbtdoGdkAvwHdrxWxJnazss8dJJAkuV315Eq9D0Fzg8d+BigRhK
8PtjuuSK/HMa9pBJ7umw3/jVjRU69yoKLIlQKGdZmu9knM3PRqTXpLS9YspdyDLH
Vc1IcUgQ8//dclFUlOKrwMrkUxOGYOTJXARtv8urLgl41xpGfTrQgEd+7wQ6lD8M
TsE01wr5pxFFWr6X3wAi85CEgmUeN4DYNKPy3deACCBxi/qzpRLEvOgWYbrkW6JP
f22Xjx4doGls/HLyYyCN093fiRwOP9EoSAEQZBMWZ1lPFPjjYGTd+iAJ7fxwMIcW
ztE8+YSc6BTjuoaugVTnOqA1s4wsNT3s2z4bPBKf4bNavRy1zbGJQ3ItW4B4DADq
TBhkFELwBM/9gPO/hInUiEcko0+bPJSmJjua8Y++uSFk8jA00oer+SlYPuBclRkE
HOIbA6XHqs+xbJ1qZt3aNjqGXOoDEPNjXg+iMo+yrl9Idz9bxQH2MWQs7kOKYu3N
bLVeT9AGTL8ko4qcy8hYmujBoH3n1RWamxwv2q/SGoFbfQeFAQQKJ8nhVr+uh+YG
5SZW1UgJqCjiHsbRDWoeFcUScmW6hUZa6YA9ilT1uSkHvDdRyMB4tAp0xAHd1XsU
cK6J3/lzRbARwI0x9xK3MvmFhXRbTpzrInuKNNOTNfixhSJF0Oyr1oN6Y6KYS1Gs
Ln78vo2TYl2XMKM4DXcfLoy73yLuZL0ATojZbMZB1xYcZ4PQ1HxVfexJAA4aySBu
8o1YWcoHcI88S2klmEDhxIIKyg57ElBjyuULUHiJCrQ6WZwV2u/yI74HpWIfzq9W
LNhG3P/VzMv/6rNWmCyNjliB33lNKhb6eXFeJ6n98LqwtVjIcOmRf1oI4SsagTdP
XB+wvYGnQ6CXbYy+3/j8kW760A6lL7XhZkB60WC+k77WqrDDyCLMCPdFXcLQZeYy
wPo2jtss7t+vceDnPiL3f1UUlT2WwGACiYxnVLwppfeIgnPzK3z/5ZRcMM7IcVZm
2OJ5ew8MDwWltgDAcbexeqSKD7gUVE73dK0je6UX5Xi+AhR2bTyGHVWC3OE3DiWn
6gYm6co6OWjndPPSigzBTG6+W7yg59cGKP72XS8u4Pvd5WrgG7g/LfyBVP7A32yw
P+jalT8ljdXnFYcGyFuFE/Ujr42aaacZ9bbq/17Hlho5YVMpvHmZMPYB0agLo/vn
UKGRDNr3yXg4mAXwsiCmlVTbLN9xo/3uvsei9ms84jzGpw2LarGMNXqzmYk+a2CM
oCM7kPRlAklLW1TD4qLqXpcl/l1Mx5DCkFHN+E0Uj0HprJYl/58d162JIWBODbua
kJtJJt9nLJ0TIATGv69u5UUzXBlrLnnxTS3FPRNVbKmcRmlwsO9KyegzTxSiPtYW
RJ4fRq4riHjzeAWtRk/sksS0m/Dl892qkS9t6U0L7MBwsyjq/dSIKKg05S8GAs4C
vHMq4fsNomwc2lplg5ihnqh6N8lPDg3W4Tc2pFTG3HCoyph8eID8hzasbZz5RCqF
V4ptVyn0yP7rrQ/on7Q3QJBEZ0CpdLY5PQg+KPg/cTpAOIN8XkAj4CUHSKlmXCZO
KqUdj05jEgFtiExahe0nn7qMhasITSu9p6knC/c33tI7McyenwFkQVEV7BhrIwTt
QcjmOYqmBYCC87qugDlI/upVHXh9BhFIgdAUxAThzS3xFWrvejJTrn4QIWbhLoBy
rptVeQ7Zj+nlTYkTLvH2VnZiQMKfKI6LxNR99H3vcEAXTg/kGTRDjz/3sJH9cufM
bAyNSntCOjthg6Mbn4qMCWyXXan1qogwqOBwmQYwNTd5gitSUxZS5vmVL6avRVw0
DOxMSC+V1VCKqzEXugzx3Y9P1l9adynDiQfEeJY4v42tJ18kb7NDuhiK5GL08qDG
JIulEju92liZii3f7VfHjqzeR1Mw5OutaR9FNO0SHi+rfc85vybNKnAWHiYbCRTD
stTdx7SOGFODMkDH/DUR0cCxMkIIkcZp4pDOcQLnd/Xz1MLjEgUycoCDF4hX+xmx
KWb8vs2i2kBZtxJp8wtO7bR4aEHkwIrT/HTwHxEjq8S3rlR1ZYIj6cNicl8NDvPy
vDKbAH6w2bhakEdzhsNr3u07kiywnK9/J2XGHctXePGx6om7uysT3dMHRM9SdJSm
EHFQ6DcKybA74p8eFCb6xhpa5a7rdvvViKGOU6+8sLoDcCMpAg0htKEHZ0ewBOVy
yyTsh/6KeL6S//ptyA1wj63fJ/N/VklmN9skjhukkJAepPR3MvdLJ31weiiukTPD
0OgYT67Ga+QWNN13X2t8lijbRlvkNf5I2kUH01jYSlniRr6MoOjlDPkZRYntj8rB
MV//Ej0bVUY89K7PidqSnqGLF2nqD3o2WQJUVuy/cobsWWHOGka7CmQmj8tajId5
5+YFmia8VlSSib1sRC3qLoYDZ+p59NVuRpkoT/IpV/kyu4ct8Th+UQHV4PANElu7
l3vty284n8227o+pL0MJGEc07vWvAj957mPcnx8Yrc7+XJ0zEkyrd00DPqGzC889
QdA2qbS6Q+KYKgq0DO2IVj0FNGJQgYLvcjMaTWWYI7TsFxcZt9For1ANee1WwCMW
0gE9CFka/dWi1K+/a1iDdUaU208DuSQJsiwoIAsUQXrOMGEGkldUxoFELlcHu0yd
GDFpw2P9pxGTWTlmaSUrWYO9VTYqx4XgLneI04TaWr5CGS2nUipmn9z4PADY0GST
6yT4zWgxhQRRlgMUirIrw1ImysAqCrPGwFpWLleaBuy0qShE2zm8wFcVbmw0t+R1
018C2Ju3rKybexbAIS0Dz3eM9M6rSgVNMf+1l60PDMVfN9UPjG5ahInvBFifxvXF
CYeg+b8vo9Q+/qW+9wZGc5/QurAc3Df0MV5iLN1M/PfEL86+5QgCU0Xd3scB0kZP
Bt3W8K8Qqvmaj6j92aAmnVoNzfQHK4IRqd6CVomADUNMOzUOfc3wsI0maMPeml7V
ZRVt5Vh0utBvHwgIeCaK0+GKACtgbNW65Gse/KiEUEWedq6HyfleQJth8Vo89v8d
kyaPhW6XCSONufpEetIKuOf4S5pYjExi3tE+eAbkUHIfnREBb+2/Cxq1OzGzMx7f
Q3OmdKZ8lB++79PyK+S4o8E/emIv7DQEUCCyUuaOhTDXWLGOaTe4ocT36CLe2Uq5
nMq3h9bSNpjdq78W6DhVdiiztP3aSADA8A9RA827n6gggs8CnHSnyLMhUlfGl3vi
HY1xzx/ZblAzcpc/idlevNEieKuoKAbrDRnLZAN/fYPPs619EPE+Uo5L3Mfzg5KV
26Ec6cqvkPnDdyMm9q/l6P5xoPBEOUQMzAEU4usa4I70PtXQdYUMuu5E0SzEiZf8
vhkF+ea3+168U2RDSz+EwmOzyr5gZ2VEyOr6opfgeRmRfGgF/g6d2ZiGKtOBjtj4
gxCGNncyW4BUzmLGBdhmzc4RUgny3kYnkjjSkLrIuhlmFQSHOShZ98UMgTV+1Adi
HH3RNPdU53TN3bCxYsIu/IoVdiAFxZf5ApNmrUrrP+DdIQLuwb917XNLM3kjMr9l
xz0iyntKFabSBwd1TUMLr3mmnA5nWLHhD+uJ58EmkUiGMI98FoxdY1CFShZ8wbT4
30p799gs66knI29Ee709HEkQbDPNypeMRwttc7ZSGrK4SPJ79gMm5BG6OWarhzEk
VU1GOFtIw6jVFmDfZ93GqsOe5PC4kiAD3WEUDe3v63GRbArSov2ycgjunlQb8V1e
bTU5fWGodKSUCGHLIyvzYFk03At3c7dj567fhK+lnEqcF1dmImYRebGQElRuH51R
+eC/M0G7TcDImTay9DSyBghR+aHRyZLj0YbBZ7HQTqlnfIGAv+xEPcVF2l8RLQb6
LSMLcaEBgbZKiZGbPYN+EO5knLZZWf51mob7QBW5gaBnk6gxLJ45fa3BFvoKxIq9
WtITzC6loC/Au1ItUM5szQTkOr1wTxMcpxNxNmf02bdzYlNIqU27QqScQFnb490O
FQOojEz8lcN0HRErwt/h9j/AGedy2J3pUZL5ZOJ1lo6/ppnfQSx8iq4u7bchpC0E
QhsCjBJbXl/PEu+fEQ6ViRNhHSszGVyesq1yGO/lKmPlCNZxWaRHGEq0VQlkuEVL
S6BLVvpM+BMZnPSB7mRou8qP2XxB1K9ZnmuadDN2+uREYg0B5bJjEAXSh1kJakrQ
np8ilKDj2CQEqyvLehzeD+NDsVQt4ND5srO0Wz+jBeiLbvSdchE/OOCwwbzrjcrD
UNuge1k7nvB6WSSBsprMG8vLy1TVljRfhxRtrHDkaHidzfATUPl+ZKsxctLTDeuk
ZffAd64DX9S15ixsCZ3DzPF6blAtOR2bE9pDuegMpyQ1sOSQaDxaqZWU+KZZy/2D
jgebTdbwOJnRtO7GYNKyASXHhFNGImVRjtheYA3BYIZchDvEgTzzxCPlfduOW2CC
qhfMqNl25njl09tMtJf/ssYAjePdqTTV4sZ3zPFnTAAkqK64wGnfW+OLledLBw4X
9Nz0ggqCrazfwLDDmC7UAQpyt46X4oFHQ8ONW3B4yPdVAOKsVSepYb2j9mzsPVry
RUhWEqj+kbhccRmF7K/E2X2kjSRyfO2OwSXH2Is1AGSVRcLhluKRVJBIryGgZY/V
fnxHnYjJH4QPmkGej0VySkVloBkpl0HcBFy4WrsPAIn/zWom+EYw+saEmEbIxLat
HfUkZjtGM3ShwRDSitDbRK8y/8ykK07BnHkUF/2RupdmvM4Loqzmnj/nGHQXEaUd
hmfLNpGIrWAFuvFEQuTGtUoEuueUw2FePYnla1IvCHl0270USJGUkFxRZPe0m8is
XYTJ8ZiCeJ2AEiSA2RIaiG6nx7aC9ugwY4hU6fzLOpK4fMzv1Pk/GjGEEGnARLJi
qR0ymVNyFyt4tHeC4782j5RQLVYb7bIeKP0oTQpG/tJY9mL18SG0joBSJgUOsgzl
Mx3xUN54oH09BQpfSDQJGNdHaxwATYKUv0El8HfCpVSELeEM45johKJYBTyNMelm
Iab7fVGh8uEHnOHyBdnMOs/hOwgkog4QTZVkWWopPHOgMlCYv6N3PN0hhK9h1e3T
GGJczrjDC65gOplbT3yog+12zTzaBNnfVNK1pIx7uinLDNnJEUI8so5+b4x2FEsT
C+I2TdhkQlRm9S9sLEPbxw9ypEFj/XmBdKtsTdNiHuBHUNiWnHylnPgLA/JhmF1Z
sHIPJJ4ghfUcNlNJpee6+WN5qFLrhXC0pSDiEty9PbnQceRU3hVwDF1UOMKZ4tBV
Ybzidzmfi7QN7LpW9xT9rYlOCKsIO8OpUUAyyLVWsQXunIm094IYqje97SFaVwZ+
SouQ2zJZbZF0nL2gWt/vii9V4K07adtjq9shdSNUPYu9n7CrKHcupIIkEiSDDGQj
lO22sHo5bH5yKpJd/t5qjJntUoMtFtiyw+n/Zsxqmxu9qVRGxQR56xXtHx5t9NlN
1N63A4YYGFFSMvB/OHagT9AdHgaOipDNLA2h6Sk2ziw/UW+zl+4iJxqgIJCveHX7
wdOgStcqgTToitc0rKkMvQItvcf+FH1ppEuUU+D8lJn0zVD/NMvkH2l7h2EigbvX
bvxtYyV0MFO+Kq9E3wVjIqmFvzx2iNsvNkSYL1SZ/4i3ti8dldyuj2+E/BaVExmC
5NhmryAb4K+zBA1GJlg0aKWpsDNB/4JIblg2uAyyjwKEN1woEau7jNuoao8TbQ2m
NoX42Sq61D7staBwFfZWrQ/5BQLLQVWkdtqwLb6Ha3ecmDn35YnpqZ6w8guY53HI
2BeToNjk50JD4bXZwNQb1BkE9Wios+9JfD7PXcdy1UXzRfEWs5cOXijxhgbduJe5
CBkcYMpoVUEYYQtqTP7Q/l1a88e1TkuBel1Tew/+2m7E4t/TLtMw42H55SV1k06J
ntsPtVqPgCzbSnECeuyOxkjEg7Prg7xCH/C8MlbK0SEPa+iG3g+eG3thq68KEH9a
zRPLGVyhew7F2xdHCEr1I5JH8ARhKXKlvVZWA0JndldBPQGPf7CfVZW8e+mNmIQC
RgpSxb6eyyNzgz/9ySko7WoQXQXqttdIxGEvRFfyNaAUN76DrA8Q6FHIal7IlnoW
eWbVPUsx5E9DhjO/NU5ux2pGD2LAEbkTqvUFmfR0cUyUtXFKAwYPUsi3GIb8L+Bu
FuIXk7s1sCR4MhC3kFKiT8MJaBCCe3rFkDpQpg2MGagC+1VU6t3e0TpTkjqPdJBK
NgXsh2Lr36eKbfHJUvRPElWWkXVj1TkxbZqTRRSaCfBMWmgi3Ly2PYDRljacwv8g
CdSKTOi3zrE/80ZAKvjnItO0fgNstDrASHWS1V8cV9Wq2+trSI3VpVqL0Dcz3q+y
Rru6y/uFKa4LU7RL10WtQNEMXk03qu05/9dRlkaK/GE1nMNMojJ8u9MMZ1lrLvEQ
U+NzjdpamtHG3SJ4Cm5uuCedw+WirByARlbJ8QEhsWaT7DG91XNJN1YTwpFfklyR
He6ReOLGzVWltq66PATWDOr1dANgrh3HqBFwSATSZs5Jf37eXDijJnr3M1ZF8Str
Qln+17GKQDebMw+c6URDmw6lBLlLMBeoQjx3qKJBlTWv64yPLJ7H0Rw1Lw8lLwTF
AP/VLwEqAgpr4/vY+5GGgAVdUfqxMe+UUeQdwECnDYpFzWZVku5KppDLpf5N8hd5
cKU5RgroV/QXn5NXrEgkQJi0OZWTOje1aQT+X9ZV22q6K3+lHZyD69J5Q1ClYfFT
1jdKLnE+TvK+6nOm6X1WtHMM96pFw4EfWQszPsvfChEiJ3DTPRpfJtNAzWu+fcHM
O+BNdWppNHSRzF2GB4d6DwwWlXirNSBNtV/MVETvaU/Vn0XU6Xa5xzHpxlva4Q9P
+Ml83hJcSxb/1+BMz/LqFO/2tU13L9436r17X6N2QFYiXA1j5tBGdfbbWXaki3gM
uAXKRUisgL17Iuc+0ruYKaOO1KN0+9/gRyT27DKAXwnIJ5q2A4XIZODKEcizlbLQ
Ypt0SCYEIEBQdlMrVw93GSJ10f9CQEyV+VbCNPMWPlfEgOSr+yLdvizh2mVYHVO8
beGtVo789pEo9NqMT0yWdv+k2Hs/qqfbsUm9yKhR+CCofveKQnXX6M8wQXL8LyuO
6M6soegOHnHGL+z1cX28wN0bb4BtV+b/YT+2lFDeUXqWTgVf7qansh/R0H6cw+dE
dKq5tIUU2cDi3cF07JLWBnpNj7d9o1IxuawMntCU+LX/M65VykvixGpe+DMfamCY
5ZUafkepiEKnx6i3bgz/e4OSyJiRUh9zrJr5v9rRUrJhqlePkeswm2Z2YGFao25G
vu+u6IWY6VFJYhBOVfUERQyJqmDHlXmGwFBBK5LfGOHFyYw2jYkYwbEn3Iz2K4bK
VbZO5Y8jF4uxowHq/FIR+aBHj90Lk2ugfTXTXvYQYPPpKRZtHyHh79GL7MMvpAND
pRg5MkKALuQYcY1ArBN/vQSjK0vPL+ZAjC2npnGUolBYJEtq9JOjDQ1mpN3+19o8
huNbtefTOivF5fNFI4rzyzwsc53jd69AP5OmLIeEgRpXV5p0yHegXGLH5rqUan+M
Kq8dG060pFGjgLBpvtKRk7HmqBu6fE4eAdmjUeN7HlpBWlR1oC1ADDIgCB4XFgl7
E1OfaaxmeR/gptDIkBcJDdJBObHYyO0sT7GwdXyUDbi7qHzbpV9rBy2CRxyU1ASZ
xAzs71ELxYZjZ3t4u37+8qpkJ5+h9/Y8t++MPWWY63a2B+8pVYVxk7gpeQwFJ6mx
x+Fvyb6DnR4iCA+IG5JDbPT9fPgQdSW+yw7FUoUuO0YP1nkAHp8ehBeyFe4NgN4A
7k776M3E5KI4VHs4wJ4QYYDdT4ENcfYfgKH/YXPpeuTqAlqGeKWYH8TDoq+edjeD
7oAy35nqdJv2SDjP9dl2UFJ5d6ev6hJLIDWMSFWXi4hbPW+5WX0B3ATyngPGhTEj
cZM6V9Imsr67dggk+speCUdIPv+N4DdiKXEDQ5rtq7vKUrifNYfCBaRNrgZW3YhV
JCvClQXgBSqBFUSeg+kzL8H5KV8CDvdh+YkX3zTQE71KW/JaAvyylikkWqsHbO93
XRACJVY3yk54yH6E1HJakupalp3ukYR4kOf5JCEst1r1NlkUruTN7jebqRxzHlCX
amYdeFhvoAxZCMVGO0oH0DFqx6UNlyhoZV0+rML4Xpd7IenY7W0bLKCHSdbVdwm6
QY0AxypeQquzBsWEoFAiYDvQrXjZewUBYuvoAe7FKTpcwvTtBTUbAVdVPueGkLNo
R2b/7jH90A8aDjlr3h/z3okHSeMvwbesWH4ZqfTHQbY7RMSXIUsSXQ4czoiQeoqf
exiziq087OgxLLQlreLCtZp1jP36R2rbpmvyRj6Hu8WKXrJCvQPUuGdzvJ6bLScF
MnDKsFMUWPjF6IGNh5Af+KPBm+0rw22pSoGNqEndd+tzV4+lnSF29UqKh/H252AX
djOEBKbnjis9H+rMiw1ayWX1rTOpPh72vvXTsetgjTGkMA4cs+y7zWMIFUayE8CI
3VKNkIclzSX0wQt6yOdAX9q9TwL/bEnypkMroi4w8/wuKjLRQfePpp7l2Ika/1kT
Sq3dvD3Kd12VmxfBIYn/QgSKRWZm1Dzy8oaO27nuZW6LNtaLxaFaETXP9I9GPXaj
A2vgG3Vzv0viUJanSHbM1wDj4Y/F6He1cSkkIB1D5BiMGORLEkG+NpalB2kZZOBj
hsEPOFmzl8a+KwOxSkgMCy7y9pyvHmUUPiQhAamlJ62RXUgEv35iVIvVeodN3F9V
c8Kb4iJ/P4Q4KYdtHwTRsYTIUWMTEbThV6BiTwW7G10HUHy88ok034vwieU7QoDN
iBtIlHgV2HLTPDB66UIF9EDY+ZCwhTQhvjI1vKGVGob9BEUsAgn8sXHgIOW7LqKh
RlpqXUBWNGMjPBgmzD7Mq1CgdjBQgxiQwmMxNRPMMYfy1it9KnHEQD6sPQiqO7A/
MEEDZCqL//MdgiYTaaCUNXgv4SdAo/QdXl5TZi+aHMCo2aVBzgY8acBMpCuc/pWX
Ol0zhazuIQ5nl2uhK7OGjaRpY9+pjics6a+eeqfrgL4V0zHG7tsjB6RlWJMbbhuM
CMro3HSBP3nk/l6ZO1JW5XpWOc7SEkwAbJUyR3Bp0kaOH1GiAIFI1OOXUA5OQ70I
c32FZoIP0eTrLad5bNGbZaS/VAm+/L6zTGtP+OPffXw4zmujtfcO4lIP+Q9E0wZl
RECmSbJ+T0QTTBTkBK9eFpBDBy+R8pS3nSbrUTLHee8IkNmp+aUyc5uUdCUR1qJy
tLRfpj7he5aBltd6ZZDbrJAy3DzlX6iVr+dTulXuvu0CxTFXrUNI7UwUtM+IsCfJ
QjCYAIWT3/LhpbMWNpfjo6ifkkwNL4SmGrHeVHGKHdaxB/AR+sTrPyHWqNqI/eT2
hfPf4Xz3pJyAca2nx4EV8iiPAScf/huO0MFXes3z8+mfss9zibh82fLMHIT1mcEb
K56W4RdTIVQYPtFgZYeq7hwIRBsg9QM5mXV/BGow/wlQqARBRhd0A+KYAi1TLmN5
3vJJq/d4yVnkJ19AV4RBnJYFAlBTN0rqPczTwoMubWZz/O4Vag7ypBkYbdWPABS3
4VG+4wCbrwVDE5o3LqOuS9OGKZ8dMM6m2JiFrqOSqblwbBmr1wW+QZlQmAGi/e5i
/LXEd1pRw9ksd3DwTL/MsYTCzZYmkFjdnEfXnvpICw65pr8kEqp4pEUtEvdQBvDB
ncUIEkMxtcSQsDJoUsG+0exk5wBTdEE2w25QkF83vGjdJ+6X9CIgJn2COzYLiiFu
3RKvPgOjXdMWBkFJEUKKRjw+zyAzQCv0ax0KIGzgGNOK4eSCeuTxS0UEzuiFcZoo
r9hHKGV0GGahf/uxgfvN9B+Do1zKxzH09Fom1G1dqGh6hVuV3RR7WjFnDhk54+3n
SPfgaJMqpM8sN2vTE6pc06y/nNsDFJfEmOJfcJXhnyEzTVFrvJk+8itK8/y38jcT
tfL4UjSP6Z6gZhTgH4uBMKx3dbjY6TxI2eOKYm3wouOwikQZaEk9DfK/VgdRbrho
dOKuV1NUKGnFP1eGlbXgItOWHoCIzYYX9yzgPcGeEWezO8YydNG/fUrACpGQMVsH
UIXV2N8k3eoU0UMtXmvV6QtBZANr4SS7VTHIPVJkIvjHrlO06ZUVtwFLTi1T+Z76
JH89vctBWI0G8ENkZAV/0qHguXic+FEVEzbH7Kzw3LDMxsnJ7Wne2y3a1jr72X8A
niUBCfvRC5+rej8M62Ro05m+7HOOuW9Hy3vBFz5rCP9hUlxKG+7K12Sswir30R0n
RaqKUVvdXY0AryA/XM6AgS75q+5Oyf7ajBKnDv3ETrEKuhZh4r6oUOm7+XJU4Ivl
2iXtOSU5c3jpFXnXP7wt+2iADsGO5MEKeVJv52/Ay7vkvzxMEDHvuYac03MqGkCY
PgfpJukqP+OlyiG7DsvwEkJvKTa1QoFgCA12TvUfbQDPRt9VunNhZsqTFkoIo5vn
SEQv5iM6YUMS69/0bzOfwwsZ5uZ9JkcSEq39HlgYxTjdcglq2Dg6pHSabBpLFQuL
+teGxaMwhk51v8qt9H8almhv7ULUd53xoVoV843L987SKfX5t1lD3wjK0z/H1H1g
R8BevXX6gejspMK1BVfNBCY8j1XbTXcmiYQCRnnufaMt0Xd8h7/McepN4a3cj3fh
Xe/1qqtoWO+Ikyp31NS74yjBlXdDB6Fzh+gI0U284jBYYfvsX2hlU3PXpKR7OI94
8U7bYvOzj5GURJCldjMs1TuaTsU8CizcEYM+Cbra/xC4bKmWvX0gPSHUH5fT5ISn
miBpWiCc5KrjeAPZBV0mZ62a5q4jps9reOcFO+KySwxtcY9NwKlO6kjfxpl9SC2Z
35qj0FnRoAbFUfSQ8umR1lY4c/IqvCDFs2CLccUq1VOoP4vQDPee5NnHxP0lNsr0
Qz9muOOdcAoDTCuhQRWAQeV0oDWG7ApFBSiPmYTXdbrE76lLlotw812BwA4jKpa2
Jb2CVKVskCftTSdqXRYSQGS8RLpwI4hWN9aJE4+K5KoVXKSY75E4KvLKkjYjEiMz
zsocmoisCDNPb9BwsLoHIpNU3M5KNOsdxY4I4wv+MgrYqU2ITvCZDRHG1TltpPLq
WmOiTMcuQDNLaTpFgLVUlvnW9W8jH2LNBK3RU4/Xsc0I2KJP0W0T30sPO8vHBVup
d3LCsJyNSKpSfCyHhmZqFSr63FcHyUbr4w3InqLDupWLDYblzbXloKWYQa3h6hNY
hEAqYHNQwnpjgpnTxEaDiqWKPX9JFrS41TUXi78sZo37oMKG2QxJ/lTDKHDFWR3e
MDuVoUu3xlsykko6MGCeNXzJTpx3uTR6oOtuuEbX/tl4PJc+87zblTaE0Fo5MQt8
5493g8r3TXxl1cTKuXNRyL3yBO8ZSKOw3jEw0XDJulJ1h2/XFkHbKjgozUO9WgVq
giA9Ui57Q5hkoJMPKikarpOFVuIiE1/+X8f4WUvAktWG64eT5Ah5OCX9YPYV/BA8
4CLlKWzRQTOImzPnMagBp5EVJ9tZqPDLmhxrDMHzC5IJehheAlgNnIBDwCeDZFN6
id69EyzX3hO7y6FctiZWh8gQsAuxmNdx9aHflJ4pM8Imd/hUWbyuPk71Vtle7s9Q
5IJ8tdbB7oPae19L3Z6P7bRcK6h4W5Mvty79Dzwja/RcV6SaexqMXq94gkmzOUP8
OKno4LKhoysGKHgTCaaKWPFfcCP25D62c2yMHQhyvCFFo889pANKHrzFh26tai0g
7jf3KZRjMAkenGo1+4N0Sklz1US7ole2b6eGHXoatbdBMGt2ood9r1dSKZrtPUdr
l10OWdgh1R8lGk72gdhtj/xFT81AqwL1D8ZDznNocFPQeykPPcZN3QBioI4DXkXl
+PgKnRYjyaJxM2ldsYOGaNFoU0Qm/zT4Oor8tbnewOehwCDOIt5+mRj9xHaQVPhP
K5JrV5vI1k1v49QMFfzNl770yzeZ0LwQb9ooFw5CxSJIKeFPQd89subxlIG/fVdc
ikGg475f3vZX5GUEfF0eDmm497QEzYX44NtTcHUqveTVH4ELsTx+f+/JN+ghlUKq
ifGhWtQuTKfxJhd2XLcl4edz9O1nsZDI9QxapMDVX92QXr7Fb2H1rlXwm63ZqkHB
6qRUt67NngWlMial4T6OthagP5Be65gRWkFAi0I03dIwasH9pKQ7E57ispSIni7W
PW8GVZxOakBA7FxEpZ2+rVdMuYDp7JRc6Ob/r2BEv2UZS+OP9Vzow9pVTgJN3vX0
Ya7YdEqj2Ay9q1Vnwhy6dDowM60QrpQAUJ+NpbZyILP+75TLM2H+Kp/u90Ea2VZF
F7dXkY1Fu20isWcmc8vS59SHX1HytgNX8yaVlPE5v+WIQsBugcqtP7hUIQC+Tphj
WAKeDqd31DpxXdpth643W/D3Tie6wmrKZLMZ0WEfYKfxSQm0EjhyzJ1IftXYk6nh
hL2cVZN65+UDAkASyMAfmT4Ztfiyo7VUxhlKL8RGZy0s+N5ccs7YTOJh9vGFkIha
RXkAntgVTngRZrYkSj+N/SIpJnBzsD9/JD3ekHj80kORKbFGcwZlyssmfW1VqZWT
o8uXqQvSVO4vLHLnkCZx0//Bovf25FW9mKnB/mlB75+sIiOlXFZvHYaHILkwFeFw
cmOIUXjtmMPVO41l1/feXjPHbwGlzh4WaQUnC+hBudN4yMB3Qujjh21QWIMWKky2
GAg7cfPjipypDvBbdSgABWyesS7DCpPEhqb/rO7ulj2XaxAQ0xEEnO7+FAEB2HcY
Kgew6XKDmXQe4BbNjwcQYzKkutjonaWiXGa696+VG5j89XQPvzd+rlrhnxxWMdaj
RYhk/Y5sIDrAdY/7C6CfX8fL+N22uql5VeXVTVUde7NKJQlQ1Otxnsvs1KQTsXUY
d0kQw1ePmlt1goNGCfYKJkxDxW5bd35uXqJnreEXdWRHxAczovhwdiCr2LG/i2Gm
Rfbsbp33DkM32x+eytzB2IW3HxdHVB8HbCw4spgKucsTmCWsWQYgYYJ5bmdrcv7q
WF0eCthrc3Q9fIbaAj3Bo4qcInM92sL/GLvzY92GOUoOAazmOH1iwmAXu7AHj8UO
aZ2lAwWAu4PSlwq5GM13xNRY4oPOUzs1IyyjMAHORJDhRORm2kVbeUh7YroSte+j
3yJdjswdXB1VQVSDRMCI05Vt8I7JFP4xpfxoGAEh6XrsKEOWC4T7Drsh0GLKusJL
fTUzWqeozmv0nla+ayL4T05wPPKKvjJfSWCXB7Xqmtaegpy6Sp6Pn0PVx6Q2yzTC
/qw6YWKmYWEcDE0fPZRtm+DkgRDJi4x0Ata1x9NboEZU+cJLORUubpN28wb/TJ1X
69BKuR4GK94o74KT46AUck0dexQd23oSXq6IwekALx7zUNDySr7EmNWTc44d8wpB
AEBlCif8BCy6fRVTMIBfTJGIzerrFd3GIUP2Htnn35rkL4WA0l3EMvl+KdnraOuc
rz5gkdwwYV72ZciyvRkdrwvxU7td5J8lbBDPa4BD60wQ82nv8HmWQ77/7l69N3WB
jBOjmtqh+iYGq1p8ZkwMUaZU67cAEX1WYh925nyeUXYN2MEM4QmqJcl+AsirMTRa
lne0tM1hJGoMfr1F1/eHe69OiB+I9zEb4tYbiU8r2oKa0k00wmYnf/gQ2L+VEZEP
J3yoc5KFxbwxf584BwLR19idTyy0SwfDyfvlo9QOyPOsSZRUoc6s6JqOfSMDU9K2
HQWG1m4bBZWnzI0yWYhWQkaXLQlqzefi0Mk9Hx/s2F4G0ppmp/K0CnKfQiMEzXqi
jcj09mA6KautohXZpxVvhwBoh5aR1mavC9hpUyly3abglU57CT08R18BWXoq5GzA
0v3jA/4S0Y5RAt4mqg3JwJTaKzEgnu0fbKEKK5n9vxl5HpYRZB6yTh42tDLWU4+y
qlBKNzuPNURxC2cGka0xcdbSdXjNPF9fv/6YQDmyoiF0vm4RjXVaZGGpPAY+oV7Z
uPrddAQJfIFoW/jA+oE4mOOPsYr1AngE4vxKiBTwPoLEjEgbNbwvQhnhBM0ot3Qy
dn1UG/qku8drxbUcdN5Ntn8aUMeEJiJct1MPj/S6RcGGcv1bgc3fZn44FRoD+wXS
lQ4FLgAXRWAPzOqCFRoHNeyJ48g1FtO4jKKVcoSQSii+kPYBHlX0mdInfwByiKnN
4QTXKX0V2B9heZxDHultLFwwnTC86+wNYy6VX30Dq31MMGaardFD4M71/mTXUP84
dsgRVtwwD9WqYSjCvfgVcNSzvnZOcZgMQwKTb+S4zheW4mDS5Wqf0K57DRLp2PhD
UctVrR5MOL22eEbdBTONRQvnYajUMKVURqHG8ZN2IpKXPbTtYllxZXBbviEwrHn/
wp0uvBo0Wv2ZPHhk/aX3TK2vMzS+BohB53CGbOd4YGPsJXFNOsi7mgJXdpX+Ut4K
aWn8cqssZghzU2+ZMTmOJuSycpqUuvPLqNeTrQqMcybMrfBi7FUEdnHWxkAey+7w
1BWIbpHmj+lraCF9EkanSFg4Ohgd8pjz3ATGj/2X1wUvsyuXKWBsC1amVUMtJYRO
+OU8h9z0euc6pREctzAaL+y81lHQ7Oyoja34vxHxEjexWbA+iLYO5BcE9o64C/dy
sysA1i5i1cD4cM1AT37rQIR8v+EGgJRkz556kyEiJdaQk7EyoCR+6Xdhm0HWuVZO
cexHVhBNUPMWMbkJYGdSlm6C2U+B7N5j+z8qkA3dEJmjlB91wKERJTwOgbfeGvjf
RR0jbyn9PXxy+W1KId3DMF9SCypktc9iUWNN//qYisT1aOQBpO6EFMW1efcqv0oG
Hw+36fMRaPc6lAX0r8v8fVskCfuFBSMBxERCZyCs+NC5PQPJ26xGtKCOkeCyf67U
I4bS5KG4vPLOfFzTbAmwTxOP4Y48Wfs+WbIC2GjB9fafG1julOJ7mkX/ePiDxKAs
ZlW1CRFf14RIRTZUiGm7oRXH3JlwtcwyX7SN6M4PmnV8hdMqKgJXRcMzZVEj1woK
f5rJYIWUu6p53yP4/kpTtWrgzgnVBmtE7W7vFPgacwJjDCvBH3pwq6Mj2bxJghU+
3DChcdMdrbk00AOq6BOnwuwaDCM4AS73l8hyOO1eeu7c6nqC0ldkwsJ3pLwnzj6c
RXyledOYdYftAC+lJUa5rcaMfh7kiKmbAHkWnI1+8NSxWCXNqCXl1vpJOdUnZjfk
2YKvkxPtllGsZdeIeI8j+avfiHTI08Im3dngRnwuZnIh4//4i1hUFLV1UVJ9Xo7h
dhYQH3L6DMoR5YVH26tn4Pb08VjWJ1MKUhT5Mf7q7KLcrBD+lst6TpW6g/EURiN9
pT7+Mv1K0gR3t66rsH0FYBMFOlcPt5gMZEhNRdFQ5eGVHZ3/GH1iIqX+x+5bD8iw
sRkMw8ai6SSGwq6LqpM0A1KvABHwvAYtW+3uHQb0+OHTkPXcqKayFlt6dUQ5Ptl5
vf1AudiSYDNG+xePc39UnGIA6uF56feBaZRQNNmaGOsqrXLBX73CK5TEuYy4vUWC
7U7DJ5NxDKZb3UGsR+eFUgjhRGxcs8QwZ3zGUA1LkzS1jirahoVCCVKW+5GZEpOL
u0XZxcaNVpR7lDHmzDtmoj7/NQ7R4rAqHDS3yIYdEAD1zFbiP9XoKrzhhl2rULXG
PjegaW1Lc05VS7TGQxaPkPUwCNYBiYD8oY4Wl1WGqK/qRgvYIuycjgxonhsitBlU
3PwI+ZlNi/ellZcp3Os+XgneCOsXvHir7PUWgr2AJccrOAH6CehNpXVZy12UGq/g
N2YK4XCl6f/Z1iZChAK5SqzhrANqDt5c5gu1vEk+b8dy1q33sngne+HfUcuIvYPB
s6SXeu1Xqomn/YdOypHMfERrTh9XSvAcAY2z/pT27uLl+wkqrKnU0URTb+roZ7zu
FntZl5r+0/+4vs7661mLA2+xsct8NHo8xRcEDHI+eFjb5TkJMKThI74VhNC6kzVF
GXLspeZxDyvIZXSK7EaIc+oR5cjhPfZA7XJ7/VqVHpQN1si8nKQ2TV2v4yq3tLFZ
dHaRq9JdBbeFWfuIxqwXWfYl+wFKonjaSnTeyL1FsrLIf/j6bbWa2KFe5CdtWEp/
+gBSemHCHnj0CQ99+yIxfDaVvCKJOT/PxuSukb1f/BdFnxr65XRbPpwqIo0lmIYT
AsIS6onyhNmR6FnJ91/Go8APygNpIU9Z22gWJ+ZZAkOhWc4OSfj5DvK39ubH3/S/
0tG76sHAhpZrIFk8wtd/5fZmmjL79iACw7ddReJgIQYZZjMXANtzjP3iriaZG3Jw
+wMUnDpOkz0FU2dk/WS1Me4+b85FdUVIns1X+HvC2Kz95OfZUyoyUc73u9l9AXa6
Wcpyn+QZ+A+yzq/oA+zLn3yUX9plBBNCDhZL/KhVsTk1UFA/ikCeAxOCBy/dquyZ
XFqz+gzy2ffrOJ2BkvEDKz6aUEQHkHSssmezig30nDHDzqoW54aeYhTGoBEvoH8x
uTOfMxIc+X46ohKtZGbvp1ZKmDZVCPOk/YNAbkpXzFEbnjeVs0amUB/YIzfbfN4e
Ugh7TfulT+A07SiaQ4rdq5uX2pryV61MaNcVAmDNtE2CVqc6gzuAvCpy2YkzCJnM
B6VfJqy7ejAgy0j55AjQd4dQJpE/OU0S7p3yRDxtSGwlY9v87G5bVclJ8lbDzGaH
vGmleGQS8abc21IGOYSWDO5IxvsI36iwWlfCVmRj1UQ4+IyRDMa2paEDGQRESS1m
xI7ma67i7O98fBzAsQ0iBorPf1YbL2axHWJys6ufImdiSTWag4DjrpseBWiqChD0
kUIv2/FRomjmmJBdm+0EH8wrYSCmbGZU6sAm3Qudl+6CEdBDVvhstPhiFYjXPOtG
SqXtMPBcFfCtzn/RzGg42KKsGSn5lIPgHLqIXD0eQMywqyaTtyGeHC92jHz0qjyr
SxN3i5Gm4CDHwJ+oVeoHrqObf0ZpPjXG71TejxHb1sKbCXBIv8LVQp9x1U1xd9DL
T8Y9Tx6ROy1QG/MhZOcfble2W2xXvIZZKcIuG1scfv6MxQbfCGIcR2tn7qS3KkvC
DkbljFVXVbcbBwfAAS8lkdi/eKczp750PqASzDfnuHKGc+dK+St3S/Fx//MWbi04
0L4WVooAfMdu+c5NjQHArdJzVAQkRewufFjL5NOvpo1ynYofokoGD7SqTIXSEFCe
P1WEvTTSle1f89WqBGkjOuti1vMekQlr1uFJfNsyLS08J+Ukb7i59MnHM/hD7GlK
h8cxxE5NnxvUUtFuRpeFaSY+DT3NSKPN5ybA9HHV8CdNUtVhjPStVopPygYqanxj
+ywxC9VbdKynUGOYiepInAL20oWNAlVi4UkL083j4otYEPlS0Mhc/Dd9a0/6l394
1DMZ/mF0BP8dDGkVf5+jGr0LlTdm95kmBOkW6yFvME8mXwZucHNYcxhL5pa8gljh
Tx8eCFlr2e0df59pI3DRXS37mMzCMQffSysv8xAQqh79o8WveE5ms+1P2UaKljmO
CUfmUyC5pVW7iyuCpdQqa99YSipi3H/n0jKVrOEtkQ//NXhtIW5Ja1WnE7hrwLSy
Od6eZujqygemoE8G45CkKwmPuR5mgJAR97zKBf/1CKmWDC5gCqNtUbfTdX/bL9N8
Iop8VjlcFaqmp7U+Z0uRJLKq+Q6OBJMkLxNWHWiAXt6mfN3a5SMRYycj3djxX7vW
ER9vTIMAyk+ZhLM7IBAc96aFnnoV66NQWsqWXk3iDZRGcwqQmOb4gVFdX5Agx9zs
NHGHo2UNWkRz66FA76y8OcWjKHPLxsAKN8CZZoWG6YAzZUfPjM8jsVAYJJTnaaVa
NFLS5gzYZRcUSqY6q2ZDa0lVTG1MayV+bplp95e9K9p2HDXOPov5FSYPYAIQmqzZ
tdTQryxn0yG545NwethijoiBesmgN91oMS3m6qVsr8zd+OjdnOKc8DsFZoo73PSN
+Mr+7ffQl1r8Ns04QFK24j30NlQ1x2Z/jzrsdWtp8UB+KurKQja4NjUQDl9UTyeh
k3saVZd//Lzn00aXQvuMSAKz2tl/O87TuBZqBJEOJ5mNx0uqivnzH5BhCBk3jYlP
8PEYHP/6sHs97/QXU8aY9sAq3HNJNbWOJZjGtqYICoP2nfCKZTDExUcH6d6TmVLs
2RHS1e4O4mWfKkPoKwi+kHB84FEsVCpavpVABoh3ZKeIOjN3cF9NQ2FYGPec5FiE
/Vi/sIcxRxh0fVOi4mm9DEKqGemVxrD/KBnY8vVq0/8NJ9iZrJrPAjynzuKzljs/
z5wO9/YetlABYqxnKlUT2Zqo4FJoUaDQTMKs2xxNPXfMjhC8NCUOgxrjFakSCUp2
g4NTB2uuMno6b3Ip7PASC8YuueN4sY48x0k0yDQjllG21FBYLN1C6cX2rqNwEz+r
E0W4tiklcY30YWHRe/aw/NDdJueRHs4+EF2Yv/QGbIahewmDLHzWK0k+6OgJNrbY
WMtn7hMR28sW1oTQLfHN6yh0IrEMwie0PE94G602UBx9cpKcXH0wLD+R/lBnihAO
rymlEZJJfOjW3qe6PKVxlN0l18HB9FH1IHbASfs57LrvBFIAspOQHJi+eu7/mmYN
HMRCYlxTAbCT4pN/PWgnOG/aPOX5c9swjjsVuCaaTAAG7zl7bkz8KjcG66ae34wP
Sd10F2bbziSEETDFrTw2g6O8ZQCuee0xfPw4vKRshjzPrh3aEsCavG08ZOfXjwaV
JWoONrp5DCGIvixSzJqQ3k/stdUP57azbrEQJAaRMQ3Oy5Zp8E6duKbjqwnwS8ct
G+ixTUqr/zc1kxuPMOtxQRLrdxcrutrftmcVU3qL87L6GW+1R0zZSne2io0SP5U7
l2wbSWFReZSN7QTmcBgFHwqTFE7Ib7qFUvMH6/e4vZvN+r+VzKYUnxKkKUemvcKK
NczFVRkUkANqMlgKuRnEE8IetrHJwqmWbqfKoGPAfq6Kwp2Oe2JZ5CxnQ5Q5ghMa
6aM41KqXPX8wffzZl9M2MPmt6tnGheg1X6+OfITKLexMaTV54Ll49KJs3YaQyneO
z2LlH2Y4RXuUB/dO4ylXBwrQda6v1jP0IR5sIhCvo1zeZBJRfX3xiwxYOwzrEq6X
IryvY0UwKawCmZJVtvRHflC+1dz+4yGLLpaBkaUYGpatOjxiyFz2waR3qiG73Asc
E2cWPHEGtaZVJTjQMboy/50VqP67GK5A7W8PjzCjoR9xsaQBkDGx+kvSrOpwNhy8
WJcsVO1pcC8/SiimfMJZeGVQ74eKeBMN4chOuFaZfhtTWC5RdfoYZxgcML8vaVnS
gH9caUdWk9v6ILupijBPx73v4xaT86ODH27HfpmWwut6F9TzwI0UVbx1iFd2fnGJ
FuSctp9W4ymzFswVGCaVtxC0YnwYHNzCDNTCI03gGsI/b6Wlk1tY2BSAKTCyHn+O
5RmMIduUAs2ZxSY81uGfOFO9C1i1D/sBG9OsMRbxhXUBpObph/4uVvsGVtc+bz4Q
oQq9Je7Yf/hG8Ip2LO0ZKpdVGuHunRGE3zpn8AWDZSmIMShKckEBIj0j8pECHwVH
y5tIrN4/l5x/aNmPyTeThoZnHuBZRQd/2j/CAwVJavkBoImvl/+qh/GJ9NW1B348
y+e+n6ogmvB/dnlqYUARzIN41u1IIygO8ZkC2HnO+vzD1Ii+FuknxdWL0Cbcv3hW
pf2OGyriZmqvRQCf+f54+G+A+O8zODgPpcebZG1kZ961RSapiBUdRApyoVLvQdtW
SRrgUp+7s/7chc7kxgTamHKwCmUNzmAUlZDIWacyVwU5NSFNh1NC72Dib1YhiUq4
szhuM3CKMh4O9IbMuetKatFTyFqSSpgW7p9BKKMkTcnT/c/IwisdzvpX8hXjygZ1
vYA1IQerae3DRSpN9CXZ1TooGNHTGm6RkVcIw1khtzQPI4eL9JKJloM4JUFtGotd
1ARDxnlersBsDVIWkDBMAQ2/EGvhb5M6gIhE9sg1IUtXS4+x9PFuCHOTN4Qg/kbG
UMSjcxbF5UAdiw895ARd0Q0qj6azu4MRCBxvcF9lgL/Nyc1/F8V9HRQugS/t1FJT
JL0FZAmATdJV327W4Euqy1XrmNb0xrna5p75SHaeRUrHFaglLV+fyz/Xz/qrdQXn
FudgWDhdl7UVyuchvZVfsURwCc/X+JYnXMNNT7DObJGrdqmhHcTFD2x5bH2+XkIt
ygIKJebkw3quq/xrbkGddAHSfJUAItw4T8sO7/mfkeu2C/g8tbotpr/lt28yg2OU
T80SplXqU1E08lhRMioDHvkXfLgQp+MX/j0j4i1cLN2j5PfHnzjSTWoeHaZehE+L
i7WD+8ddGM/ZmeZdwy14J89XssEtzVpyaUl7m0OfQCgXI5nw3hbmdiFobBPDBHe4
bJLG6c6Nn2548wX+ENZOKY4wz2NTtf3LsnZrwsxG/ZQaeKlSvN+B8ukuQADMeTp6
QIWYtYohLkwTtQz+c5NEiNth4DtLJjNCtDKGB+BbOlZlxwf5cGR5NxalBOCm1j+K
lxlTptwWU1j+I266IraLCAZfpDXwstsnN8q0mFtZEApSV4pUswfxTUCr1RietenF
x5Hjh77tJTIEE3sbqyzygVYru7Om7rHjykdsfmbrQzrCWCtUCbkGzw3MVCHWvF4+
6s3L+n0miyICwguHTp9N0ZR+J+c39tqNJE3b5IxN2egaX159UWskjWFW05uToxKa
iQcgDXY7KZjZ1Yu45xFYRGeTOvnxBTGxgj9VqREqmoaP57O8KYiRFRigVshyTTxQ
OTUwUA5zAUelzIx60/laFrag9vn/uvj6jR/W5unB7PDIMs3Cqo2xxLRq7PDDcOZi
hUTrvUR/MWQVEzRfeWX5DS7xml896Vpdd87XXC2x7gNxGJotsI2H2kFeI+95+lpC
9M21QhFO5e3SOX2C2dnc1+ZlAqk4eU3aVRmbs6sr+oADKBDp6M+71m1lwJKLMpO2
NlJrokZ+taKjJR5Thfuu6OVGXNPgUG+PEjFrDkVNW+aMZCNpPKy2AX89mAHLCy3Q
ZcXq4F30WgURs7EtQYlFYsLb+3BizSv4GZMHN3gOmZObK98aIoxi3Witlm9oF+4W
GarlXVLBsQMMsH8s1tmSJyELMlpxs00svsASOioWKOBVBsYUlpKTLC37EOPtJPJA
EIJ1Jc8XDAzPdbcLrsjNI7Qz113qjdwniRNS4HIDJHfnrMTY6a1K2bVsg3t84CXq
5ex9r+7gW4Xd2zWWzHbl702tDTaYIe15UOurDJf+CcqLec5mX9KEmA6ZafE1zncm
SGknG22vcUH2TLekI2XUJpvhjO3v70C/wMey14VjkrFjbkm42tJa/yY9Gnc4gfQc
Lc3mkV5tsH4JaboLcUGl4/Jdd6UUGQBGR4xIA/14Na2XEbap+e7lTndXkWImlmlV
0RZ7/mQn5UvqC2bIJ8fGRexnpSmbEpjkyX5VTfftHIy97OKEMAYb67/ij/XE5JO5
4Vmo7xhCCLJWvWBaHNX7capdOHvtbRV9dPWmckAT5uYXU9XhCleLJvDzLH5toYDt
SqY6EVQI9L9QMSojcVRNryNX4s7IsPueTG9OgmFHQRC514VQmT7JuOel8qMTPMlT
JviASELg46+oicY0HQRKd9b/qFPu6rVjjeDTuVOLc51QUTxM+wyQE3YWIhICSlYV
y3POg7mOwqe3jNvs9Utcnd4Qds57d56J/A9wpTN1u60Erh1SVXdrr4do494DrG4c
TYlhFgktHlToCFTZPOl4SOK9utNP4trhWHgZF7mTGIWaPNQHAczWtwgamyby8PlP
zX9HaAJatqdqTKnOD3velg9ZMLQ6FrKaSbwRtqpo8fIXz5S4xdyHPpN1len/EDzA
MLETYFbdtCQMU310XSTfOQ+9ngyIellkvkVLmUmQk8xe3g94YnbBlNOQyDPkzsb7
NCYrL0CKI5KzTaa7spa27cP1v/uRL4JRO+c8jZzP3z+DxzomDGpFcWPULGbMjQ1z
FzzfOgn1348xHFDMV2dfQtBF5T2wWUHCmExnO2lfQk/tLUCRlt6HXSBNvd4M1Hjr
CGFTbIR51IrAlk+LxthKf9JaK5GCYcYTtrQfc28rRxl6V6Nc/b7yChQLix2Xq78O
rCSeWVZDnHdjJUvB5yHDpPA37gFNhpJeavLK4zkgMsLhRa2IpREVM2s7Al8if1Zd
eaFZgmcYvXN7oNY5tDTEIy7PrdIu4RDSyas5eJi+Gpy8UOMkWT1Ct/r3rnIa2r1R
5UqPhHGud4ZnDWxQxFB/JEkXelMn5kzs6RZDqFzRhznixQlA74RSqWlP45qS59WT
g790LX+iHoKYR72tlA7XCVYryeAe/RpfXPNUPw+Yl3Dio769m9ieZVZ/+SdXIyiH
NKDtio1c336Y2Y2PsK1LZ4moadk/n5NOXaw1rSU5yzlriSHlSR1srBRd2xmS5Qca
tDhFO1F9C8w9rdCcHX08I9N4NkTWHCfSPCJhD8rx9guE0bFFeL9FyOfFsX4aU+OE
z0vAYOSeBddKVKFaor/I0rD/0i3IH2fLdoGUUGsKdl17Oi65MPcG1Tm4R1irXFed
yoAQpyNVrcN/dDU9pyTVQr+De3i/1OHyYYHcfJXdPct6b+9mTmxzixi45+z9ita6
zxqdYgxnzjXXVaw3GsnyhyNYJXmCzz6F3tvaEBYTOJZ6h93O7MFVd0L98BEcWpao
ULKh/KJ+wfpL9+eVMzUaGsLXxUf4CKx3xrHfYkDWGC6UCuo7Mn8JYnIOIVZ6teEG
o9IFGukrUI6BbtHFR6tW5igtawSJsldMF+tl4nwuVcked1imZXOsnulPvDrdd4h7
nQTEP3na9gcbeo5lQ/FfEw9ofVg0zuo/x/fNEiiUgJnjQITGdwCufT09xKJcGgsh
go7cJiOCdhcEAP9JlvvLOZDrNh0/ZWEVj27mhps4coqAvc3g/2i0DBSQqsxSMVIZ
Hy0uuILLXZbpSBhpm5GuN2tSodOJVXDfBGeEu1WUftPooXt3Esey70TPyp2Q7WPn
YBNRUCrOPOTi9OgAgsaLGkPBeN12rb3XxmToliE/3wOFJvUpWVq7JuepRL4ENfCG
C4dL17tyePeaAleyW49ZDQgtEosV7qbRJ9pMqJhpc6qmRI1HwKhJm6sM9EGM9BN9
aLDa/T4e+ZMnztaFJXSaA/DQaxz03zuHaTEG8u61iQtmnu0rL0y/lQuEj89NxANZ
rzdG6qMfXlDB/oVDPG14nKW8Ts0IrrS1uIKmvLFGFcS+bJwA2+yz7u3OrPlNFI7i
aDkpxqst8dXnhL7E+uD2zY3JWFjrXQT9Mi9v9cZHM2JjQg7CEqZ4T0aCCjPx3K5E
R+wv75pd32tf1F7ApcQ/CExlhMw0EZHoTXemArT8P89dUDItmjmbQgcj88j/AR6D
wazm3e2NYZNq/hc3TaXTqrcpPefHYzMJpyQtD4AHoHwm2Gaf9QKOVGzUmK4mtLO9
dwweit1OtaBYAICVlkBdaWNXRnI44Uppaj7Iq7Gz/WYMLH+PslDLWpii72kCEtB7
fuFqAqzuOCZCdj8uE1T6gEIdsP+fU9QOZEUIm+TtNeoY81GjP9/bamiN5dtKXxQ1
8YeZeS/FtO6PNBEcKgkmJTVjxc6ppkBmdrXXtNduktxYIIRLXkXVkxs2mwlmdxCv
5cdGoBkj2MpqSCr/Kv8xjKAN3opLsTWFwJpcNhmIDpDY0atiiM1wYoDRmvGKEIQj
CiwZPSlcAq4D0ypqNaUSBgtz5a5q5RvPGLVBbvimCW/36n4sG3XyE7TIgwtEbpdF
5/fafvLeumcPvkWMVHFbHStMz5342Ob3LGRPVmzp37qIQ5FRCs86p7OGR5FsXCh1
GuR3/D0jGFFsSgURMf+vj3XAVSXDvpKUeacegjXrF1Lk/HJO7kLBHOnvoxv8XUbu
VYcjoOosD/bgZvCVhKG9AC3xxzsob7ERE2azM73ikPBwERwUWZI1EZJ0dNbOc/ue
aULBU1n7eiXCmYZGolF9MTEcgAQLBgCIVMFL3oBQmcHMf0hICHtUCCZ9UswKd2Gc
T8a1wjszOQjXJw4BfOD/ttynvnqT06sch0JCe6TTQ2uv65iJ+cPr31xQESish5PE
sti75l2m8b0W9mePbEBjwhXsOqOV5bej5goiFj2YA88hHIubJIGTeddbvuksrvYN
I2Lo+8Gazw9J4eCHgOuoz/sCwN47IcMbFljYCB2ArigwaIB6wss5cnw0K41nNNPk
wKi+gGdjNVWZX8AUOOIninzmUk8BoAD6mQ5K3L/CU2f2SnqdyoLz9Lr59FV+t+M+
Z+UTPSW4HQtB0xLHNto3PKWo2oXUBsGu2+B6vEtjOVy532Plwhlx/9bqCk841gbX
PH+lXi8BFz3KVZWb7dH1CQjrgcN3iQRe5+9aOVgYanW8fugAPQkymCOixW9hDeq/
rGSd6cFaLriXm09IGGmcr4ksEpnzLXmCPrP4c8+6pes+Z9FpfUOFWvLordhhpPm3
Xe+TCXqbNA/VWWbKcNlGDSAGoE/tAM3YlzT5nLO4PXfu4WWKzKAhUADxh1Nnmvlj
7v0F4eMhp4uQK2nwuUsr5ZgCWrBpuCJfd91nm9WKGPU/kJFoDRJe1gfZdaF5WfXX
omD7rRm9FyVcMEyADDAQewQLwy/CTLJhYbD5eNFuQ9UJszTEdqxpPHW1uJLVfoWM
s0g8xZCjgdgs1EYWBG4cfx8U+XyD2Ka3N0ZT5uu6ysydP5XV2TolxI3GK7ZEspsW
CneufdShoOkw5f4MLiqLu4YnL18mHkiS+leWP9BJk3XD6cNKGSyN3WH+JnGGw+nZ
OX6DIGtmMPsxuC3l5THlRFmgSW4dKjJ2lHX2S9i2Bbuw9/S1o4T/D7MrDG8dBBl/
4T4WufZqOXZzTqA6tTLWBB2HyrAR6EdgjBE2ky0dXYexa7mx4hDC6/EAlBOPGOtR
eBYF/HkucnDlw6RZbGbfbEHQTT9K9mAVnEKu4IZ8ox9MRIZNp/SqtAev24w3IBhJ
h9ztHvX+/7PrIaoZL+ljz76th1cZGCHOf9HkqY8VB2w+GfsVkOzmrIlR2wJ68n7K
BRL1SU/n7h5HQ5+Tv+rCQJSwQt1NOrirsyomraHO7vLL9WEHiVsRlserXmqpO3ZB
Oa09cABmjKR2gqCTJTsPiS4pljqpyaO9IzfdwYOX8L6n0S+SBQiIwRjy5Icie/jV
Qq8qgyz2O+dLzFRPniek3YdM8rwsQdFoB/3JsEGKDQQvFOXSuhV10ktYzChrFZPh
p5a2AYRv+Uq9UPwIcSwYRrrZJmjVBJ8MaUB3gn/MkCvlIUmm45TlLBMa5BUTe0Oh
lCjTT74cTQST3G1D496q473uIsU8PFvFauMdRYyw8z5pv8iwrxVdvuN3Bgm5Przs
SagLoOrLvQDrwRQ12YiqVYYnSvRbdLGEQrCEVRkJqMQuq4AFjfwxTCqto/1Tq6cP
nhejEhr8JwxwNmbGIrZhE8u6dTNKOhpxZZ6rZNk3v/j6sHBmPv+/iK1oQxJpqc59
0Y7/K8pZ8NfbEBG2RpDxDFa37EY/NjdrwON5r17CdR/S6txkFE1oAPgzP3tSOmfq
qMq+kXtu8c81oMvB+0e1ZPW5ovYqPuIdCgePCt5nSsznRiDRlXjKL4MpZig7kFXP
scflVrii5SpMdevigL+skhmcGECDFHbE5rocdivI9Ift8aPf/myvYcOH5hs2SDcF
u49pwXd/jo57SioynFXYh4EkCKwwqbgVaBor54Rv4kKTCbMXkAMnxzQr+sXwIoHv
IRJ6y03k/vhbtpv7MjE38SY2EBuQGIck/A47ha+1Tia9xlN7osddFWhb5EgOmCPw
LtH0h5Si7TLkt+/e7I+ovEId71ihyEvnJ79QsRAiPL1nbsYqwHlAiKD7MQ2NNAvi
2USShKTkUM0quNAYlYZid1+PGkbh7h5ZdZxZfSxwBwCbGixNEyN1T6fZBNIolJyR
GRxuk0HTIXXQkuVB1Orc3H7FvCrDuvWpVvpfUEa329XtU8MG4kQn21rTkBV4butf
qODuVt74WNVjgtlBnxfIibGB4H4BiYhsvg2tVXKyVdkGxkJvOohlBSEoIfVemZJ6
dJeocUw/kiVRnnefYKb/fhFAfS5EEmRGSWxdooUXQtTAq2tuwesWMSOWIofTYGQc
Lbml4tx8ooDm1oxSwa/dvMmRQUaiydVePbUI8acna2nuTcxfCib/sdigQiLHg53F
N4bDLx5gVZclj+1/kbLpBeWgNiidAAtQcTcV91IeDy9LoKqeaQtQvz4IFL4+sXfs
9+x+Azqq2LbiCohHw750y48TTklnDTJH4pvhYCJKyx1oNlBghZaZXwWH5cIhCyEd
8GdFBsEWpsq5X0J1Q8RwLT5u4Uh2hG5GKJRY6jvV4oYLiaSc7lKiIRw2/SB6Fdwt
lack6GAglzX69YNhOeZzQkCZaYPtnJx31ayD57nytxuQhxnqrUibimf2Gp/KQoLc
gIvzNZ95Av59jRLuzIDQN7KUr2lqsKqjSZLWOR3MHAcsvhWm8McSgIah1kcQ+sVv
bwEkuw3e9UqrYpXbV3QvvVLdojoEBL6gwZxeUJw0LPziff+NPPlVI3k3zzVFaGmO
NJdCUF5/7nQjkn1EDWppa1lPVFI+reMC/Glu1lVY87mr+bgRwhZcAjRBKQUjAcRd
ZoeX5mdA/0SNXmBY3zodnRi4rQ9Kr+/hQWvrNGzo1cQ05WM7cNYpKzPt7dedYDO1
zGcnVbk1lEfBQtZoNTUz5ZCpoPWCG7atuU+AFKIPSg5bdXNTtwlB/1TLEEp+32Yx
d4x1IHTUYJZ7fpOFSFzQ7lJaVP0zGQ+jBN4J3vTpWF6/gyjGeDLDadvpp3rPOKar
605gX+tNt6hvco7G1B3Y/bXWRwn5e6/Qiq6paRZkktuImYZC6ZlLu+LhpzqY7a3O
IW2JRUJnLLKTgH5qCjkYyTMaaUBgg+lYEPAbHDC/BwUcz+1Atz0cZVAT++VPi+Hn
yXflzrsV9dWHgPIbYbstLei4Mrhj2pZWXq7Hsb73UO97GRl15S6mOisPO9mTvqBf
AMX5Aths2RU18CEXRcDdOJUdwcPETsRsbZT2CxAYD9vasRr0RmFL00CQ13YMF4Dy
Xmie3giTZ/Cfmq/TAjFYl8iauQiL4UFkNeCHSyOU7M4tSgcY8xIjxWPhzV39TMWn
ytdem4p82cmbgMTs2fX6w/E+16UshYvM4HXcXLkY3h5DdTP8dDwZ06mNk17eKUgg
i+zaRr2wUQKY6URDYB+r7IdVl/fnxEpzeAjCDWLBbfrCekXHYWiEUQ9T98cxh8l7
uOe6ZWeWh6vUBnwmFShS0Qw0E7tejCRji5nzhhk1oR5xX00UXpVZjk/CLfHpIBE5
H4qYcYjhg4Vj4D/XoMOhGFbR6NIz5AqkTkavQBcDAqdR/IX41akmsDw/1Luw5fvU
75wZgPXCoONDKt/07JTBzEp9fdFjeuvuOSir3+XbrJCM8SFt1BrmWmEzZ6XSNthJ
ap0Lgc4IWlS50l4fk/7w/6MLTcY7bXFeIaCFPN4aMOlPQ/QZ5hRRSQYwKFRBoyqS
g0V9G1kTefho4z09IEYLT84tSCYxmbxZlkYdxWXK6znIW20Cp2Zjme7oDTX6Ej7r
8qjZMwkic7wDW0QAXmHxtdxALG2pRlhvX5yBQKtbX1j3nHouK9MPNvEqg5Zzq+0K
x4m5b+t/CSRQfUKSXqGPuY1UBnEUJcQ1774hJt9BWWgY01duw95vnYOd6cMddgy4
IPAfAJY7TqxSbjtNMpnJvp30848UwmXn9SUIP3GN01MKPNiaANO8x4C1eZZ5y8HI
SO1ZsSTuG6oG8JcrPf2ce63gY6u0D3Q0+adkmaGlnYaew21aHMzFtXS0N78htnJA
bxDpizaIPt5zI8GoY+cMfliF7PWTx9C3dG3/XC3YSDDI+hThxwRPMEsrMu+eKqfU
Bv3rbG2NafSPiGzipRg1DVuWMZhju8YRbBrZceazHoayLk5yNd9GroGNUOZ5Iscw
aQNRdx4eC7HYawucVM3v9jJEFYYje1j6FGNUigtQGeUT758AnfUjPyfcofceRboY
IsjevmeK6NkVDNx14g/O8RgB3ykB8TEC8eRVh0nNYWShMrmhrJ6nPRmKzw2UCxSP
OIWfrV1s3nwvAoh4fd/lf8OJe2XxaSPsf56rT4JSwy6PJ4QRMOgeXQ7WLlIYj9Lt
sOYwKrELdoSsuLw6DiQE8ctVWPFq49ZkkEzC969V64WTKPHcpjwT0QxD0n80LAst
cXrFAiKYmA4qQ5df6JE/Nqq1GJ/GY8VFj/82xK4BoIaVwLxZMQmxVYpV6Mdparec
7b+iuVy9joCBp+234n43MolN+eEQvZSvS8fHgjNcgA6ZK034Lc+cwpTkQWX56kkj
V1/R8VGsg7o+Lmr2wCtT7eVIphxWbNykOIA/U2aWCvNUy/598ORJ+4B9XLiKk5qM
SJRet0txm5zGk5lQEGr01uslA6MnW/wKE79N+JN7/dQ6M7CKtnhzuG1cDmhDJ13X
i+PvA3OX+3kX9RsxvU4NNT49XbBX2eX3+pfDD6mU14QfkpNg44iM1WYA09un4jNE
Os9Ofl2GA+1Qpb3dnTOVa79cCoX8g1IbX7k30np8RLNkWSYIWYecfhwsOiVLCitp
Q3Qe5wool6SDOY1HnYVCqaSY5Ng5tTwxgNR8ONN1XMWzxsZrPHCqKNYERSBDlunO
R04RPncVeyB+w0Z5MsLLwgFZ7VkNASNSKhidjDhqypGA0xE3wdBl/qAZwQj5pdKL
hrafHa3kS4u2t7iL+939fzjG+izcJ8F8yE9qx2DX1VMbAEQbhOHftYTO1KBNI+QP
XBBtkaFmX2S7Z6UssqBLhYQ9YksT0BunIjG22kHMgZhcRMvnDIvgnF56CQb2Zrsl
J2JkqZxEPOQR2bfd1JJOFjSGbLTgpvHy3ULjh1UsPYVn2PY4JkwoqYKKGpFhP2qr
u5dfRlTn0LuB2sRLUnSpKyLjEhOYd05AL53BQPVhGiQ+tghX4XFAdh+UveeEEejA
EjBotvcBpgeYK2BEjdhHTrmS+3r+WJ51VOQrhpPTGg/QhkQ4nVrnJKKSC23d5TTS
MjKw6MbJjoT38bCHjPnjptD2vBda5shJDbMOh8M0tu1q+O2YwfHUEn3+CsAfyTnP
sKxE/b9aL2Lw/hx1VfhXVGgNZ4Q7PiuGqJ2+RHCoAXdnEe+tQ4oL2kXkn5QpVXzN
ty8G6HbYa0eSiXxAH7mV8Zl5/Br2HQAL+BXDpEs8P9v/934/aA4JOBdmQ1m2teVx
nB08VQyyiXCUpWhmhZ0LEIutLh22gf6n+XH9EF4elSDxy7fZCrzKhHDX3t6f9+z7
3WNhV5wXL3Q27Y8wS+Ouf737jR0LQpWTir0AfdzqXSwcEoxvLw1US6LzRxjgPE5f
9R063LO52JaQE67dGM9+NXZkFudRxhubfUQO+zKZTUhYsevgxvUgAoneBl4u56nP
F5VvVKFSo8pacwHbj0JiL2QZMLeM5ZPY/JQAL4qpAi13bZADOvD6wBkyuXobEil1
jcCCLmCWwVoVghwp543r/vMuKLnGYWR91s8OiLR+/J3cK6w6bOEc5oli0kpgVVjC
YEmHu5wVhRQV94vTuBNa9Lg3+wuTVp+1hf1Jwc821B/pJdPMU3RhMdfrTMNkKytV
WWh2dzPT32VPXGhoeCIuno0kGy+8q7wZf90h8iU4WIGWP8OV1PY2wSUlPSDI0ymX
pPDMwyfMl8ydwPUdJ8cT15Z8zDlpk7iZHtfXBEddDoN8onjRrqAeMDtxPF6dmIrX
Kw/b/uMoIO7dVnceeQa45rzY1VZqONKXIicMUtMCBJjeThm9IUb16/NDDpB8qPgn
A6z5f8AvnT6HIXoQWNbYpt8WtYpY37d0Jcbq9vQO6ZUChVDO/0mLJgVJPcxV/fqE
Us1WjewzuMpDRj9gnsLRcPyAKd9jZ/oyClLV0we0LjrE6CNJf65rX+uC7GX07bmf
92atjQdJqIjFz5TREq0SdXseXY+lTKVG4RTyqRQ2Qje1i0GnElmoE/2ukkg5jID+
a6oOerpff5iLqO56u28rIxIW+DEZz099aDmkDaHBhpT1V36aSOml9zDpEW9fyML9
vti6Uuk1pvcG1tucDQsfmInnX9HD2jn5sCE23JoE7jvMrIZhzmPedlL9gxFTlC15
q3GeNtvrzzHQPC9DL3VjQ2hxb2g2vT4gjhJiCkjdaVBVKBuaSXge8ElZPHgIl+Yj
FC+A0svDCpMjjQVnbUlCvAYR/zsLTOlF6p0DUyY52wWRlUAH0juIpX3Z1DMcfqGq
pa0U+GNsyn7EFvJw51TOtEytOWNJ3xDeRCg+3pLmkvTcFk648nVhok7kBK5huP2C
Rgivj3ufzuntDuqDJHPZZJcaVvbGSIbN/h0qKsfp756lzyd2qOn2WWG/DT33QqTR
1q7LiSmq/AzYH+BuRer84xk15eSQ28P3/nmXf32p6BVfrsC4u2YjcKuCQSFLUaIw
imVOTJI7XBD/82yrm9HnWJrEgVyAdMmysz2S04jis2L15w1FX8yGW2Ec7lLC8j3f
VCWj1FtcLM2uiq5b7ZCfPO+ECEby4TUs4DAWE1e5HSlFS6YDqVJTlRaPxH1zJHjc
dhoXhqX8cyrqAyr0X8n9q3H1kRrCGXuJoF26YzBlLGtQyU2bYXLlmp100lOvsvvj
bbxvsJrFZ/qEJfLEERuhSBmDOT0YtKajxEHPgPjm+svUrAHTjo594Qh6+Q2qQmhm
XQQMhJi368g7Op6aQ0DlMH7XkSxldV3qk/0ssVPw20i5IX6gahhMcUtW4OX3AOLJ
ufeDbZjyAGWqrVDxwPv5+VzDWibX8T19QLk8GqWALG4ZyM0r1ZkUPxM5boQ7XQ8o
qurxIEin8JZZDWD8UKbAiGLShDC/vE2UyG4ATIqLlkCWRVlzcwhG/2xzcto6cR1x
98H4NFl3KX8/46zrfT6k826hcHtySnIIJ5MYwG2xBT7Sdf3/RVOw244P1+ZKnfBw
5Ww31ZVugEWk9Tl+VELEaD5Veqzrc4c8rKiKEITr6LY00Alkqjq8gi5HXNbNVEE4
tBlRT+ghpEj791DYx9psJhFmF1gOQVJzdM+/UmWqcESm3idwXOg7m8ffutcXCwOt
zkYm1xS+ER9w1UYuM8tS4E6cV2rlDyzm1uQoWknbxnUxbfGbf3laWgktjJkwifsx
fRbItyPZaCdkN34f77mWhoCsG1Ld8NMyN27dFWjgmjSuqMBfLFBpx5CAhBmyhmmQ
fXgn1IUSc6Bhfw+GscRBVRWrgZalaM6BppkOjGyTCHWHGwktliub2xXRSPQLinR8
753pI9BjiuNlhILdK7OTErn/c/VMXTsYw5QLKRcy7pVKqwip55vt5v5Ues4n+Hno
45nR5vNrHlJG9mN1tc2wb9PKpna7xqa8TGrBC8OOSFisy9fru85vNWVosfMcuODT
D/Ct1RZMxsWCBX5pftmKtLfp8tmbGX1u0lIGx3zbH5pOlkGvqH4sD/IrXmUjpt3K
CY0nPuITXpdv2jsvBzW1gIcCuKfw6z4/ErVsMfXPXY+OecAsppHv7xyLGQv6qRTW
THADcj9kRvb5DitMAnfhu3YuYL4/aPI2jhSO7aEaaaNGXrbRaoYXspejDZCIEfQ7
IFvVyvmmDuqj1YW180mY5pYYYeNrtzXpqfD/24lFFkmNyLcMlU+DQsEcXfRnRXSi
Wpr+hl9I5qO5pbbxzQShEXf5NU0wWioke5N8KdplIRuk96XRwSgndmt969whI15h
uDX71J6o07K/0BNjvy1ACmTQAFR0oiwxJ/YFF8RLZK99bR5XWzsrahS7/lNuxLCq
HXeyxgefKAFq2Izc/OxC5EZwoQD/3idMbDe4rz7RiuLfyOHBz5A7kvwMKMCEL00i
E1yYACY7Z80Y5xb1sip6ykLHGrgSaUCHB2XXIJBI5FyEG4FVakPA/a1tatfGK8t5
b+0YN5S7M4wNRQjeTh1gsebu4zaTskffyPyijVqHjzLA/MdKDOx3M5AXh1WRKF6+
EqTjziWsK+jS/AnCQdZ0X0H2VWqVB+BwJkbuh2kR/jX5M+jXM9hlcp+qbUVb1Og8
+6d/rv2mHUyCZ6/zqsgk93jsHb8A+pNUqvrFmbXYdMjW0iTTJu8PfwiufiXRNco2
JMPViE9p9NzMMlmHeG3kvP79dlSAFfGGc7xTnbVUrJbETpfixXQ+6kWzboGLVR+u
2n9HotyZHH67iGHm85rbX2LOwvvQBqQX3OlGtOdPSmJ4E2HvRWSEmJKnzZ1EyiW6
BAZYVIJt6Y8rKxK/C5OwWdhQ5NKqVpGTsytrqK4RyFfHmNQvvQRTEzpCLf1Xrz6C
erivsW3m6UF42C/Ik8Q5hdW+j5lMbQCEUggCjWY4QIyHXg1eO8MY9bQ4LaZAhxL4
+C2ctEos78Rln9HMEbbirHNtHHR9SpaMZxQPldma/xE71jgSddtVfybES7heH5DS
CnK6BPRJfDKsOtOQqNThFxrFsQOOXDl8hRl7zLLcg6SdUhvan/yKb7nB9JO0VWKZ
8y/643MAnJavPWE5Uip+ucGgXzfXHt8QDEwSD3zuutUQii/QlDiCokt4ih6B+crZ
oJjXvToDKFRiaKEQBl9njnS8/aKtfh3/NAeRWd+kW2kQ1Ek4vBM0Ek/a5wa/zJVo
B4AUEqJFxqYcQGTdm6nTYgp2zFx9UUecJ16yXozD2R1WfMSGxB7djTA9fMT6heQk
TQrW5NmZNjbtOrC36nnPdz8yZSn4WL4yseo+Ux75Jb40//u/XpOOlqX9BeiXM3Vb
8TLf5FYDkbK18o1oEbqT23fpf62jJG4fyckJ68J6uLQh/BEeyKL2QBmGRcUJtlbK
g9ffnCPMaBUYc73IbjeIH5Z4OobueDWfuodlezdTQML1oyL/C6i6kZPsBWnb67V7
XAT56qKQ8gKlKwI9YgkWEW+FSpJrSmSWTR8ZNMQK/7dccHJrCLpnOORiMVmEyeDy
Tl4H5l1yzGG0xSefUErc0upNLCd8j/TRuUaWgRJQK2m5IDeJKrmyyNNCULzpYF6/
3LXwAkWo1JIjovuG/ry+dD8z/ydj/71jnZiKKCun6AGqMr2OhqSCAM3QqTghGY7w
WCQqUjSnbYZWAcPol8hdwkVhBSQip6lScVjNv33G+5Fkbkl6ZjJo18JvKx4H16AA
gfPiXDZhYHknuGaUoAOIL1XGYnTLH5/+i7zVRGXHN+2WswZY5mnjgJtUOKMfN83h
nK2gbH23qwb/jl+lpaL0du0q1ce1vH7X8u1ljFyR1NhK2FoDpy/PDtUtjMJK6T1R
TMPqhiC1+fKk9J3Z7Vbe2cSKaS8KV3J7bpZ4BB/HEoowZ81ptEv/ccDqiB/FLMJ1
DhUB5IbigUY17E8vQp0CN/tBCKT5qjzksSeOOMgtJqlldKzKYqdlSN/3e/XEyFEm
5k313T7loUol3KULG/QdxnrX+YfZW/zq8I3juLZuwDh/BBXHTT2gdEnlxI6V3S/+
h6bTVbYELfncwRTCF+ZAUDzlemSv+I+pIAQ3YkP/8soFEBBs03w90nqMbYDyeRK+
0Sf8rNmAczb+ZnQq6yepEBrlEaCZDpokrSjMENlIRvVoJDCa/rQmDkLgbkiHPFjQ
9sBllV52m0pdZE3etUaevSyplqf8iNL0SgjImAnFVe/PVMhsO9oaBUottVzn4vIs
SNsCtQs5eNy+l9D7XYDFP3RVUgKi1fAE59uMjDDYJ9pJJCFX8Ecsdd5+9d7ENsuQ
xO+iPFbg70pO6RwlRPKiFTB0AcGdAsx2iKduhepxBXvZ8PcjIeatTxQVtQKCYQAg
iiNrDdBEIEvqfkeP4vXCNnwNjqTXslo1EMBRWGtQLg7+M4VMTHO1nRpCy3BepQ4D
tDjpScJe/ZBeJGz+rVhZmA85t3JtjXpM3cFt2O5eAs3V2ppVdi7fI/75UIy4pqyk
fmje2n0MBmDPJsZpWTC/kg1er5ahWHgJ7o9lOKPv9haUfw9t8nP/N3oWXcWQ5c4D
U5CQup1txBTwVvgjzLiyGT5z0joBQY7bkGOezmNy7fbYc+S61n34Rgl2VlkjBjcw
bprItEvLn8onEkVeTh+iwzchFJQOya0FS8WPeSqRCTVH/84hmF6iuglQ2+sPbu5v
CQrkC6hXW+twG3XPvzegqkGrKGZL1TmqexIL1ULvc559yjiLNa3VhHYL3a4yFURS
bCHQJdgQBNCrgZ1gf9+BhY3g/45xQ6J7kwG1AiydBjL0Kr4lqJyv1wV4Okk5Bx7F
B0qGRjH9M64D5xJR3VJy7FnGsxDy0Y2yyFKP8uNuWiE+LUTpsdsfzhnzlA90kdUH
PzG42TNgOC5ijzKemVQyGlUdVwbl/gDyG9mhy8wP7vCDsd1UgrtDRB2LCGh7380l
22CaHw6Tn1snFNXZ5gUJtJlBtuwv1DVp57ISVrOH1uIAeNI7IH3Qd2pS5JLv4rtN
37m9o/5Kko7kFySovaMVPWroCBBzd9Se0IIh14/3PUC3WrJT0kmAEhevNPEVM/pN
dEcihEOd7X/ZbEk+Loh5nVdUiBcPDu6KjO96szBGTlJ80cvGg2rlvQtn4ulm7ptc
miBr3Hc7X0z4EoWv8MR1BJXN2lq3D4CS2RCj3z2MmMGeRa8tbhn/DFBfOK02mFlR
CXXmINZfFHjwbbNQZ6h6altQdM0Q7pN/gVURPmPBaf+lcqnBza15ic+os/K6xVR+
nwWOYs3Vh3SGmdWavWpPO5fvrKDFetWGtY9nvTnPm8hFI69jfK4Q3NAfmAr8knxh
o9D4c+2kIatQW3L5CBvJOMKsepM5sXPFETfE75zEBnd34L9And5Rp20tTpJl9C/i
6KDSi9lUj1d5ul7qggflTcoiG03xgVqDfyyUfsNGbHnNorSVmiwTryH8QjQPoWD3
1woXzLlYr46zlVXR9IfYEkOz2Pxi1tvrAN451F+2Gmi62tOU9z9xbmvivfZEJHKH
eU6pLu4jVDoQcY7q6b7AT6yN+1E0zaDpkTIVByJcmiGZTt+pfuDfDPyWJG1MjoaR
NJbr6uQ5RjPuY919V7w4ryDga/u97V+9YW7M8g54VtA5C4iPewa/baShwdAXQtfX
spyUmqkFedRhaCqHc6u5/7cgZU0WoMLLA8yepMF4BBkPmbjZRByah5zbzvscRFcb
1MszJNNQTGQZ9i0VsxZf4JCSWZEqqv+/Rjzs/LAePbkrcUQKPrly5/3YkavYkUhi
8CvC1jnCeD5AKCqiaAnUdXG5pTELFpgrcVZXuiqnKdt8k2AJKwaTk8HQHbWQuiXS
75aahqidqKmzqTNMsps3nFmDuCarxJr2fZHROE12SqCDhyRWd07kdJGBpfNykVhn
zZ9kUFe9Yi8Hrb+SxYBVcy69Z9M+S1vggv+Qsqa2IIRyYKsrRmbr32WN2WyKv2+a
tCABMfPM+wQjgBOcyIpT0s2U6k/zBwjXHhRwzbfhCmNGrVfTlTiw95ofhr9/hwG+
+OmB8XQ9IMHpBZp2pyrFp4ew+elGECaJomU7jJTmlznLPUGlqqS9NdTgyWDVXzG8
nAle/ZIp5y3De9lCPs72PFuEksk6PupogTC0QIMhby/9T4SWpJ6XYLWeJ7dXkNPz
bo50BK8/pOiV3O/SoqEd7hrzqX/TmpyYqTei+CJKrkC6OFU0tfzT7h8Av6oSGtJP
O+bSSJYLvpne2k0koP+5liQ3Gae0J2mFW+b1b9NuB9rO2v9wk4nK8WmcKEOW/dfJ
WeUVWIZqXtYt/tGLmuSl2BoJY+Wl/DRpzOznPjSn9nVzrjZRpAEAz6VXa1TghA3+
2ziFgGGpdmevmDDeliJ1OokWAjJ25Lx7OyWwofzqasoXMz+lmehJWDKU3qAwIn0G
0YNdP/VRKm9GErsI0VGaGOIAH2sEXtY888Shd0dWoi1OZw+vxxRI3oL++xaMTn35
qJj59E9Ubs3UHR+2b/ZukugVPcZVApFUUbSBSQ/B0zi8jz5V25e/r07nGy3HSYcV
u9jnCXW2ls/mxh/Bw4owszXefZzdBKFVeb1GKqDx0Ohb8Gn6yJnIqNuSBGlG4CN5
QdRwdEeF3TS859lb7Rl9VoaUWJInKTWTaXaahj2vilZjAZRj5DxbgM0azz4szF+k
UVPv0lftlYyFOiuAHfr2fXohlkl58/OqliluePlUASajDl8brh/yRS16SYJgXuTi
W8WH0QHMvs8yh71YGWPwRcEa9okFUpVEbJUAl728K6dGQmVNhtLE9KimVyw6osKE
ruVctQwr10nE7b7WUOIFuiUurCzCBov3b9MXVhnQ04X3/5/1PKTbZx35X8L96NWp
S9tIHaK33ggoKSoMAdyWyl6t/T/USW3tHkfTVVS9mMdBh1i252rsnRJdvhz4A546
GTMScirL2Z+KX9TfyBFdmSGMLHA0hkA1VceEkYc9/ct0yfmQsnD6+dt/H30ro7hk
R03M2GuiHhRpPesT3d+p8Xi1uyzbGWTIQLyw/bUEUPJww8T+7FDxGZsIKdJ+pXzJ
PLr/bJTpJ8gOHee1vVHqfDmra/vP1QxD+yvnseAlmUnuyWCXbDp2fAU5nV6F5Ady
auBM1mOuu1IpJwpcY7sFCQVxyfGoI8sqK4/6Ta0MbxhLrSWamujhpj0dwB4oQNxh
oA1JCWZ8bbGC5oKNqshafjT3PaSqugtH5zccCjGNWy9I0wXZxfC5i+zMTtkiAY+b
qIC+8C08Z5CToLrA0YFL+wLJnWCX5Q/hbE6c4m88eHNRhW0RPfjh2NavX1c2gGlh
r1l93aZThse558EUixN8Uc5XZ4uu6Q/qJm4uo7y5otZxTc0ZQwmXLomv5j9AfRfP
pnNgSfgFQER55kn0rz/SyS4TmPjVNR3poCwcEl3R0iZJgoeFYWuz9unR1KIPDQtk
qWR23+FM4VqNoP7dxDUBIDz4Q++OErVeOiZsDAWPknTi8IN2o2eUBlYL87UcuX97
eat+0UR8M0EPh31/64lihenYf87zeCKx+/gxYDLe+2ukpfl/W2RemW2IeWcyGmMw
XdqJhmSVI5HRas57Wfbk5EE1iQNr7WCWJFM8VwoRSpBkXLXnlWYnztPhArA2zBP2
7iNMRtZGJ2+FULMUTQpw4otRWiTr6EePFxZNTxofpKb3Pqn3DtPNw+8WdC6npGXn
d5NuUg4L5v8vzaKFUCWXuk5CRNRvFa8rE06Na7rujZoJxZn4ZRy9/a9tLbKabsL/
Lm5j+WWaDTMmLK2psMsJGigswyHTsrmrqLDypVhc02QsVFalCzd7XtTmc4we7A0d
L9Gojc04MYNDk2frFjLHmqSwUz1KxzG98guLVrSa2QoUG+C80hIWH+CYInqxrSMx
OcrUD3vnSythOC/AkvNBhceMXUNMtBEihKEGjWrgJJ+2775THMOHD5k+zTqtteFe
EZrzzOQJgMxvxPZRy5JipTNaeHmklbg+ANOd7D2ghNSt9x2POtyt7yERyfhUClsh
fEXF4pWAXtGmmdv508+YY7Ze8lQBe/etpNbjEyvYYljHJ+qv7kDrVAPNRlHhtqAo
f+YVlaeTyOlpQUbToErCWNXrMPWt93n/gBjH8qsPMe2JhX2EvYbDEN0sWBFjhMam
0UzbIGJ9YAuyh80NFRaGISDnvSQhpdDjVe75HOQlseDXp90JW6tKbcIzlBHEFJ+V
olVXHkzu9HO5nFETUEO6f9I+l7mYOIwJmGxCFXx8j+gEwLouPbuoiZbR/VuDTQfV
0GeYoD/FDh914ZNDu/GIQOohtb6PrhJG5/0l5VbBBq1dyHP8NDwUaQujPwoWVgBg
yBvTGK4o5lOHo7RR5IZHvwFMs8Y4mgLGSHqFiyeuSTXiOi1N2IzXcAAJNOkbep+9
NpTQGOE01N7Zgq0JL0y31vC/YacZ+lMw7B/a4vOR+Y+U0aye41B8eh7WKb9LdesK
Q3k5JiyKaCS0nKjqDuiHHZy7pUDgdo3cQT37VMtsOsECDskPh9GXJiC003pRuBON
E7icZpFPyT6Mfc6Oe95MAXQzhAMR2m/LExs52dMvIKxKlSnV7W7FR40eI/QkCg6o
1HzLKBCoj6ALX5VNHILM8vl4Jse/J8nIynn5ATHo6FUOc7mLzNbBCYQIUvrLlbyq
RWlqbEFHj/AqAoRSgK3qdQfDjUGnXSS4PRH/6dC4ugJL2Mr7aqX0qrq3SIyRh3Sr
SsTa1QPouzTWbEHtv8BTaEzrzw0dNbALe0JjgaGAFYJoSSEYg71puyKo1lYNg5dR
LEPc2NRw2W7ZZxhQ4+89YIRHmaL1sMckYux9I6oMXtVRkjun6AxUzCjlLaTtEYd3
I9FhUXuNz3zzwI3mupL0jEb0c8txwNQQ4hKvL0+1wJDlUphfBXpJdte8NrR6XXDS
heiRG6GaKUYWEHzTtLe8INj79W+tGM64SPZouWcqX+nvQQgiWdAzgiv75ui4cqOs
tV7zIpYcpFUp02Hnk4BR00GH5qZBA97tA4NW1xYYSV5ydusyo9WHDF7K3NZFxdYE
gij3NiOvgqgD/MQISAJSEMupeMtifKdkz+72EsO1bIBAVb2GGQecvEyulnM1a5Sr
EwDRjx05keHEpg9+Eybc59NGczYEoocmJ5pMlk+qvFAZWgiTkmYPSgYj+6AiN7kR
J4YPmHGAkvicf4kkgrR0QtWuIIl43uZ06o700MkLEDXBbfmDMfNi3E1PeGVmWnev
5wjHmiZKpRk5tfZw5WsoDdO55ysFgHyLkKV6lp7bKixlVjfm034UCLp1Hx0SmzEr
9S7mdiSdze4tOTi/1aXug3Bn9/2ixI6yfnU0WF+Yh5+hGP5M5O2lZ2Yz74qo+PvJ
Pd23ZUmXigSOrWOwyZ5d91On4eQ+fnh4Fh9ouD/4QRYQwQ+6V0MxTJGu+iik4D0e
9hJZRng61pOkrgo/9tgA70PmJ/OkhlZQ91Gih9r6fqF13tS//MjLsRCackfFn/ng
3szAGim43CJPlQ93KRV7iqycmZOT6Pkf90VxjHf2nF79grucZ2L6HF9TvHY83kbr
IWJwQhnQ+8zd8/jgnsPJzmV4RsI9OQRlaiIqOpLv2CAbvuJIAzAhgY36eLzeox8k
Ipz2mDmWZ4Qi1qB0esyZP3bTgh78CiG1ILfe/ZenoFJptnjiqSUQHtcj5VFwX4c4
qTWZmDhAV8aOTAw+94mfJrVVgGNGWoNiPkj3rHox7vJeE12U/6QxliLS05DiD2/c
KgElizSlox5LieR2tyiStCbV7UPzrFSVtF+jPX+tjK43V3RraMl9i1Halbd86hlv
GB9I71R98uKEhJ/lw5ynIUi1Qyi7WxxZm8m5O9+3Qu0cHM2wyVPqhPXuqKdsjHFN
/ocJEeZWeezWvwT/9k7dIp/q1SfpeEZj4t0UfeQAVgqDU6HCI966wJ3IChG9t7on
DDm1boRNoYHPr2dHUCGR2/cRSDXD/5ozNAyTTYenCeV/rLpWb7EkSqg2ElqZ06nj
W0MKZgC17Ezu4EH3ZP1yJxiQ/dtxrILKNfv5pi6+kfGy6Pm5TiGTWGvPAAlY2rMY
NMKKyLQ+fNp1MS9m0LfLbgUAkmTLC40sVycd60tHAkOmaYIlKeQQfP4odH8e81Bg
eHba9V4bf7SKzj68JTepiKBg3VIKCkei1Ht9TW4ZZJk3I4iG6WRMUNrG3fkH9/Xy
RvBaIcnSw1S11uc+jUfLnFEZpBLdVvdh8wuwypOwExNH4DJmyQj9UuTItM9Oxcfj
2LGN+FHflc8A+OrnfydFzTjFSCpUobpmF0ROPIA22Oy1Yp2I/h7KmX6Www3pJ3fC
ulbDoD7d67bqiSWItC51hOW7hMSI+A+lG4WucRBL6hfa2EflAOO0Iu8tqeciFkIj
3RvsfVjAyUkPAWi17F6dZy309V/vuUew0pI2rRRfzZfAW4eRD2NNpsG83ZQBm1gM
JtxnsHWwXrxd//Np+HwB8d4OciX7NVSem1MJca3w3zNWSdVtKUi/OT6V9S6nwkY4
JP4QhZImv4cJJx8LZpla3AqS7N65c2xlna0dK7OK3N0VsJx+/7ChEBFI66/9EFE8
ocKbiS8nZX2Dkkb+8CpoHKn35lCMbIr96ENti4WBDeRwPUubtO3x0YEbCSYTlo9b
1a5SiagA7xk2D2nn/KtNbUaoZP3cSE5b7QNzOoF0CLDlswrdQAZjE9x1SY804zJ7
FCfwWCLc3f8E/XWIq9MUpPB0ivG+fDoj72Lns34IT/DQA56Umjj+0swHlBrDP1an
mFsnfMEZwUclvWw1p55r5Lni0RwYhxb89nx9lQmfJhopwPXa+yAY2Uigh1Wg9xtC
QMNjZ0R21X/7YOsEjlohgnCNEvV4HzgKoslvdVvDGoLpZa6I8nEZpYkHPiyB4qyS
I4gc4kiG/3UNP/Gqt5lZXKDfb94qwL/cB/pKhYL4JLUxLr8UskMtyNqBcWOWqVOO
y1S0L5jzeHhs22ODxXZFUvXBXvDSeLxWSkNPPkW+vgHm6DN27bwO3XsP1dT7UlUn
TdjYz67YIrT2gsO5dsxiCbwVbWgU6Q6cO3vzbfdimEY2K85OsJvnnSwUEMJ7ro3V
dYSR/DExmMPPfuYFfdK/yrsle7wttTT+5JSkofAT9sZsUI4Kep23ew8eKDZVwF3Y
11ODu9LJToKKCL8vr4re24zFJ+sKLRTESmBhStnNsn3KdYppXpvNMDQUEQnJCOjm
A8urw78uQMdJoDrpY08OLepfx9F6tXzcI0HZ5ccc74abzNes8L9WNuPrt2y1UnP6
JVw7LHsythp1A+aLgOpF2t4U/kO296x0QQJP9uaQZTWq8V3c36wjAGNe4wP6+f2h
wrf5/ZA1wsEt929DFuD4cI7j5CTmgntiSnQv8fRfz+4zbkki5q5Rb8C5ipxlJrjJ
XEUx0ezTY8HT267JtVrsc2YpyHdHQx9fJRgpSy+WsK2f48+Jx+4rxDiozTrKlk9U
jra0dXZy8ower89jwOS8+GTtntQaQMDj53UHSQeHV584owNeXaUvZo8+xQzqt1zg
SHKWTTiOjOsmuB7RcZuxdu8DsUZ+BVV4S4rluFIaMquV/LGxFgVIDo1SEumUceSa
5Pk0lLqwiAn0SHUJgajmz5fNJRS0edZ9tk8uWUmbIWbxT9Y1cJj3DFxo3q9JBt1C
hRsErOjTf977hvitycPL2K9SiFxeggtL4cAlyTwJjCWwbxBLDo0Ko9oFojOmUIm2
QVBoxyPXnyu0wDbDJSRaNYAjy7NIgL1g6SSyl35lBNNSDZpmHzKuxi4lQoEF/7QT
Mcf4s5UFeHmTOvMY/cyhwE5qQ98yz5WIvXdz2Rp3JelHSY5l9mJVrT3Jhl4drLEW
Knu+lYJOp6Nl+PJYxrxVaA4kC35jV/KOTYkus7FDjwC5Fv1KKUCcr+LUUmDvF1/P
Ubp7POTD5tf4kkUwejfmdXOp1KSU6SQPwiUaexVIr1GjuhcugmElhsn8MBqepxzA
z/5NLHXk+2+xQN/UVn5zaebo5ZCcmtHj92YlvHE17MWrKg1xllC9M7RV3OJ8hULU
sM/QVFq/SplNAX9b1PT2ZZr/nSTW2IGPUIjdjvitFHuM+ammRPxHBVRhctJz9Pqg
6sbPRTvRqh6CWZrFr4Wz84ovbOsLgkgiQwKjciz8CzvBFmpZompkwrSbRGrUwmAO
uQlKaPGSW7HQj673tnkHz3bI82inaHTECUHossentyAjAwdMePO8F4lwM5gNRE3G
PUNMDSB4EStbDDs454Z0Rj0XpZjFwdSSWR5/QSXsFH8iQkltlwPG2mT9Kt1i8Ibm
DfPof3oPi4h2Ls63ZQd7w1adVerq/O8ECeNtEi4OBMp9gCKtixUo7xrc9bWXS1pp
P6Zd89AvAt19RdObrlnE/rQmr54JXovpQMI0k5aojWqKYOdyHGBQpP+jN/9JoLAX
zcAOYJb6DNNTJXS5nRDIXDjcwgam+mTNHiJpWe5CR0Dzbi3Kc/JiVQCFkl/n2pVw
s3QivlxfM9iCnk316MAicm8V7SONAR+DqPG6Vq+YDQAbAmyXN0MsOBklWDnVcelq
v/PJ2GadlI0e6bTkJ8EZorPKeJ7T3yWXYbKR/dX+jYZFdbt25HphQjknmCf1sDF2
xrbTwu5khB5XW0pKfr3RkjV11Vzp1JqxZQbOjNhVTHfpQMgBBW/lhsc90VNwAGJH
xS6qfH1ljqS66zUZha38eBeTc9U74NLWX/DWjdz3S2qOymXgbCOTEqcDey+uF8SU
CyL/fvdBNFGT1N838JaWbEApRL+u7cNYK+qAmE4APnUe0eUeXFLklJBjLygvzZ4L
mirCuGUxQO4HpXdTTMkMHSyhOeDGARe8QSiQJ0iJj6WT0IWp4ApdStdl/x+/daZ0
qzUFg9rDzDGpJ3ag4XEeraPGvgKMWfR+s/e+yTBH7yc5BuQrU+kRAaYwlJT+AEke
fdEfhmOnnBuc1JEh2p+6sKHUlbZJ6lIX4+eInCbTNxbFQeAxN8jh7EZfT60RXBlM
8Fqt8t2vN/ZfKwxUK0wbEd3XO8FZDRbocSYl9B0FANcNaSj1ktGU4XVIP17RyTjM
01jZb6WSaRx2H5fP+hOgbQcI4d4GKhs6ObDLlwBttmVdZ0Df2yWfRhbx7L0oCvtm
A0D/TctQ8uBdoCfwKe+M1b5iB7/eN2OQYVrAJgxAj0xHkTrtiO16yIUbomDVfBlQ
GRNLNZZY8EUl0H2zKlck25CFZibSuYia1MWN15CngMiSo+G5D22fKIvocfZKIqsI
XrKXqsffE8BuswUF8FxX0rmtn0DFRGJn+y6aen+wo0JZM2O+IYxb6ksrfGfsbXby
uK52VGi2FCgbDlwrvVtlt1rzE+5jnF4DleCUpCZ9qFeEt5MQm2nRiSVAho+W0Mk1
RsMPjEMn50WKwZntfbC/Ideg/9sukPK5GhADFQdNWYHEUXZoQckcwYoCOJjhibNR
YjkaF2Ry9mkfu8A+5qz71AI78NAnGnAXJqAPBjquKx2oEKg1Xp8Z+buTDXlBsmgE
yk6ljgQ1GCqBJfykp8Qz0hksrBUwezprJ8fMv9cJZH9Vyi/JHychS7EVtDwDKd+J
IrcSeXOdQmGsXGxb7cJoKFnVBYHCTQO+ELJPrfE11OKFidzByXYiJGfB02LdAuax
CX1hsWEfZDqKMPdVGoKDuSDy8tv74BSfB2RflURMSmhrzM4zNwmPuNAwIso6aIt6
GVOsjgVscGbPpfAYRbNXgGoCuQy9GzzWLNphgWpHJVYoI+pIk1rJpJMPMGR8nrMu
+liYzPiL76XMJ1FnoYaBfxrZXotaEjgdWNsgiVVZp4QDGYXH+OsCDQWXHiB1ELgu
/OBMLIAFZ0SMCPE4rq71QiyQfQ7OAref0OLlDDxcpEPrnaa96gINI1hgiCi+C7ke
Bd7rJD9KbPMu5Aj9G1N43VcnZ6qegzap122a7JJBXvqek4TNEVHTSets0Qoo3wF4
5axDGR5XclVWswFfxGJz+hUBInPjh6bEF6GZRKkNBvW43ID07R+WTvPsdNs8qL9S
sz4OyrWWnajG7YlXfTFEJSm2wta1gAmH1A0PZ8mK7VNPMa89XcBnErG+vxnaGm5Q
PsEKZ/4ps/6eeJxN96Qnu5kBt3uvEu0u3jcuq/YOEif+zWZCO81Rr5eRbQYCspqx
W4SIsUYtAH6xPb6nG9JJmWVctZlHy1mSfJ4UoxcIcLl25REXtZjI6UwmJcpjJF+7
eC7qguOpnjcoUwRRVboOdap6hP/HTF14RzlVkOxdMJ60rS2v4sL4SOhfrEqprmAw
xdlws3btSd8YXsT475ZFtAVqMnv6GgFCVuBrHR98DhmpZEIzWLjm3ZeuDMd8QRtr
GEFPgywLIj2nhD43nSe7DoMgE9PdW06Qw2A0HQSfhRCueLhMDRoJ6XMG5MUOMtVg
cncgeVxVTlEdzuj85KZ+sd0x0OaWhA3v+siDabTDYck5U6FaW6RPctt9cZtyQF0w
lflCpvLsPQvbBM9vYGeFaGiYZLfR6wsSlJCrjM+21JncNgQhd3+azmKyLAdqdJvq
QySRA+BL9il3IxZqcqLLf2yxQwUhyXAmsNsjYSCnslPIZqSxKI9iHAkO+P1Jmj8B
gWcwxbsWWZNcWBf97IIg7+KR0FbhzGXhePDMJnjtHDPvbf+jlx9S5QLt0wB97jUe
Pm54Av7Aw5m9DBOp/9LUWqWOfOfvKrCLKDoWsj+A/3szwkVajf1Lmylo57R6kFiF
sRv30G8P7QEClvR6ZUUEA3VIUO8O5pM96/S6EHGYr+B76VyUmuSg559o5UveYQfr
ewTwb2xpZzqH5au7CQ78wux/bsMi0WwNVBa39blgie6VdolkBDHWeQX001Dgd90s
CZNhMbzfxgYfgRe8rP7ffE4TqKWyc/RuI1sD7SYePJr4ovXbk3JB2cvQdimCTmra
/XI2QiVcCJ/LA6i2MBhmFza3RwTqvD87VCb+URvLbG8C59JvNNbeRai9K2dx9cmW
s7pVLXBA3OYukYXOHXlWPKWregDJDxS5fA4NBNkBAPWKmOCiuSQV2XuqdFpkRcV/
deFcGIybvDwz5V2fPBwNb808JVqrf/ZVJH+IrEkCkTOfbKeKDbBLP+eVGOQTDaVZ
UZfhnaIVwu78SoLJa3MirYTT5f6bB4jyq+iTw/LshVBidcibzCgZekNLLtbq5jFy
6wl/luskYulUt7NQmurKsvjq2I0RE8tE4yR6ByY5YQ1JwhCUWyF6NK2nG6jE1E/k
n9DUa5ZWt/JYqah2o6FvkJBhExcWFd+6wLBnE25Id5Iq8GfKqmOT8nxLCVcCrRYq
KXwLteCKw4SDyNfZcd+ixwtg28s/Y60vrftkeBhrqNuVIQXJwT6s1cYww/ZAUiK+
8U4zGo40AH6DUGEB8oBsEIAR9eGOe5/y4D62xz8BM1m+AgHm6FLFOvS3GqDGstzf
7FvobuVwfo5Urt1ehA909MifT5Ecif8UdAvlA+gzl7WWtXPq7SKes55QBpDlC6Fo
Vj4uIvs1pFnUTYs/A4HDmQfBYifD6f7u5CsbhExiMj0SHACurmdqvjL4oPUKFP1u
kukCVauFi1eLqcrHqL6HTaRMjV3Xqit5k9cNVsdt4DusrXrFTRXdKaXWps13CDKl
8O5J+TZ4jbJJdYTHeRwcC5ruTmOup5YXOEI2K3t+5V/UdUiD3jELO9YAsGK3C/V2
YJSkW6MkGRuIalTwCDfMTJqKht03NPREHTA3Yurc0uPqDnNLviy3wsbqlbdQ7T4n
o7DQvC3Mh/ETSk2qifdk8V4D1WvnAlH0YUwxwmUlwQtWzrcmlj6d+otpawWkpRvg
vcmjHRhoX7Bns5Jwkp04GMOlpzZ0m18yrtGYlgkD2PvgV+sQQdBdh3+ZZkumG01m
Y0XRJE01GWAEUPQLBv4zKhLnF5qC7xeUqUVneXE/ApLe/oC916fwoc59doRUBiTH
2XvV15WemVElQFPDHv+EMmEZ6u09yakhj9z5sg8Os4yA5qbkTSxLIA3l3iwd43ya
utnCCzKkcDLsOK82VM65SknV2EhoUXuaLVzqZeiTyUQL6ga+81PheM39s+hYQQgX
sGE0o0sDZ+3agrfd1m2F2ofJdOCeXcrr8Ajlwz2DIZAMITI23G33Hx3PQ2MDXEhG
mzSngjA3n3J/z6CErNJ+52vIaTOwCENJNOfe+v1oAV9lzMDBoRkZsmDP78F4izlO
9EVQ84pV9CqPFNz9tSZrglkq9hw9bfw6RoHwDtvV6T0cgYu2QpU9nzK2gha+wpAW
GHWJYBE09yGihhmrNW0GGShfoJtcaY0JeNvZTDpr5QNae1pawAPhZnxrL4a03LkV
9xVOPZCdlgRpNOzN6I86wVLFkYpalaxC25rTZRpwS/MUy96tUJvYBVqyc6+6sDYn
XX/w/CYBrwIrTnXzGJ5l416JBZtHy4cXC5fV9ehfW4gj91nAOdD60HgNae/tr5bi
fNylEFaFw0iliQz0fGHbQJkgFhxhERaf2SeAbMoXu4XF7pC5uEibZGdIGwjW2Ulv
qirP65nTaRECK6k2oHoZAzGj+EfOarb1x3XBsw/HhYh+Ni1FtfYdjz3yNI8aqg4Z
0o/wL1dvjuEg9X3mHhV3RtxtGMC5BAToy5hoQ6rmCokGaBsNKMj3CDcBXEGdilWh
JwPI3OUWS566H3b+8DrWBGFBoj+4OzkirDsMvRNwx5JnhZtTopi1r6kd6knwh3EO
NuHWHEWnliRnxA5A99n8juD/PnaMcUEv1toYqZYzWH7MD3zNsb5oUh2Y0ZXO+mKq
J6anej7VLySy0lChsPxvdOXBjKQUztceuLCvUyDBrwaFRuQ6v0BzsYSWu+V9f3F3
BASFVkPQWNz/FfpWKoJcCWhucGm95cqb7ZUx6HyyHPPUGbsmWUwP0pEykKbTEQs5
KC3hFOB/aLkbvKN/o9Uw8lLdMAy8jGM8oDq4VELL2bdDNiKoHqEwEoGHW9Ru26Q0
eoFa057OmfWN99Xt2JF+6W2/WainAPvYp8nxfAb5k2dn7pR1IqeMMGaBLDGtWk9o
BbvD44m1r6D85ZNZhbEffkr3RIIAPHXF201FntE8UScwAXYeRbWKnqdep1YauQtg
ZfHITjGRgsuDPnVLoPGsEpUpAM2fJqkCOWbWmbUzPAgBwHf8o9l232IygVTYlCAi
aQliNjGnLlqwN3rZ51d4BOeDqLznv8FmqQLBw5kzKpwQZj43bjFdEZmB46bQ3QT9
Elon5O/AVYkJV24fcmfkd5CzCmN1A4hofx/viQ3PtmcpkNyv01QUvu2VHMXPybve
rLaFSbC2Zd4NPP24P8kH5AbcyPfXm40RMvjh1Fl2ibjHeGofEW1g9b80s4AN0bUG
eYfva8CU5R5MZj98W8uSOWupz4fwvecNtZvc2/wA23cS7Q3K69SZyV+64qmmma5A
ehBizuUaVZGKbRLz0+J2HLTE2tKL2tQe7jMvGk+2sSiauqyGvJQ8u+faP8xZ+wL4
OElCE5xbOik0B80QNl7WCq2J4fS5CSy0AS+BKbH8/az7FZJTi6byrMAn4qjmVtFO
zp/4lPD7id/c76nPE7p14I2j1tOQ3RH+zoBUmpSbMd9H4ODET8t+umgrI23nYo8L
IzB6uSFrABN+aBuQc8W4vX97E6VtMyc3CaFGdbBcgq+BNvDTsrDZEJbPlM53axtM
5Cx+MQ2iIK0fDN0VOyNZ56E+Y+706gH1sHKHjIoxCZq2CUPEpmPwbsH/O9pBtEZz
JzPYYSzxz5LbN2fix+y8azAgiATKEPyQlsICSw5v5GsM/qCUVseB6KzSbsNK9P9n
ZY+8S6zOBV9EhYK3fTDzxz5z+Tx3cyI3aOh6n2t9RFo+IGhFMWcxZdQiKwrBxCKt
/doA3407PWCLB/SdehYF+3CTIENHjAxTwPmDEX6oCI+hAKg8NVtMrcjhFpuxBsxc
pMmpFs/Zp7wUKsmPLs3qmFhV+WNsDB1ZyJEai9feDNiIxy/NgAczmbT2/ry9Kh1c
AS0XAmZf6rjulsoApYgr4JJGiwjoqzMs8KFXbo3fylCoMyrCR0qZpePnvIPSRnfi
rnLUl93zXkAm/RcQpj5sj7CJtfNhcRbkbxlf/ae8ReIMXUmUW6qFvmyJXqY6OG6T
0GqZNpRsY3jvpRdenQDHAiCPVx1HE725pcbX1x/MUVHVuJWPIY35RsMMZK7PVtiW
mLJgPuFpqw3J71dH8ylPOHc8YnoZyuzCdIYxoMl14aIHJ6ARNhqJO2g5yfI+YzIC
bYmAoAUimoYtELIlaZd4zH2H4XG/hmnvfmw3rxkfUZ3e4MaKlb17bHOlT+8C3HqZ
VJoiJ7kt1rUXFS5eqZ43b2TAVzERZ7WpS3aW9rC8ZRQTueaSSWA/FzyVog+PYlsL
9qL2gQGcHcDfPFJYG3ewv0UppcYh12qiwTsuOStPDa31klBHmdSbxyto5puIB/PB
eiwbfFbF5WQovP/2TyElkds2Dlh8PXt9qzv7IRdANheKhPCuMXE1bPQNf2KXI3G4
d3zyPJRkRZJiUBTlUDGQJjUBRQrupBtiF3K/glJAqUPtrAGkrnnpofa4txpOXzO9
2fJw6/h0qlkFIQAFm2T7GdygSc5t1zQbsU2arjP01kPmW9p6Z2dHYZkLJVnL5AfF
Jyk2K2dRK3h1Pnx7xJ7Dk6UhwLxLntguZ55vKxVshiCRW/Ag7UZyI/kWmu7Ft3IH
K8mXEWs6fDxTkI236PVRhen/Z9QNvvOehNjXS9oJWTesHBWszG9z15YBOpA7DtYz
oM3chrxqejPggu9+X2g5lJR3X2VOz4CSYsoKKUUxSmwyHc322lJO7O/0dPfabXDi
ap/+AT71SDZr3BYheNOSm2vmjE/zehtfLDWMn84Se5OEaqfJ6XnHHfCHvIDy1kBL
N97y1KmljUNfG7kK1laU78dRj9TSHgcY0FDqDMId4tkUZr2U2cK6d9ibU78+uR6u
IkTVHdt7AMy7U6WPGsQmduc91XhxHw1ossUqTULSDxnr8KBD97Xdz05kv1RY/Y28
a0/RjhFUHkceYXK9T9bj6CwZ/fM4xXpTBYjtLihKtAApTr4WGkH3F81p3Gnzqd2U
OgQbrGfCahBYGxLinU1j3+bLhdpxbn88CpL4BdT6qzHlchmViU1RZrsKhrD/Txk6
WYCJkwV+k/Wx0Lf8cLdnQ4ue7f3VxkRWfi57KzIQqxH86Kyka/u/1XhygX0YQn05
3VcxyDE8qya+PJd31NKFrukuYLhGigYhoqmfB6SdfTfEFCQ4MhPIG/3Z6OsLHAAv
MtEuNcWZA6CtCfYfgDcM1uFFrhzyUlTbJ39RxFtg3AXHfXFexVB38wBLO9rirZGz
ql6vOUomsdOW653JRaXEA4OBUfgn59ky9+CxhGKzwL2pVtt+MPa/EnkbQiv3GAs1
FxNGY7XBojIwAhkoxIQXfoCPME/38TIG0hRlPkw2KShQUd/OWiDNrBZIRYU38cKa
oF+L6pcH1fq4W+QoNX2baeI90a+5S56bQ62CJMXB0G+YtlaC278flbKXY/4EPAzp
jKiSoImHiYv3HW/2OYN2fOphjfnMy1G2S3QW6az6XKTjSMBGpZdJmL/mpyhZCsg5
3V/ekhLnWjhv4YttSUKLeW9r7BKtfCLPqHD2rQ/dmFDeWe1f2ZbGpQ+uz5wqXbil
w+zOa9JTwopHnqmLDgOg6iVWdl/7PUA/Q/CxN268autcdVxdf0CqVCeVMWoJlZaf
BjLEq7XpNXWjn2buXCOwqKCXjVMwb1YFpCh+Kto7ebp/XRHcHAularlJvIhoh6Lb
rXg2K0m4GQLI3I5ARJaY/QoLrb9RHtDZ1F8uX7u60w5b9gMo+LRt1Q2H2WX20DIN
TPdefWDXqQ5MgWv5ftESalHFjpBO3QJS6LKkjdZSLfk3ohctXlWgaJhQgJ7wERsE
xpMsTNkdHgfijCnSrbp/hziqT295jnrD8tsPMarszH/CxKwiNEAf3Ll46oJHgMJp
jr/aENRkJw+m6BPDe1NFBnVe2Ir0Z/0y6mLgPGpRSEndd0Qj/kCmOLoHIhx8w5I2
9eUUbKJ5Nv8ZWV8Tl18t/dRVAwYe00cRiUjpBQ5n+db7yOsF9by4CiLgd1NXJd1P
FgfSMiLHsScXhYKpz7wTAHmHaW39h3HTm+y2N/FiXSXg2f2dCtNiP6NfTMYR01Wm
FS7+NO63iuPokGxz8XY8GNVLnOaGL5Ts31pMf7bLkap/0oH+gYk8v73v2BKFMrmn
QaNfjpTh5z0aCqKyZXHPAxXpYe3H1Sgsh+D+CnnfNGEKMYrf8usuzgDgmAJ+nDL6
Bwj0ELX3Ri08bKd7dfR9jWOOAQxNa0mCUyKTZE4eWjGMO51OoBHJq+r576GLrs1g
oKwxFB5/wei9vM31nXtCdoqddfOwI7fFyLBxY2s8g7VPnzQvMyB6r8dpEimYrCFL
ZC2JaEOhCXmkcnbWKxNj7ONhsjsJXForhcR7qT0nZEBAf/vAjmVw3F3ZCuO6cSEC
Xomi8MbbkWVwO1noXKvD2bf0lKkAU94FfOO/n6SR2sB/FaEXsToB/Flszmv2U+mn
RT1fwjh8+i5JIkeaDz+qKbUL+ioyYhBG/D223DKnjrX9xe3jkY0JKXSlP7XpwYp0
ggxYtmqzKA0A3G+CUfw6qNEVULhq7RUTDXF4K3HXL5wZ/y5eXXlJg+3jZUgnrUf1
e8u0hn8fU0Dq/8E6EIotjld8iBtajiMB9ciA6BVOchfA56RiwWkEp822yXKAUnnE
ZmQs9luaSx6dOC0idj/8MsU4PdtCAdOrecbs4hSK5TWF/664rUZjbpIfaZp1Rt+6
kx97GtkTJOWInsh5GaYF+nZKO3+A8PzNVboBExTBTUAqXuCCWDUcgrAWlXh4Kbx9
rH7EC2/jDtOje4qsxDdiN0qcFR08/U2AoVCPOMMQeZ9yNyTXll5mbf4AW7RWd3tz
sk+uJ5jt5b9doJFtOnFdqA0gh1q3YEWGsP94jiTSnOyqHsA2Qy75UIXHMjdBZf1y
wMMVNfEka73hwqOP12MKqWcQJrqT2uMXQy0g3YSD8Iwv8r/J6ALwXtKlEh1+ch6K
l7InLza/cSbQ/fE1qBut7ZqOIL0zkzdR3DBU6Gde1+ly8OzzblAx/aiTXhDIuQG5
3KWqhkbYAa2GiJL4SW4p/cxYMY7/NQfw49rRG10tFi8KDiSSd/ZI61q2IEj6nOfr
X5zu13tD+yNl2b6w5qwQklGm3PezdWL1uvGUfDIVX4iBuIrg3GHCQ/VOOO4j/ABP
Oa9bjqQWp9HbKt43KesHOkTLWgSLlEt7JkZYZPxUwNd8x2yWdxnvicopR9bl4XAy
zr3oXGk1A7voWU90XZK1+h1d9eUUyai+qFO26LgiRTSTYdBWR8Ay2jNlTd9wuoge
TUPV5r9ra2/DroH1UTGYvVXgK/wLXK1VZTEQXdTOKTwI4cOEidvi9z/Wd23Ao6jO
55BFr70kRt2B8ADt7PErFo9vZAtfHddxKmbAZrkDXIdz0QDAyFlzAjgqpgEjxbRp
Q4PDXHPBdrHvUZ3hsy3ZPTFfF+G2s8Pl3tz6uyNjX4zx9IzZQlkngDuG6SqKL3LF
njP+qBvTqCpD0O01FMqzNns8D4KPIossjlmZdP3eyw6WzvO8igpwI5WOzE1UesPW
HDAkjBz7ZAeYQaX8XbBfn4MllKhgsds07JvISFFUrfwgUlz9J18xNDWeE+2yKdcl
DJ8nEo2t3OfhyKqRoot6ivBcWe/EzjOUTKxTDj56y1o4i28szrNP+AMie5jybje5
RFWvvzM754PHkz5DgY7u5kLnB7rHD0uWTSic/vtfxANVlazyCr2zqgQ4y0Hw0+bU
3LV94C/geL8/5dRtFAftVDuqechp5I7KKkuGCW5/qF2WzcJNUN+Jn63t1rRwtkYd
jewT0ZDzJpic9WzK7IMoQfQhlF4Eo/L8OXffiBRdX6X48lpWpTVp+d+FMo6r98Ar
qLVDn28aM0m5kHM6t2vhXqq2cnSCaKokOei5nR0+ocdaPtLV9d0QRxry+zaJvcnM
yx1FJUhekl+WxuaGiUA0CWFYjWSuwH2UMo+uOpLV4dvNZEay5jVU+x3ANcscT7xP
7frySDIf4JOrbi0kmSyyqw1thBdzSme7ISyk3U0EjJgZi3ETntiM2rcyxzZRd5ce
qf7KP8i37CZA65u5fXItrOVf5QTLH/qvDkmrlHi7rzxJQTOO7ty0SYigYxJQzdTg
SJ1d8SxZ9qeP2A4+V7DmcT8jpFnPFqcn7r77dqgs30yBasYJHmERiNKLf628S/pp
gOFwptmqvGE45uk/IRhZ3VLae2u8j4/mWoUIK1gelTaQu5eBxpya3ncafwScmQau
rZuQSYJDJYvkyOGDPg8VmyZGIfidOa1NHMlCFGUOJBvv8XcnyDfiJYItG9op5+dH
iShjYBP+vtwlN7hqgE8fiU/sf8+1SRIxAtucjdH9HP+ihcNRwY2+vmjcZ90KKYTa
h9XffrAVi0312aIVkzvjH5TXoLGQROC2TkfJer/dDCPaWs8W+0UWpUW3L532VV5w
JMqoBJesX7U8/PgbREGajgjVD3oTUGuChO9ddVFCf3thJU1drVxCSIXrigU2nQaX
vARYcoKttWbnUz0sPwh0gSq6lhgVNf+MhkQURmM/mudX4zwEVYFkXr8rWVZTYhwr
JeTu8SsBplHckd5MqAHfzJNn04P/bYvq252j6Bq8FAkMRG1PMDVt6dyhBWCLEQMZ
xhAzmG4+K00DQO/SrKLs7+2ag9G6lfwFqudLhr+ZYKpWxmkpHAS9Ck13ypvImafQ
zZpM3wBOnZKmQFfklnRoub+H0+IgHCE/mOLE/O4Xlr9i4QDlvMFm9ht+5per2a2k
XfsBlbjG1vU1h3N3tmbEykc6WB2wCwUst355AjhPd2c9HCJnPMBKjVEK+q8w/xnB
EfeKcfXKj4UcOZfQRpn5IdBT6gsfO2eoQKLJePdHXz/ICSwG0ksd8nMHzdj7HbFO
pO5P7td1AB8Sg9elu+sUrleg93Ljzu8qoQBWQBeacIT2tkq4Z5V+K7yXpYS1deNk
EBk2z8nWO57pIh/2JTh60YzeGy9+SKqDjjyeJ9TqzPVwY59MUFdZSslaj+frdlei
JCovULLIwY0sVXcmF4cRd4MOg5PeuKwD+fjAavbsEJbXyioV9GWfelKyEUQxR5e7
OgE5ZdB0Dlg9Q7WMiZR0kqBjBi5+dkk+aP6RG3E2aYiwmhNj1o/fJmVcminelB83
2QWXoWALEpta4/xa6wfIwXZ0e/bNnKHgWUMQJz6yF7lXuE4oZ9wSMcQDbnQDpvSo
2cfUNkoZS1aIP96oqj2e13Bu5zDq+ry5rBvN+QMbJKf2aY6k/41nl0ZjF9IniZIm
`pragma protect end_protected
