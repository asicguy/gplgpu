// Copyright (C) 1991-2010 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus II"
// VERSION "Version 10.0 Build 262 08/18/2010 Service Pack 1 SJ Full Version"

// DATE "02/05/2011 12:53:01"

// 
// Device: Altera EP2AGX95EF35I3 Package FBGA1152
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module ddr3_int (
	local_address,
	local_write_req,
	local_read_req,
	local_burstbegin,
	local_wdata,
	local_be,
	local_size,
	global_reset_n,
	pll_ref_clk,
	soft_reset_n,
	local_ready,
	local_rdata,
	local_rdata_valid,
	reset_request_n,
	mem_odt,
	mem_cs_n,
	mem_cke,
	mem_addr,
	mem_ba,
	mem_ras_n,
	mem_cas_n,
	mem_we_n,
	mem_dm,
	local_refresh_ack,
	local_wdata_req,
	local_init_done,
	reset_phy_clk_n,
	mem_reset_n,
	dll_reference_clk,
	dqs_delay_ctrl_export,
	phy_clk,
	aux_full_rate_clk,
	aux_half_rate_clk,
	mem_clk,
	mem_clk_n,
	mem_dq,
	mem_dqs,
	mem_dqsn)/* synthesis synthesis_greybox=0 */;
input 	[24:0] local_address;
input 	local_write_req;
input 	local_read_req;
input 	local_burstbegin;
input 	[127:0] local_wdata;
input 	[15:0] local_be;
input 	[6:0] local_size;
input 	global_reset_n;
input 	pll_ref_clk;
input 	soft_reset_n;
output 	local_ready;
output 	[127:0] local_rdata;
output 	local_rdata_valid;
output 	reset_request_n;
output 	[0:0] mem_odt;
output 	[0:0] mem_cs_n;
output 	[0:0] mem_cke;
output 	[13:0] mem_addr;
output 	[2:0] mem_ba;
output 	mem_ras_n;
output 	mem_cas_n;
output 	mem_we_n;
output 	[3:0] mem_dm;
output 	local_refresh_ack;
output 	local_wdata_req;
output 	local_init_done;
output 	reset_phy_clk_n;
output 	mem_reset_n;
output 	dll_reference_clk;
output 	[5:0] dqs_delay_ctrl_export;
output 	phy_clk;
output 	aux_full_rate_clk;
output 	aux_half_rate_clk;
inout 	[0:0] mem_clk;
inout 	[0:0] mem_clk_n;
inout 	[31:0] mem_dq;
inout 	[3:0] mem_dqs;
inout 	[3:0] mem_dqsn;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[64] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[1] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[65] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[2] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[66] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[3] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[67] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[4] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[68] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[5] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[69] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[6] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[70] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[7] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[71] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[16] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[80] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[17] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[81] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[18] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[82] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[19] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[83] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[20] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[84] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[21] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[85] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[22] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[86] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[23] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[87] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[32] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[96] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[33] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[97] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[34] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[98] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[35] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[99] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[36] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[100] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[37] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[101] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[38] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[102] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[39] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[103] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[48] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[112] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[49] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[113] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[50] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[114] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[51] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[115] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[52] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[116] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[53] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[117] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[54] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[118] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[55] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[119] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[8] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[72] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[9] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[73] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[10] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[74] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[11] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[75] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[12] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[76] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[13] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[77] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[14] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[78] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[15] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[79] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[24] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[88] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[25] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[89] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[26] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[90] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[27] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[91] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[28] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[92] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[29] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[93] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[30] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[94] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[31] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[95] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[40] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[104] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[41] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[105] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[42] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[106] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[43] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[107] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[44] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[108] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[45] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[109] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[46] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[110] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[47] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[111] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[56] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[120] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[57] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[121] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[58] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[122] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[59] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[123] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[60] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[124] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[61] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[125] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[62] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[126] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[63] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[127] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|half_rate.pll|altpll_component|auto_generated|clk[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|half_rate.pll|altpll_component|auto_generated|clk[1] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|gen_odt.odt[0].odt_struct|half_rate.addr_pin|auto_generated|dataout[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|cs_n[0].cs_n_struct|half_rate.addr_pin|auto_generated|dataout[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|cke[0].cke_struct|half_rate.addr_pin|auto_generated|dataout[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[0].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[1].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[2].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[3].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[4].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[5].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[6].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[7].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[8].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[9].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[10].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[11].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[12].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[13].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|ba[0].ba_struct|half_rate.addr_pin|auto_generated|dataout[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|ba[1].ba_struct|half_rate.addr_pin|auto_generated|dataout[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|ba[2].ba_struct|half_rate.addr_pin|auto_generated|dataout[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|ras_n_struct|half_rate.addr_pin|auto_generated|dataout[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|cas_n_struct|half_rate.addr_pin|auto_generated|dataout[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|we_n_struct|half_rate.addr_pin|auto_generated|dataout[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|ddr3_rst.ddr3_rst_struct|half_rate.addr_pin|auto_generated|dataout[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|dqs_delay_ctrl[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|dqs_delay_ctrl[1] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|dqs_delay_ctrl[2] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|dqs_delay_ctrl[3] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|dqs_delay_ctrl[4] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|dqs_delay_ctrl[5] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|wire_output_dq_0_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|wire_output_dq_0_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|wire_output_dq_0_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|wire_output_dq_0_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|mem_clk_buf_in[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|mem_clk_n_buf_in[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|wire_bidir_dq_0_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|wire_bidir_dq_1_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|wire_bidir_dq_2_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|wire_bidir_dq_3_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|wire_bidir_dq_4_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|wire_bidir_dq_5_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|wire_bidir_dq_6_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|wire_bidir_dq_7_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|wire_bidir_dq_0_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|wire_bidir_dq_1_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|wire_bidir_dq_2_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|wire_bidir_dq_3_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|wire_bidir_dq_4_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|wire_bidir_dq_5_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|wire_bidir_dq_6_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|wire_bidir_dq_7_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|wire_bidir_dq_0_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|wire_bidir_dq_1_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|wire_bidir_dq_2_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|wire_bidir_dq_3_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|wire_bidir_dq_4_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|wire_bidir_dq_5_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|wire_bidir_dq_6_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|wire_bidir_dq_7_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|wire_bidir_dq_0_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|wire_bidir_dq_1_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|wire_bidir_dq_2_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|wire_bidir_dq_3_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|wire_bidir_dq_4_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|wire_bidir_dq_5_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|wire_bidir_dq_6_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|wire_bidir_dq_7_output_ddio_out_inst_dataout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_pseudo_diff_out[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqsn_pseudo_diff_out[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_pseudo_diff_out[1] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqsn_pseudo_diff_out[1] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_pseudo_diff_out[2] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqsn_pseudo_diff_out[2] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_pseudo_diff_out[3] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqsn_pseudo_diff_out[3] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[1] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[2] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[3] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[4] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[5] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[6] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[7] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[8] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[9] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[10] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[11] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[12] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[13] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[14] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[15] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[16] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[17] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[18] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[19] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[20] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[21] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[22] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[23] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[24] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[25] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[26] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[27] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[28] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[29] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[30] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[31] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_buffered[0] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_buffered[1] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_buffered[2] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_buffered[3] ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|fb_clk ;
wire \ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|cmd_gen_inst|ready_out~combout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdv_pipe|ctl_rdata_valid[0]~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|half_rate.pll|altpll_component|auto_generated|locked~combout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|state_machine_inst|int_refresh_ack~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|local_init_done~combout ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|reset_phy_clk_1x_n~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|bidir_dq_0_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|bidir_dq_1_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|bidir_dq_2_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|bidir_dq_3_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|bidir_dq_4_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|bidir_dq_5_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|bidir_dq_6_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|bidir_dq_7_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|bidir_dq_0_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|bidir_dq_1_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|bidir_dq_2_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|bidir_dq_3_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|bidir_dq_4_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|bidir_dq_5_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|bidir_dq_6_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|bidir_dq_7_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|bidir_dq_0_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|bidir_dq_1_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|bidir_dq_2_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|bidir_dq_3_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|bidir_dq_4_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|bidir_dq_5_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|bidir_dq_6_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|bidir_dq_7_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|bidir_dq_0_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|bidir_dq_1_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|bidir_dq_2_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|bidir_dq_3_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|bidir_dq_4_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|bidir_dq_5_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|bidir_dq_6_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|bidir_dq_7_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|dqs_0_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|dqs_0_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|dqs_0_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|dqs_0_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|dqsn_0_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|dqsn_0_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|dqsn_0_oe_ff_inst~q ;
wire \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|dqsn_0_oe_ff_inst~q ;
wire \~GND~combout ;
wire \mem_clk_n[0]~input_o ;
wire \local_size[1]~input_o ;
wire \local_address[0]~input_o ;
wire \local_size[0]~input_o ;
wire \local_size[6]~input_o ;
wire \local_size[5]~input_o ;
wire \local_size[4]~input_o ;
wire \local_size[2]~input_o ;
wire \local_size[3]~input_o ;
wire \local_read_req~input_o ;
wire \local_write_req~input_o ;
wire \local_burstbegin~input_o ;
wire \global_reset_n~input_o ;
wire \pll_ref_clk~input_o ;
wire \soft_reset_n~input_o ;
wire \local_address[8]~input_o ;
wire \local_address[10]~input_o ;
wire \local_address[9]~input_o ;
wire \local_address[23]~input_o ;
wire \local_address[24]~input_o ;
wire \local_address[22]~input_o ;
wire \local_address[20]~input_o ;
wire \local_address[21]~input_o ;
wire \local_address[19]~input_o ;
wire \local_address[17]~input_o ;
wire \local_address[18]~input_o ;
wire \local_address[13]~input_o ;
wire \local_address[11]~input_o ;
wire \local_address[12]~input_o ;
wire \local_address[16]~input_o ;
wire \local_address[14]~input_o ;
wire \local_address[15]~input_o ;
wire \local_address[1]~input_o ;
wire \local_address[2]~input_o ;
wire \local_address[3]~input_o ;
wire \local_address[4]~input_o ;
wire \local_address[5]~input_o ;
wire \local_address[7]~input_o ;
wire \local_address[6]~input_o ;
wire \local_be[4]~input_o ;
wire \local_be[12]~input_o ;
wire \local_be[0]~input_o ;
wire \local_be[8]~input_o ;
wire \local_be[5]~input_o ;
wire \local_be[13]~input_o ;
wire \local_be[1]~input_o ;
wire \local_be[9]~input_o ;
wire \local_be[6]~input_o ;
wire \local_be[14]~input_o ;
wire \local_be[2]~input_o ;
wire \local_be[10]~input_o ;
wire \local_be[7]~input_o ;
wire \local_be[15]~input_o ;
wire \local_be[3]~input_o ;
wire \local_be[11]~input_o ;
wire \local_wdata[96]~input_o ;
wire \local_wdata[32]~input_o ;
wire \local_wdata[64]~input_o ;
wire \local_wdata[0]~input_o ;
wire \local_wdata[97]~input_o ;
wire \local_wdata[33]~input_o ;
wire \local_wdata[65]~input_o ;
wire \local_wdata[1]~input_o ;
wire \local_wdata[98]~input_o ;
wire \local_wdata[34]~input_o ;
wire \local_wdata[66]~input_o ;
wire \local_wdata[2]~input_o ;
wire \local_wdata[99]~input_o ;
wire \local_wdata[35]~input_o ;
wire \local_wdata[67]~input_o ;
wire \local_wdata[3]~input_o ;
wire \local_wdata[100]~input_o ;
wire \local_wdata[36]~input_o ;
wire \local_wdata[68]~input_o ;
wire \local_wdata[4]~input_o ;
wire \local_wdata[101]~input_o ;
wire \local_wdata[37]~input_o ;
wire \local_wdata[69]~input_o ;
wire \local_wdata[5]~input_o ;
wire \local_wdata[102]~input_o ;
wire \local_wdata[38]~input_o ;
wire \local_wdata[70]~input_o ;
wire \local_wdata[6]~input_o ;
wire \local_wdata[103]~input_o ;
wire \local_wdata[39]~input_o ;
wire \local_wdata[71]~input_o ;
wire \local_wdata[7]~input_o ;
wire \local_wdata[104]~input_o ;
wire \local_wdata[40]~input_o ;
wire \local_wdata[72]~input_o ;
wire \local_wdata[8]~input_o ;
wire \local_wdata[105]~input_o ;
wire \local_wdata[41]~input_o ;
wire \local_wdata[73]~input_o ;
wire \local_wdata[9]~input_o ;
wire \local_wdata[106]~input_o ;
wire \local_wdata[42]~input_o ;
wire \local_wdata[74]~input_o ;
wire \local_wdata[10]~input_o ;
wire \local_wdata[107]~input_o ;
wire \local_wdata[43]~input_o ;
wire \local_wdata[75]~input_o ;
wire \local_wdata[11]~input_o ;
wire \local_wdata[108]~input_o ;
wire \local_wdata[44]~input_o ;
wire \local_wdata[76]~input_o ;
wire \local_wdata[12]~input_o ;
wire \local_wdata[109]~input_o ;
wire \local_wdata[45]~input_o ;
wire \local_wdata[77]~input_o ;
wire \local_wdata[13]~input_o ;
wire \local_wdata[110]~input_o ;
wire \local_wdata[46]~input_o ;
wire \local_wdata[78]~input_o ;
wire \local_wdata[14]~input_o ;
wire \local_wdata[111]~input_o ;
wire \local_wdata[47]~input_o ;
wire \local_wdata[79]~input_o ;
wire \local_wdata[15]~input_o ;
wire \local_wdata[112]~input_o ;
wire \local_wdata[48]~input_o ;
wire \local_wdata[80]~input_o ;
wire \local_wdata[16]~input_o ;
wire \local_wdata[113]~input_o ;
wire \local_wdata[49]~input_o ;
wire \local_wdata[81]~input_o ;
wire \local_wdata[17]~input_o ;
wire \local_wdata[114]~input_o ;
wire \local_wdata[50]~input_o ;
wire \local_wdata[82]~input_o ;
wire \local_wdata[18]~input_o ;
wire \local_wdata[115]~input_o ;
wire \local_wdata[51]~input_o ;
wire \local_wdata[83]~input_o ;
wire \local_wdata[19]~input_o ;
wire \local_wdata[116]~input_o ;
wire \local_wdata[52]~input_o ;
wire \local_wdata[84]~input_o ;
wire \local_wdata[20]~input_o ;
wire \local_wdata[117]~input_o ;
wire \local_wdata[53]~input_o ;
wire \local_wdata[85]~input_o ;
wire \local_wdata[21]~input_o ;
wire \local_wdata[118]~input_o ;
wire \local_wdata[54]~input_o ;
wire \local_wdata[86]~input_o ;
wire \local_wdata[22]~input_o ;
wire \local_wdata[119]~input_o ;
wire \local_wdata[55]~input_o ;
wire \local_wdata[87]~input_o ;
wire \local_wdata[23]~input_o ;
wire \local_wdata[120]~input_o ;
wire \local_wdata[56]~input_o ;
wire \local_wdata[88]~input_o ;
wire \local_wdata[24]~input_o ;
wire \local_wdata[121]~input_o ;
wire \local_wdata[57]~input_o ;
wire \local_wdata[89]~input_o ;
wire \local_wdata[25]~input_o ;
wire \local_wdata[122]~input_o ;
wire \local_wdata[58]~input_o ;
wire \local_wdata[90]~input_o ;
wire \local_wdata[26]~input_o ;
wire \local_wdata[123]~input_o ;
wire \local_wdata[59]~input_o ;
wire \local_wdata[91]~input_o ;
wire \local_wdata[27]~input_o ;
wire \local_wdata[124]~input_o ;
wire \local_wdata[60]~input_o ;
wire \local_wdata[92]~input_o ;
wire \local_wdata[28]~input_o ;
wire \local_wdata[125]~input_o ;
wire \local_wdata[61]~input_o ;
wire \local_wdata[93]~input_o ;
wire \local_wdata[29]~input_o ;
wire \local_wdata[126]~input_o ;
wire \local_wdata[62]~input_o ;
wire \local_wdata[94]~input_o ;
wire \local_wdata[30]~input_o ;
wire \local_wdata[127]~input_o ;
wire \local_wdata[63]~input_o ;
wire \local_wdata[95]~input_o ;
wire \local_wdata[31]~input_o ;


ddr3_int_ddr3_int_controller_phy ddr3_int_controller_phy_inst(
	.q_b_0(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[0] ),
	.q_b_64(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[64] ),
	.q_b_1(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[1] ),
	.q_b_65(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[65] ),
	.q_b_2(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[2] ),
	.q_b_66(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[66] ),
	.q_b_3(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[3] ),
	.q_b_67(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[67] ),
	.q_b_4(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[4] ),
	.q_b_68(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[68] ),
	.q_b_5(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[5] ),
	.q_b_69(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[69] ),
	.q_b_6(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[6] ),
	.q_b_70(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[70] ),
	.q_b_7(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[7] ),
	.q_b_71(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[71] ),
	.q_b_16(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[16] ),
	.q_b_80(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[80] ),
	.q_b_17(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[17] ),
	.q_b_81(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[81] ),
	.q_b_18(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[18] ),
	.q_b_82(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[82] ),
	.q_b_19(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[19] ),
	.q_b_83(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[83] ),
	.q_b_20(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[20] ),
	.q_b_84(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[84] ),
	.q_b_21(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[21] ),
	.q_b_85(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[85] ),
	.q_b_22(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[22] ),
	.q_b_86(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[86] ),
	.q_b_23(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[23] ),
	.q_b_87(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[87] ),
	.q_b_32(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[32] ),
	.q_b_96(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[96] ),
	.q_b_33(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[33] ),
	.q_b_97(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[97] ),
	.q_b_34(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[34] ),
	.q_b_98(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[98] ),
	.q_b_35(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[35] ),
	.q_b_99(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[99] ),
	.q_b_36(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[36] ),
	.q_b_100(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[100] ),
	.q_b_37(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[37] ),
	.q_b_101(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[101] ),
	.q_b_38(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[38] ),
	.q_b_102(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[102] ),
	.q_b_39(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[39] ),
	.q_b_103(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[103] ),
	.q_b_48(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[48] ),
	.q_b_112(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[112] ),
	.q_b_49(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[49] ),
	.q_b_113(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[113] ),
	.q_b_50(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[50] ),
	.q_b_114(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[114] ),
	.q_b_51(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[51] ),
	.q_b_115(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[115] ),
	.q_b_52(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[52] ),
	.q_b_116(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[116] ),
	.q_b_53(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[53] ),
	.q_b_117(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[117] ),
	.q_b_54(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[54] ),
	.q_b_118(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[118] ),
	.q_b_55(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[55] ),
	.q_b_119(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[119] ),
	.q_b_8(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[8] ),
	.q_b_72(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[72] ),
	.q_b_9(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[9] ),
	.q_b_73(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[73] ),
	.q_b_10(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[10] ),
	.q_b_74(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[74] ),
	.q_b_11(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[11] ),
	.q_b_75(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[75] ),
	.q_b_12(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[12] ),
	.q_b_76(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[76] ),
	.q_b_13(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[13] ),
	.q_b_77(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[77] ),
	.q_b_14(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[14] ),
	.q_b_78(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[78] ),
	.q_b_15(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[15] ),
	.q_b_79(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[79] ),
	.q_b_24(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[24] ),
	.q_b_88(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[88] ),
	.q_b_25(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[25] ),
	.q_b_89(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[89] ),
	.q_b_26(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[26] ),
	.q_b_90(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[90] ),
	.q_b_27(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[27] ),
	.q_b_91(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[91] ),
	.q_b_28(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[28] ),
	.q_b_92(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[92] ),
	.q_b_29(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[29] ),
	.q_b_93(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[93] ),
	.q_b_30(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[30] ),
	.q_b_94(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[94] ),
	.q_b_31(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[31] ),
	.q_b_95(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[95] ),
	.q_b_40(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[40] ),
	.q_b_104(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[104] ),
	.q_b_41(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[41] ),
	.q_b_105(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[105] ),
	.q_b_42(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[42] ),
	.q_b_106(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[106] ),
	.q_b_43(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[43] ),
	.q_b_107(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[107] ),
	.q_b_44(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[44] ),
	.q_b_108(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[108] ),
	.q_b_45(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[45] ),
	.q_b_109(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[109] ),
	.q_b_46(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[46] ),
	.q_b_110(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[110] ),
	.q_b_47(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[47] ),
	.q_b_111(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[111] ),
	.q_b_56(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[56] ),
	.q_b_120(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[120] ),
	.q_b_57(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[57] ),
	.q_b_121(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[121] ),
	.q_b_58(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[58] ),
	.q_b_122(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[122] ),
	.q_b_59(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[59] ),
	.q_b_123(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[123] ),
	.q_b_60(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[60] ),
	.q_b_124(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[124] ),
	.q_b_61(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[61] ),
	.q_b_125(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[125] ),
	.q_b_62(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[62] ),
	.q_b_126(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[126] ),
	.q_b_63(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[63] ),
	.q_b_127(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[127] ),
	.clk_0(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|half_rate.pll|altpll_component|auto_generated|clk[0] ),
	.clk_1(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|half_rate.pll|altpll_component|auto_generated|clk[1] ),
	.dataout_0(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|gen_odt.odt[0].odt_struct|half_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_01(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|cs_n[0].cs_n_struct|half_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_02(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|cke[0].cke_struct|half_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_03(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[0].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_04(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[1].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_05(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[2].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_06(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[3].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_07(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[4].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_08(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[5].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_09(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[6].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_010(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[7].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_011(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[8].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_012(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[9].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_013(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[10].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_014(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[11].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_015(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[12].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_016(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[13].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_017(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|ba[0].ba_struct|half_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_018(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|ba[1].ba_struct|half_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_019(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|ba[2].ba_struct|half_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_020(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|ras_n_struct|half_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_021(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|cas_n_struct|half_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_022(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|we_n_struct|half_rate.addr_pin|auto_generated|dataout[0] ),
	.dataout_023(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|ddr3_rst.ddr3_rst_struct|half_rate.addr_pin|auto_generated|dataout[0] ),
	.dqs_delay_ctrl_0(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|dqs_delay_ctrl[0] ),
	.dqs_delay_ctrl_1(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|dqs_delay_ctrl[1] ),
	.dqs_delay_ctrl_2(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|dqs_delay_ctrl[2] ),
	.dqs_delay_ctrl_3(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|dqs_delay_ctrl[3] ),
	.dqs_delay_ctrl_4(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|dqs_delay_ctrl[4] ),
	.dqs_delay_ctrl_5(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|dqs_delay_ctrl[5] ),
	.wire_output_dq_0_output_ddio_out_inst_dataout(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|wire_output_dq_0_output_ddio_out_inst_dataout ),
	.wire_output_dq_0_output_ddio_out_inst_dataout1(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|wire_output_dq_0_output_ddio_out_inst_dataout ),
	.wire_output_dq_0_output_ddio_out_inst_dataout2(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|wire_output_dq_0_output_ddio_out_inst_dataout ),
	.wire_output_dq_0_output_ddio_out_inst_dataout3(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|wire_output_dq_0_output_ddio_out_inst_dataout ),
	.mem_clk_buf_in_0(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|mem_clk_buf_in[0] ),
	.mem_clk_n_buf_in_0(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|mem_clk_n_buf_in[0] ),
	.wire_bidir_dq_0_output_ddio_out_inst_dataout(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|wire_bidir_dq_0_output_ddio_out_inst_dataout ),
	.wire_bidir_dq_1_output_ddio_out_inst_dataout(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|wire_bidir_dq_1_output_ddio_out_inst_dataout ),
	.wire_bidir_dq_2_output_ddio_out_inst_dataout(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|wire_bidir_dq_2_output_ddio_out_inst_dataout ),
	.wire_bidir_dq_3_output_ddio_out_inst_dataout(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|wire_bidir_dq_3_output_ddio_out_inst_dataout ),
	.wire_bidir_dq_4_output_ddio_out_inst_dataout(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|wire_bidir_dq_4_output_ddio_out_inst_dataout ),
	.wire_bidir_dq_5_output_ddio_out_inst_dataout(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|wire_bidir_dq_5_output_ddio_out_inst_dataout ),
	.wire_bidir_dq_6_output_ddio_out_inst_dataout(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|wire_bidir_dq_6_output_ddio_out_inst_dataout ),
	.wire_bidir_dq_7_output_ddio_out_inst_dataout(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|wire_bidir_dq_7_output_ddio_out_inst_dataout ),
	.wire_bidir_dq_0_output_ddio_out_inst_dataout1(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|wire_bidir_dq_0_output_ddio_out_inst_dataout ),
	.wire_bidir_dq_1_output_ddio_out_inst_dataout1(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|wire_bidir_dq_1_output_ddio_out_inst_dataout ),
	.wire_bidir_dq_2_output_ddio_out_inst_dataout1(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|wire_bidir_dq_2_output_ddio_out_inst_dataout ),
	.wire_bidir_dq_3_output_ddio_out_inst_dataout1(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|wire_bidir_dq_3_output_ddio_out_inst_dataout ),
	.wire_bidir_dq_4_output_ddio_out_inst_dataout1(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|wire_bidir_dq_4_output_ddio_out_inst_dataout ),
	.wire_bidir_dq_5_output_ddio_out_inst_dataout1(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|wire_bidir_dq_5_output_ddio_out_inst_dataout ),
	.wire_bidir_dq_6_output_ddio_out_inst_dataout1(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|wire_bidir_dq_6_output_ddio_out_inst_dataout ),
	.wire_bidir_dq_7_output_ddio_out_inst_dataout1(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|wire_bidir_dq_7_output_ddio_out_inst_dataout ),
	.wire_bidir_dq_0_output_ddio_out_inst_dataout2(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|wire_bidir_dq_0_output_ddio_out_inst_dataout ),
	.wire_bidir_dq_1_output_ddio_out_inst_dataout2(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|wire_bidir_dq_1_output_ddio_out_inst_dataout ),
	.wire_bidir_dq_2_output_ddio_out_inst_dataout2(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|wire_bidir_dq_2_output_ddio_out_inst_dataout ),
	.wire_bidir_dq_3_output_ddio_out_inst_dataout2(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|wire_bidir_dq_3_output_ddio_out_inst_dataout ),
	.wire_bidir_dq_4_output_ddio_out_inst_dataout2(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|wire_bidir_dq_4_output_ddio_out_inst_dataout ),
	.wire_bidir_dq_5_output_ddio_out_inst_dataout2(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|wire_bidir_dq_5_output_ddio_out_inst_dataout ),
	.wire_bidir_dq_6_output_ddio_out_inst_dataout2(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|wire_bidir_dq_6_output_ddio_out_inst_dataout ),
	.wire_bidir_dq_7_output_ddio_out_inst_dataout2(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|wire_bidir_dq_7_output_ddio_out_inst_dataout ),
	.wire_bidir_dq_0_output_ddio_out_inst_dataout3(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|wire_bidir_dq_0_output_ddio_out_inst_dataout ),
	.wire_bidir_dq_1_output_ddio_out_inst_dataout3(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|wire_bidir_dq_1_output_ddio_out_inst_dataout ),
	.wire_bidir_dq_2_output_ddio_out_inst_dataout3(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|wire_bidir_dq_2_output_ddio_out_inst_dataout ),
	.wire_bidir_dq_3_output_ddio_out_inst_dataout3(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|wire_bidir_dq_3_output_ddio_out_inst_dataout ),
	.wire_bidir_dq_4_output_ddio_out_inst_dataout3(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|wire_bidir_dq_4_output_ddio_out_inst_dataout ),
	.wire_bidir_dq_5_output_ddio_out_inst_dataout3(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|wire_bidir_dq_5_output_ddio_out_inst_dataout ),
	.wire_bidir_dq_6_output_ddio_out_inst_dataout3(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|wire_bidir_dq_6_output_ddio_out_inst_dataout ),
	.wire_bidir_dq_7_output_ddio_out_inst_dataout3(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|wire_bidir_dq_7_output_ddio_out_inst_dataout ),
	.dqs_pseudo_diff_out_0(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_pseudo_diff_out[0] ),
	.dqsn_pseudo_diff_out_0(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqsn_pseudo_diff_out[0] ),
	.dqs_pseudo_diff_out_1(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_pseudo_diff_out[1] ),
	.dqsn_pseudo_diff_out_1(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqsn_pseudo_diff_out[1] ),
	.dqs_pseudo_diff_out_2(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_pseudo_diff_out[2] ),
	.dqsn_pseudo_diff_out_2(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqsn_pseudo_diff_out[2] ),
	.dqs_pseudo_diff_out_3(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_pseudo_diff_out[3] ),
	.dqsn_pseudo_diff_out_3(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqsn_pseudo_diff_out[3] ),
	.dq_datain_0(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[0] ),
	.dq_datain_1(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[1] ),
	.dq_datain_2(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[2] ),
	.dq_datain_3(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[3] ),
	.dq_datain_4(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[4] ),
	.dq_datain_5(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[5] ),
	.dq_datain_6(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[6] ),
	.dq_datain_7(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[7] ),
	.dq_datain_8(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[8] ),
	.dq_datain_9(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[9] ),
	.dq_datain_10(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[10] ),
	.dq_datain_11(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[11] ),
	.dq_datain_12(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[12] ),
	.dq_datain_13(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[13] ),
	.dq_datain_14(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[14] ),
	.dq_datain_15(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[15] ),
	.dq_datain_16(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[16] ),
	.dq_datain_17(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[17] ),
	.dq_datain_18(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[18] ),
	.dq_datain_19(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[19] ),
	.dq_datain_20(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[20] ),
	.dq_datain_21(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[21] ),
	.dq_datain_22(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[22] ),
	.dq_datain_23(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[23] ),
	.dq_datain_24(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[24] ),
	.dq_datain_25(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[25] ),
	.dq_datain_26(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[26] ),
	.dq_datain_27(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[27] ),
	.dq_datain_28(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[28] ),
	.dq_datain_29(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[29] ),
	.dq_datain_30(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[30] ),
	.dq_datain_31(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[31] ),
	.dqs_buffered_0(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_buffered[0] ),
	.dqs_buffered_1(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_buffered[1] ),
	.dqs_buffered_2(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_buffered[2] ),
	.dqs_buffered_3(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_buffered[3] ),
	.fb_clk(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|fb_clk ),
	.ready_out(\ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|cmd_gen_inst|ready_out~combout ),
	.ctl_rdata_valid_0(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdv_pipe|ctl_rdata_valid[0]~q ),
	.reset_request_n(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|half_rate.pll|altpll_component|auto_generated|locked~combout ),
	.int_refresh_ack(\ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|state_machine_inst|int_refresh_ack~q ),
	.local_init_done(\ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|local_init_done~combout ),
	.reset_phy_clk_1x_n(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|reset_phy_clk_1x_n~q ),
	.bidir_dq_0_oe_ff_inst(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|bidir_dq_0_oe_ff_inst~q ),
	.bidir_dq_1_oe_ff_inst(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|bidir_dq_1_oe_ff_inst~q ),
	.bidir_dq_2_oe_ff_inst(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|bidir_dq_2_oe_ff_inst~q ),
	.bidir_dq_3_oe_ff_inst(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|bidir_dq_3_oe_ff_inst~q ),
	.bidir_dq_4_oe_ff_inst(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|bidir_dq_4_oe_ff_inst~q ),
	.bidir_dq_5_oe_ff_inst(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|bidir_dq_5_oe_ff_inst~q ),
	.bidir_dq_6_oe_ff_inst(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|bidir_dq_6_oe_ff_inst~q ),
	.bidir_dq_7_oe_ff_inst(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|bidir_dq_7_oe_ff_inst~q ),
	.bidir_dq_0_oe_ff_inst1(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|bidir_dq_0_oe_ff_inst~q ),
	.bidir_dq_1_oe_ff_inst1(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|bidir_dq_1_oe_ff_inst~q ),
	.bidir_dq_2_oe_ff_inst1(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|bidir_dq_2_oe_ff_inst~q ),
	.bidir_dq_3_oe_ff_inst1(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|bidir_dq_3_oe_ff_inst~q ),
	.bidir_dq_4_oe_ff_inst1(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|bidir_dq_4_oe_ff_inst~q ),
	.bidir_dq_5_oe_ff_inst1(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|bidir_dq_5_oe_ff_inst~q ),
	.bidir_dq_6_oe_ff_inst1(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|bidir_dq_6_oe_ff_inst~q ),
	.bidir_dq_7_oe_ff_inst1(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|bidir_dq_7_oe_ff_inst~q ),
	.bidir_dq_0_oe_ff_inst2(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|bidir_dq_0_oe_ff_inst~q ),
	.bidir_dq_1_oe_ff_inst2(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|bidir_dq_1_oe_ff_inst~q ),
	.bidir_dq_2_oe_ff_inst2(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|bidir_dq_2_oe_ff_inst~q ),
	.bidir_dq_3_oe_ff_inst2(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|bidir_dq_3_oe_ff_inst~q ),
	.bidir_dq_4_oe_ff_inst2(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|bidir_dq_4_oe_ff_inst~q ),
	.bidir_dq_5_oe_ff_inst2(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|bidir_dq_5_oe_ff_inst~q ),
	.bidir_dq_6_oe_ff_inst2(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|bidir_dq_6_oe_ff_inst~q ),
	.bidir_dq_7_oe_ff_inst2(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|bidir_dq_7_oe_ff_inst~q ),
	.bidir_dq_0_oe_ff_inst3(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|bidir_dq_0_oe_ff_inst~q ),
	.bidir_dq_1_oe_ff_inst3(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|bidir_dq_1_oe_ff_inst~q ),
	.bidir_dq_2_oe_ff_inst3(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|bidir_dq_2_oe_ff_inst~q ),
	.bidir_dq_3_oe_ff_inst3(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|bidir_dq_3_oe_ff_inst~q ),
	.bidir_dq_4_oe_ff_inst3(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|bidir_dq_4_oe_ff_inst~q ),
	.bidir_dq_5_oe_ff_inst3(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|bidir_dq_5_oe_ff_inst~q ),
	.bidir_dq_6_oe_ff_inst3(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|bidir_dq_6_oe_ff_inst~q ),
	.bidir_dq_7_oe_ff_inst3(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|bidir_dq_7_oe_ff_inst~q ),
	.dqs_0_oe_ff_inst(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|dqs_0_oe_ff_inst~q ),
	.dqs_0_oe_ff_inst1(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|dqs_0_oe_ff_inst~q ),
	.dqs_0_oe_ff_inst2(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|dqs_0_oe_ff_inst~q ),
	.dqs_0_oe_ff_inst3(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|dqs_0_oe_ff_inst~q ),
	.dqsn_0_oe_ff_inst(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|dqsn_0_oe_ff_inst~q ),
	.dqsn_0_oe_ff_inst1(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|dqsn_0_oe_ff_inst~q ),
	.dqsn_0_oe_ff_inst2(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|dqsn_0_oe_ff_inst~q ),
	.dqsn_0_oe_ff_inst3(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|dqsn_0_oe_ff_inst~q ),
	.GND_port(\~GND~combout ),
	.local_size_1(\local_size[1]~input_o ),
	.local_address_0(\local_address[0]~input_o ),
	.local_size_0(\local_size[0]~input_o ),
	.local_size_6(\local_size[6]~input_o ),
	.local_size_5(\local_size[5]~input_o ),
	.local_size_4(\local_size[4]~input_o ),
	.local_size_2(\local_size[2]~input_o ),
	.local_size_3(\local_size[3]~input_o ),
	.local_read_req(\local_read_req~input_o ),
	.local_write_req(\local_write_req~input_o ),
	.local_burstbegin(\local_burstbegin~input_o ),
	.global_reset_n(\global_reset_n~input_o ),
	.pll_ref_clk(\pll_ref_clk~input_o ),
	.soft_reset_n(\soft_reset_n~input_o ),
	.local_address_8(\local_address[8]~input_o ),
	.local_address_10(\local_address[10]~input_o ),
	.local_address_9(\local_address[9]~input_o ),
	.local_address_23(\local_address[23]~input_o ),
	.local_address_24(\local_address[24]~input_o ),
	.local_address_22(\local_address[22]~input_o ),
	.local_address_20(\local_address[20]~input_o ),
	.local_address_21(\local_address[21]~input_o ),
	.local_address_19(\local_address[19]~input_o ),
	.local_address_17(\local_address[17]~input_o ),
	.local_address_18(\local_address[18]~input_o ),
	.local_address_13(\local_address[13]~input_o ),
	.local_address_11(\local_address[11]~input_o ),
	.local_address_12(\local_address[12]~input_o ),
	.local_address_16(\local_address[16]~input_o ),
	.local_address_14(\local_address[14]~input_o ),
	.local_address_15(\local_address[15]~input_o ),
	.local_address_1(\local_address[1]~input_o ),
	.local_address_2(\local_address[2]~input_o ),
	.local_address_3(\local_address[3]~input_o ),
	.local_address_4(\local_address[4]~input_o ),
	.local_address_5(\local_address[5]~input_o ),
	.local_address_7(\local_address[7]~input_o ),
	.local_address_6(\local_address[6]~input_o ),
	.local_be_4(\local_be[4]~input_o ),
	.local_be_12(\local_be[12]~input_o ),
	.local_be_0(\local_be[0]~input_o ),
	.local_be_8(\local_be[8]~input_o ),
	.local_be_5(\local_be[5]~input_o ),
	.local_be_13(\local_be[13]~input_o ),
	.local_be_1(\local_be[1]~input_o ),
	.local_be_9(\local_be[9]~input_o ),
	.local_be_6(\local_be[6]~input_o ),
	.local_be_14(\local_be[14]~input_o ),
	.local_be_2(\local_be[2]~input_o ),
	.local_be_10(\local_be[10]~input_o ),
	.local_be_7(\local_be[7]~input_o ),
	.local_be_15(\local_be[15]~input_o ),
	.local_be_3(\local_be[3]~input_o ),
	.local_be_11(\local_be[11]~input_o ),
	.local_wdata_96(\local_wdata[96]~input_o ),
	.local_wdata_32(\local_wdata[32]~input_o ),
	.local_wdata_64(\local_wdata[64]~input_o ),
	.local_wdata_0(\local_wdata[0]~input_o ),
	.local_wdata_97(\local_wdata[97]~input_o ),
	.local_wdata_33(\local_wdata[33]~input_o ),
	.local_wdata_65(\local_wdata[65]~input_o ),
	.local_wdata_1(\local_wdata[1]~input_o ),
	.local_wdata_98(\local_wdata[98]~input_o ),
	.local_wdata_34(\local_wdata[34]~input_o ),
	.local_wdata_66(\local_wdata[66]~input_o ),
	.local_wdata_2(\local_wdata[2]~input_o ),
	.local_wdata_99(\local_wdata[99]~input_o ),
	.local_wdata_35(\local_wdata[35]~input_o ),
	.local_wdata_67(\local_wdata[67]~input_o ),
	.local_wdata_3(\local_wdata[3]~input_o ),
	.local_wdata_100(\local_wdata[100]~input_o ),
	.local_wdata_36(\local_wdata[36]~input_o ),
	.local_wdata_68(\local_wdata[68]~input_o ),
	.local_wdata_4(\local_wdata[4]~input_o ),
	.local_wdata_101(\local_wdata[101]~input_o ),
	.local_wdata_37(\local_wdata[37]~input_o ),
	.local_wdata_69(\local_wdata[69]~input_o ),
	.local_wdata_5(\local_wdata[5]~input_o ),
	.local_wdata_102(\local_wdata[102]~input_o ),
	.local_wdata_38(\local_wdata[38]~input_o ),
	.local_wdata_70(\local_wdata[70]~input_o ),
	.local_wdata_6(\local_wdata[6]~input_o ),
	.local_wdata_103(\local_wdata[103]~input_o ),
	.local_wdata_39(\local_wdata[39]~input_o ),
	.local_wdata_71(\local_wdata[71]~input_o ),
	.local_wdata_7(\local_wdata[7]~input_o ),
	.local_wdata_104(\local_wdata[104]~input_o ),
	.local_wdata_40(\local_wdata[40]~input_o ),
	.local_wdata_72(\local_wdata[72]~input_o ),
	.local_wdata_8(\local_wdata[8]~input_o ),
	.local_wdata_105(\local_wdata[105]~input_o ),
	.local_wdata_41(\local_wdata[41]~input_o ),
	.local_wdata_73(\local_wdata[73]~input_o ),
	.local_wdata_9(\local_wdata[9]~input_o ),
	.local_wdata_106(\local_wdata[106]~input_o ),
	.local_wdata_42(\local_wdata[42]~input_o ),
	.local_wdata_74(\local_wdata[74]~input_o ),
	.local_wdata_10(\local_wdata[10]~input_o ),
	.local_wdata_107(\local_wdata[107]~input_o ),
	.local_wdata_43(\local_wdata[43]~input_o ),
	.local_wdata_75(\local_wdata[75]~input_o ),
	.local_wdata_11(\local_wdata[11]~input_o ),
	.local_wdata_108(\local_wdata[108]~input_o ),
	.local_wdata_44(\local_wdata[44]~input_o ),
	.local_wdata_76(\local_wdata[76]~input_o ),
	.local_wdata_12(\local_wdata[12]~input_o ),
	.local_wdata_109(\local_wdata[109]~input_o ),
	.local_wdata_45(\local_wdata[45]~input_o ),
	.local_wdata_77(\local_wdata[77]~input_o ),
	.local_wdata_13(\local_wdata[13]~input_o ),
	.local_wdata_110(\local_wdata[110]~input_o ),
	.local_wdata_46(\local_wdata[46]~input_o ),
	.local_wdata_78(\local_wdata[78]~input_o ),
	.local_wdata_14(\local_wdata[14]~input_o ),
	.local_wdata_111(\local_wdata[111]~input_o ),
	.local_wdata_47(\local_wdata[47]~input_o ),
	.local_wdata_79(\local_wdata[79]~input_o ),
	.local_wdata_15(\local_wdata[15]~input_o ),
	.local_wdata_112(\local_wdata[112]~input_o ),
	.local_wdata_48(\local_wdata[48]~input_o ),
	.local_wdata_80(\local_wdata[80]~input_o ),
	.local_wdata_16(\local_wdata[16]~input_o ),
	.local_wdata_113(\local_wdata[113]~input_o ),
	.local_wdata_49(\local_wdata[49]~input_o ),
	.local_wdata_81(\local_wdata[81]~input_o ),
	.local_wdata_17(\local_wdata[17]~input_o ),
	.local_wdata_114(\local_wdata[114]~input_o ),
	.local_wdata_50(\local_wdata[50]~input_o ),
	.local_wdata_82(\local_wdata[82]~input_o ),
	.local_wdata_18(\local_wdata[18]~input_o ),
	.local_wdata_115(\local_wdata[115]~input_o ),
	.local_wdata_51(\local_wdata[51]~input_o ),
	.local_wdata_83(\local_wdata[83]~input_o ),
	.local_wdata_19(\local_wdata[19]~input_o ),
	.local_wdata_116(\local_wdata[116]~input_o ),
	.local_wdata_52(\local_wdata[52]~input_o ),
	.local_wdata_84(\local_wdata[84]~input_o ),
	.local_wdata_20(\local_wdata[20]~input_o ),
	.local_wdata_117(\local_wdata[117]~input_o ),
	.local_wdata_53(\local_wdata[53]~input_o ),
	.local_wdata_85(\local_wdata[85]~input_o ),
	.local_wdata_21(\local_wdata[21]~input_o ),
	.local_wdata_118(\local_wdata[118]~input_o ),
	.local_wdata_54(\local_wdata[54]~input_o ),
	.local_wdata_86(\local_wdata[86]~input_o ),
	.local_wdata_22(\local_wdata[22]~input_o ),
	.local_wdata_119(\local_wdata[119]~input_o ),
	.local_wdata_55(\local_wdata[55]~input_o ),
	.local_wdata_87(\local_wdata[87]~input_o ),
	.local_wdata_23(\local_wdata[23]~input_o ),
	.local_wdata_120(\local_wdata[120]~input_o ),
	.local_wdata_56(\local_wdata[56]~input_o ),
	.local_wdata_88(\local_wdata[88]~input_o ),
	.local_wdata_24(\local_wdata[24]~input_o ),
	.local_wdata_121(\local_wdata[121]~input_o ),
	.local_wdata_57(\local_wdata[57]~input_o ),
	.local_wdata_89(\local_wdata[89]~input_o ),
	.local_wdata_25(\local_wdata[25]~input_o ),
	.local_wdata_122(\local_wdata[122]~input_o ),
	.local_wdata_58(\local_wdata[58]~input_o ),
	.local_wdata_90(\local_wdata[90]~input_o ),
	.local_wdata_26(\local_wdata[26]~input_o ),
	.local_wdata_123(\local_wdata[123]~input_o ),
	.local_wdata_59(\local_wdata[59]~input_o ),
	.local_wdata_91(\local_wdata[91]~input_o ),
	.local_wdata_27(\local_wdata[27]~input_o ),
	.local_wdata_124(\local_wdata[124]~input_o ),
	.local_wdata_60(\local_wdata[60]~input_o ),
	.local_wdata_92(\local_wdata[92]~input_o ),
	.local_wdata_28(\local_wdata[28]~input_o ),
	.local_wdata_125(\local_wdata[125]~input_o ),
	.local_wdata_61(\local_wdata[61]~input_o ),
	.local_wdata_93(\local_wdata[93]~input_o ),
	.local_wdata_29(\local_wdata[29]~input_o ),
	.local_wdata_126(\local_wdata[126]~input_o ),
	.local_wdata_62(\local_wdata[62]~input_o ),
	.local_wdata_94(\local_wdata[94]~input_o ),
	.local_wdata_30(\local_wdata[30]~input_o ),
	.local_wdata_127(\local_wdata[127]~input_o ),
	.local_wdata_63(\local_wdata[63]~input_o ),
	.local_wdata_95(\local_wdata[95]~input_o ),
	.local_wdata_31(\local_wdata[31]~input_o ));

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[0]  = mem_dq[0];

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[1]  = mem_dq[1];

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[2]  = mem_dq[2];

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[3]  = mem_dq[3];

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[4]  = mem_dq[4];

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[5]  = mem_dq[5];

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[6]  = mem_dq[6];

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[7]  = mem_dq[7];

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[8]  = mem_dq[8];

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[9]  = mem_dq[9];

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[10]  = mem_dq[10];

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[11]  = mem_dq[11];

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[12]  = mem_dq[12];

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[13]  = mem_dq[13];

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[14]  = mem_dq[14];

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[15]  = mem_dq[15];

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[16]  = mem_dq[16];

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[17]  = mem_dq[17];

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[18]  = mem_dq[18];

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[19]  = mem_dq[19];

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[20]  = mem_dq[20];

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[21]  = mem_dq[21];

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[22]  = mem_dq[22];

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[23]  = mem_dq[23];

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[24]  = mem_dq[24];

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[25]  = mem_dq[25];

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[26]  = mem_dq[26];

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[27]  = mem_dq[27];

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[28]  = mem_dq[28];

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[29]  = mem_dq[29];

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[30]  = mem_dq[30];

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dq_datain[31]  = mem_dq[31];

arriaii_io_ibuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].ddr2_with_dqsn_buf_gen.dqs_inpt_ibuf (
	.i(mem_dqs[0]),
	.ibar(mem_dqsn[0]),
	.o(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_buffered[0] ));
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].ddr2_with_dqsn_buf_gen.dqs_inpt_ibuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].ddr2_with_dqsn_buf_gen.dqs_inpt_ibuf .differential_mode = "true";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].ddr2_with_dqsn_buf_gen.dqs_inpt_ibuf .simulate_z_as = "z";

arriaii_io_ibuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].ddr2_with_dqsn_buf_gen.dqs_inpt_ibuf (
	.i(mem_dqs[1]),
	.ibar(mem_dqsn[1]),
	.o(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_buffered[1] ));
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].ddr2_with_dqsn_buf_gen.dqs_inpt_ibuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].ddr2_with_dqsn_buf_gen.dqs_inpt_ibuf .differential_mode = "true";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].ddr2_with_dqsn_buf_gen.dqs_inpt_ibuf .simulate_z_as = "z";

arriaii_io_ibuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].ddr2_with_dqsn_buf_gen.dqs_inpt_ibuf (
	.i(mem_dqs[2]),
	.ibar(mem_dqsn[2]),
	.o(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_buffered[2] ));
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].ddr2_with_dqsn_buf_gen.dqs_inpt_ibuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].ddr2_with_dqsn_buf_gen.dqs_inpt_ibuf .differential_mode = "true";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].ddr2_with_dqsn_buf_gen.dqs_inpt_ibuf .simulate_z_as = "z";

arriaii_io_ibuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].ddr2_with_dqsn_buf_gen.dqs_inpt_ibuf (
	.i(mem_dqs[3]),
	.ibar(mem_dqsn[3]),
	.o(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_buffered[3] ));
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].ddr2_with_dqsn_buf_gen.dqs_inpt_ibuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].ddr2_with_dqsn_buf_gen.dqs_inpt_ibuf .differential_mode = "true";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].ddr2_with_dqsn_buf_gen.dqs_inpt_ibuf .simulate_z_as = "z";

assign \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|fb_clk  = mem_clk[0];

arriaii_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\~GND~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \~GND .extended_lut = "off";
defparam \~GND .lut_mask = 64'h0000000000000000;
defparam \~GND .shared_arith = "off";

assign \local_size[1]~input_o  = local_size[1];

assign \local_address[0]~input_o  = local_address[0];

assign \local_size[0]~input_o  = local_size[0];

assign \local_size[6]~input_o  = local_size[6];

assign \local_size[5]~input_o  = local_size[5];

assign \local_size[4]~input_o  = local_size[4];

assign \local_size[2]~input_o  = local_size[2];

assign \local_size[3]~input_o  = local_size[3];

assign \local_read_req~input_o  = local_read_req;

assign \local_write_req~input_o  = local_write_req;

assign \local_burstbegin~input_o  = local_burstbegin;

assign \global_reset_n~input_o  = global_reset_n;

assign \pll_ref_clk~input_o  = pll_ref_clk;

assign \soft_reset_n~input_o  = soft_reset_n;

assign \local_address[8]~input_o  = local_address[8];

assign \local_address[10]~input_o  = local_address[10];

assign \local_address[9]~input_o  = local_address[9];

assign \local_address[23]~input_o  = local_address[23];

assign \local_address[24]~input_o  = local_address[24];

assign \local_address[22]~input_o  = local_address[22];

assign \local_address[20]~input_o  = local_address[20];

assign \local_address[21]~input_o  = local_address[21];

assign \local_address[19]~input_o  = local_address[19];

assign \local_address[17]~input_o  = local_address[17];

assign \local_address[18]~input_o  = local_address[18];

assign \local_address[13]~input_o  = local_address[13];

assign \local_address[11]~input_o  = local_address[11];

assign \local_address[12]~input_o  = local_address[12];

assign \local_address[16]~input_o  = local_address[16];

assign \local_address[14]~input_o  = local_address[14];

assign \local_address[15]~input_o  = local_address[15];

assign \local_address[1]~input_o  = local_address[1];

assign \local_address[2]~input_o  = local_address[2];

assign \local_address[3]~input_o  = local_address[3];

assign \local_address[4]~input_o  = local_address[4];

assign \local_address[5]~input_o  = local_address[5];

assign \local_address[7]~input_o  = local_address[7];

assign \local_address[6]~input_o  = local_address[6];

assign \local_be[4]~input_o  = local_be[4];

assign \local_be[12]~input_o  = local_be[12];

assign \local_be[0]~input_o  = local_be[0];

assign \local_be[8]~input_o  = local_be[8];

assign \local_be[5]~input_o  = local_be[5];

assign \local_be[13]~input_o  = local_be[13];

assign \local_be[1]~input_o  = local_be[1];

assign \local_be[9]~input_o  = local_be[9];

assign \local_be[6]~input_o  = local_be[6];

assign \local_be[14]~input_o  = local_be[14];

assign \local_be[2]~input_o  = local_be[2];

assign \local_be[10]~input_o  = local_be[10];

assign \local_be[7]~input_o  = local_be[7];

assign \local_be[15]~input_o  = local_be[15];

assign \local_be[3]~input_o  = local_be[3];

assign \local_be[11]~input_o  = local_be[11];

assign \local_wdata[96]~input_o  = local_wdata[96];

assign \local_wdata[32]~input_o  = local_wdata[32];

assign \local_wdata[64]~input_o  = local_wdata[64];

assign \local_wdata[0]~input_o  = local_wdata[0];

assign \local_wdata[97]~input_o  = local_wdata[97];

assign \local_wdata[33]~input_o  = local_wdata[33];

assign \local_wdata[65]~input_o  = local_wdata[65];

assign \local_wdata[1]~input_o  = local_wdata[1];

assign \local_wdata[98]~input_o  = local_wdata[98];

assign \local_wdata[34]~input_o  = local_wdata[34];

assign \local_wdata[66]~input_o  = local_wdata[66];

assign \local_wdata[2]~input_o  = local_wdata[2];

assign \local_wdata[99]~input_o  = local_wdata[99];

assign \local_wdata[35]~input_o  = local_wdata[35];

assign \local_wdata[67]~input_o  = local_wdata[67];

assign \local_wdata[3]~input_o  = local_wdata[3];

assign \local_wdata[100]~input_o  = local_wdata[100];

assign \local_wdata[36]~input_o  = local_wdata[36];

assign \local_wdata[68]~input_o  = local_wdata[68];

assign \local_wdata[4]~input_o  = local_wdata[4];

assign \local_wdata[101]~input_o  = local_wdata[101];

assign \local_wdata[37]~input_o  = local_wdata[37];

assign \local_wdata[69]~input_o  = local_wdata[69];

assign \local_wdata[5]~input_o  = local_wdata[5];

assign \local_wdata[102]~input_o  = local_wdata[102];

assign \local_wdata[38]~input_o  = local_wdata[38];

assign \local_wdata[70]~input_o  = local_wdata[70];

assign \local_wdata[6]~input_o  = local_wdata[6];

assign \local_wdata[103]~input_o  = local_wdata[103];

assign \local_wdata[39]~input_o  = local_wdata[39];

assign \local_wdata[71]~input_o  = local_wdata[71];

assign \local_wdata[7]~input_o  = local_wdata[7];

assign \local_wdata[104]~input_o  = local_wdata[104];

assign \local_wdata[40]~input_o  = local_wdata[40];

assign \local_wdata[72]~input_o  = local_wdata[72];

assign \local_wdata[8]~input_o  = local_wdata[8];

assign \local_wdata[105]~input_o  = local_wdata[105];

assign \local_wdata[41]~input_o  = local_wdata[41];

assign \local_wdata[73]~input_o  = local_wdata[73];

assign \local_wdata[9]~input_o  = local_wdata[9];

assign \local_wdata[106]~input_o  = local_wdata[106];

assign \local_wdata[42]~input_o  = local_wdata[42];

assign \local_wdata[74]~input_o  = local_wdata[74];

assign \local_wdata[10]~input_o  = local_wdata[10];

assign \local_wdata[107]~input_o  = local_wdata[107];

assign \local_wdata[43]~input_o  = local_wdata[43];

assign \local_wdata[75]~input_o  = local_wdata[75];

assign \local_wdata[11]~input_o  = local_wdata[11];

assign \local_wdata[108]~input_o  = local_wdata[108];

assign \local_wdata[44]~input_o  = local_wdata[44];

assign \local_wdata[76]~input_o  = local_wdata[76];

assign \local_wdata[12]~input_o  = local_wdata[12];

assign \local_wdata[109]~input_o  = local_wdata[109];

assign \local_wdata[45]~input_o  = local_wdata[45];

assign \local_wdata[77]~input_o  = local_wdata[77];

assign \local_wdata[13]~input_o  = local_wdata[13];

assign \local_wdata[110]~input_o  = local_wdata[110];

assign \local_wdata[46]~input_o  = local_wdata[46];

assign \local_wdata[78]~input_o  = local_wdata[78];

assign \local_wdata[14]~input_o  = local_wdata[14];

assign \local_wdata[111]~input_o  = local_wdata[111];

assign \local_wdata[47]~input_o  = local_wdata[47];

assign \local_wdata[79]~input_o  = local_wdata[79];

assign \local_wdata[15]~input_o  = local_wdata[15];

assign \local_wdata[112]~input_o  = local_wdata[112];

assign \local_wdata[48]~input_o  = local_wdata[48];

assign \local_wdata[80]~input_o  = local_wdata[80];

assign \local_wdata[16]~input_o  = local_wdata[16];

assign \local_wdata[113]~input_o  = local_wdata[113];

assign \local_wdata[49]~input_o  = local_wdata[49];

assign \local_wdata[81]~input_o  = local_wdata[81];

assign \local_wdata[17]~input_o  = local_wdata[17];

assign \local_wdata[114]~input_o  = local_wdata[114];

assign \local_wdata[50]~input_o  = local_wdata[50];

assign \local_wdata[82]~input_o  = local_wdata[82];

assign \local_wdata[18]~input_o  = local_wdata[18];

assign \local_wdata[115]~input_o  = local_wdata[115];

assign \local_wdata[51]~input_o  = local_wdata[51];

assign \local_wdata[83]~input_o  = local_wdata[83];

assign \local_wdata[19]~input_o  = local_wdata[19];

assign \local_wdata[116]~input_o  = local_wdata[116];

assign \local_wdata[52]~input_o  = local_wdata[52];

assign \local_wdata[84]~input_o  = local_wdata[84];

assign \local_wdata[20]~input_o  = local_wdata[20];

assign \local_wdata[117]~input_o  = local_wdata[117];

assign \local_wdata[53]~input_o  = local_wdata[53];

assign \local_wdata[85]~input_o  = local_wdata[85];

assign \local_wdata[21]~input_o  = local_wdata[21];

assign \local_wdata[118]~input_o  = local_wdata[118];

assign \local_wdata[54]~input_o  = local_wdata[54];

assign \local_wdata[86]~input_o  = local_wdata[86];

assign \local_wdata[22]~input_o  = local_wdata[22];

assign \local_wdata[119]~input_o  = local_wdata[119];

assign \local_wdata[55]~input_o  = local_wdata[55];

assign \local_wdata[87]~input_o  = local_wdata[87];

assign \local_wdata[23]~input_o  = local_wdata[23];

assign \local_wdata[120]~input_o  = local_wdata[120];

assign \local_wdata[56]~input_o  = local_wdata[56];

assign \local_wdata[88]~input_o  = local_wdata[88];

assign \local_wdata[24]~input_o  = local_wdata[24];

assign \local_wdata[121]~input_o  = local_wdata[121];

assign \local_wdata[57]~input_o  = local_wdata[57];

assign \local_wdata[89]~input_o  = local_wdata[89];

assign \local_wdata[25]~input_o  = local_wdata[25];

assign \local_wdata[122]~input_o  = local_wdata[122];

assign \local_wdata[58]~input_o  = local_wdata[58];

assign \local_wdata[90]~input_o  = local_wdata[90];

assign \local_wdata[26]~input_o  = local_wdata[26];

assign \local_wdata[123]~input_o  = local_wdata[123];

assign \local_wdata[59]~input_o  = local_wdata[59];

assign \local_wdata[91]~input_o  = local_wdata[91];

assign \local_wdata[27]~input_o  = local_wdata[27];

assign \local_wdata[124]~input_o  = local_wdata[124];

assign \local_wdata[60]~input_o  = local_wdata[60];

assign \local_wdata[92]~input_o  = local_wdata[92];

assign \local_wdata[28]~input_o  = local_wdata[28];

assign \local_wdata[125]~input_o  = local_wdata[125];

assign \local_wdata[61]~input_o  = local_wdata[61];

assign \local_wdata[93]~input_o  = local_wdata[93];

assign \local_wdata[29]~input_o  = local_wdata[29];

assign \local_wdata[126]~input_o  = local_wdata[126];

assign \local_wdata[62]~input_o  = local_wdata[62];

assign \local_wdata[94]~input_o  = local_wdata[94];

assign \local_wdata[30]~input_o  = local_wdata[30];

assign \local_wdata[127]~input_o  = local_wdata[127];

assign \local_wdata[63]~input_o  = local_wdata[63];

assign \local_wdata[95]~input_o  = local_wdata[95];

assign \local_wdata[31]~input_o  = local_wdata[31];

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].gen_dm.dm_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|wire_output_dq_0_output_ddio_out_inst_dataout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dm[0]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].gen_dm.dm_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].gen_dm.dm_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].gen_dm.dm_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|wire_output_dq_0_output_ddio_out_inst_dataout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dm[1]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].gen_dm.dm_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].gen_dm.dm_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].gen_dm.dm_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|wire_output_dq_0_output_ddio_out_inst_dataout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dm[2]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].gen_dm.dm_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].gen_dm.dm_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].gen_dm.dm_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|wire_output_dq_0_output_ddio_out_inst_dataout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dm[3]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].gen_dm.dm_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].gen_dm.dm_obuf .open_drain_output = "false";

assign local_ready = \ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|cmd_gen_inst|ready_out~combout ;

assign local_rdata[0] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[0] ;

assign local_rdata[1] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[1] ;

assign local_rdata[2] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[2] ;

assign local_rdata[3] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[3] ;

assign local_rdata[4] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[4] ;

assign local_rdata[5] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[5] ;

assign local_rdata[6] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[6] ;

assign local_rdata[7] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[7] ;

assign local_rdata[8] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[16] ;

assign local_rdata[9] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[17] ;

assign local_rdata[10] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[18] ;

assign local_rdata[11] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[19] ;

assign local_rdata[12] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[20] ;

assign local_rdata[13] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[21] ;

assign local_rdata[14] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[22] ;

assign local_rdata[15] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[23] ;

assign local_rdata[16] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[32] ;

assign local_rdata[17] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[33] ;

assign local_rdata[18] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[34] ;

assign local_rdata[19] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[35] ;

assign local_rdata[20] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[36] ;

assign local_rdata[21] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[37] ;

assign local_rdata[22] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[38] ;

assign local_rdata[23] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[39] ;

assign local_rdata[24] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[48] ;

assign local_rdata[25] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[49] ;

assign local_rdata[26] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[50] ;

assign local_rdata[27] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[51] ;

assign local_rdata[28] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[52] ;

assign local_rdata[29] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[53] ;

assign local_rdata[30] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[54] ;

assign local_rdata[31] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[55] ;

assign local_rdata[32] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[8] ;

assign local_rdata[33] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[9] ;

assign local_rdata[34] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[10] ;

assign local_rdata[35] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[11] ;

assign local_rdata[36] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[12] ;

assign local_rdata[37] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[13] ;

assign local_rdata[38] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[14] ;

assign local_rdata[39] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[15] ;

assign local_rdata[40] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[24] ;

assign local_rdata[41] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[25] ;

assign local_rdata[42] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[26] ;

assign local_rdata[43] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[27] ;

assign local_rdata[44] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[28] ;

assign local_rdata[45] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[29] ;

assign local_rdata[46] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[30] ;

assign local_rdata[47] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[31] ;

assign local_rdata[48] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[40] ;

assign local_rdata[49] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[41] ;

assign local_rdata[50] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[42] ;

assign local_rdata[51] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[43] ;

assign local_rdata[52] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[44] ;

assign local_rdata[53] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[45] ;

assign local_rdata[54] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[46] ;

assign local_rdata[55] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[47] ;

assign local_rdata[56] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[56] ;

assign local_rdata[57] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[57] ;

assign local_rdata[58] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[58] ;

assign local_rdata[59] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[59] ;

assign local_rdata[60] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[60] ;

assign local_rdata[61] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[61] ;

assign local_rdata[62] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[62] ;

assign local_rdata[63] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[63] ;

assign local_rdata[64] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[64] ;

assign local_rdata[65] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[65] ;

assign local_rdata[66] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[66] ;

assign local_rdata[67] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[67] ;

assign local_rdata[68] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[68] ;

assign local_rdata[69] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[69] ;

assign local_rdata[70] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[70] ;

assign local_rdata[71] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[71] ;

assign local_rdata[72] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[80] ;

assign local_rdata[73] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[81] ;

assign local_rdata[74] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[82] ;

assign local_rdata[75] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[83] ;

assign local_rdata[76] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[84] ;

assign local_rdata[77] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[85] ;

assign local_rdata[78] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[86] ;

assign local_rdata[79] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[87] ;

assign local_rdata[80] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[96] ;

assign local_rdata[81] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[97] ;

assign local_rdata[82] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[98] ;

assign local_rdata[83] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[99] ;

assign local_rdata[84] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[100] ;

assign local_rdata[85] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[101] ;

assign local_rdata[86] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[102] ;

assign local_rdata[87] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[103] ;

assign local_rdata[88] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[112] ;

assign local_rdata[89] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[113] ;

assign local_rdata[90] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[114] ;

assign local_rdata[91] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[115] ;

assign local_rdata[92] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[116] ;

assign local_rdata[93] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[117] ;

assign local_rdata[94] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[118] ;

assign local_rdata[95] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[119] ;

assign local_rdata[96] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[72] ;

assign local_rdata[97] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[73] ;

assign local_rdata[98] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[74] ;

assign local_rdata[99] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[75] ;

assign local_rdata[100] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[76] ;

assign local_rdata[101] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[77] ;

assign local_rdata[102] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[78] ;

assign local_rdata[103] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[79] ;

assign local_rdata[104] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[88] ;

assign local_rdata[105] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[89] ;

assign local_rdata[106] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[90] ;

assign local_rdata[107] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[91] ;

assign local_rdata[108] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[92] ;

assign local_rdata[109] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[93] ;

assign local_rdata[110] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[94] ;

assign local_rdata[111] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[95] ;

assign local_rdata[112] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[104] ;

assign local_rdata[113] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[105] ;

assign local_rdata[114] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[106] ;

assign local_rdata[115] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[107] ;

assign local_rdata[116] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[108] ;

assign local_rdata[117] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[109] ;

assign local_rdata[118] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[110] ;

assign local_rdata[119] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[111] ;

assign local_rdata[120] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[120] ;

assign local_rdata[121] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[121] ;

assign local_rdata[122] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[122] ;

assign local_rdata[123] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[123] ;

assign local_rdata[124] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[124] ;

assign local_rdata[125] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[125] ;

assign local_rdata[126] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[126] ;

assign local_rdata[127] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdp|half_rate_ram_gen.altsyncram_component|auto_generated|q_b[127] ;

assign local_rdata_valid = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|rdv_pipe|ctl_rdata_valid[0]~q ;

assign reset_request_n = ~ \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|half_rate.pll|altpll_component|auto_generated|locked~combout ;

assign mem_odt[0] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|gen_odt.odt[0].odt_struct|half_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_cs_n[0] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|cs_n[0].cs_n_struct|half_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_cke[0] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|cke[0].cke_struct|half_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_addr[0] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[0].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_addr[1] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[1].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_addr[2] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[2].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_addr[3] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[3].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_addr[4] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[4].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_addr[5] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[5].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_addr[6] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[6].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_addr[7] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[7].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_addr[8] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[8].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_addr[9] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[9].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_addr[10] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[10].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_addr[11] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[11].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_addr[12] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[12].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_addr[13] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|addr[13].addr_struct|half_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_ba[0] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|ba[0].ba_struct|half_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_ba[1] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|ba[1].ba_struct|half_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_ba[2] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|ba[2].ba_struct|half_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_ras_n = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|ras_n_struct|half_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_cas_n = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|cas_n_struct|half_rate.addr_pin|auto_generated|dataout[0] ;

assign mem_we_n = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|we_n_struct|half_rate.addr_pin|auto_generated|dataout[0] ;

assign local_refresh_ack = \ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|state_machine_inst|int_refresh_ack~q ;

assign local_wdata_req = gnd;

assign local_init_done = \ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|local_init_done~combout ;

assign reset_phy_clk_n = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|reset_phy_clk_1x_n~q ;

assign mem_reset_n = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|half_rate_adc_gen.adc|ddr3_rst.ddr3_rst_struct|half_rate.addr_pin|auto_generated|dataout[0] ;

assign dll_reference_clk = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|half_rate.pll|altpll_component|auto_generated|clk[1] ;

assign dqs_delay_ctrl_export[0] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|dqs_delay_ctrl[0] ;

assign dqs_delay_ctrl_export[1] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|dqs_delay_ctrl[1] ;

assign dqs_delay_ctrl_export[2] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|dqs_delay_ctrl[2] ;

assign dqs_delay_ctrl_export[3] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|dqs_delay_ctrl[3] ;

assign dqs_delay_ctrl_export[4] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|dqs_delay_ctrl[4] ;

assign dqs_delay_ctrl_export[5] = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|dqs_delay_ctrl[5] ;

assign phy_clk = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|half_rate.pll|altpll_component|auto_generated|clk[0] ;

assign aux_full_rate_clk = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|half_rate.pll|altpll_component|auto_generated|clk[1] ;

assign aux_half_rate_clk = \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|half_rate.pll|altpll_component|auto_generated|clk[0] ;

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|DDR_CLK_OUT[0].mem_clk_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|mem_clk_buf_in[0] ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_clk[0]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|DDR_CLK_OUT[0].mem_clk_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|DDR_CLK_OUT[0].mem_clk_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|DDR_CLK_OUT[0].mem_clk_n_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|mem_clk_n_buf_in[0] ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_clk_n[0]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|DDR_CLK_OUT[0].mem_clk_n_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|clk|DDR_CLK_OUT[0].mem_clk_n_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[0].dq_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|wire_bidir_dq_0_output_ddio_out_inst_dataout ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|bidir_dq_0_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[0]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[0].dq_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[0].dq_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[1].dq_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|wire_bidir_dq_1_output_ddio_out_inst_dataout ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|bidir_dq_1_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[1]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[1].dq_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[1].dq_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[2].dq_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|wire_bidir_dq_2_output_ddio_out_inst_dataout ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|bidir_dq_2_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[2]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[2].dq_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[2].dq_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[3].dq_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|wire_bidir_dq_3_output_ddio_out_inst_dataout ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|bidir_dq_3_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[3]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[3].dq_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[3].dq_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[4].dq_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|wire_bidir_dq_4_output_ddio_out_inst_dataout ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|bidir_dq_4_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[4]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[4].dq_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[4].dq_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[5].dq_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|wire_bidir_dq_5_output_ddio_out_inst_dataout ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|bidir_dq_5_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[5]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[5].dq_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[5].dq_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[6].dq_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|wire_bidir_dq_6_output_ddio_out_inst_dataout ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|bidir_dq_6_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[6]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[6].dq_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[6].dq_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[7].dq_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|wire_bidir_dq_7_output_ddio_out_inst_dataout ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|bidir_dq_7_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[7]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[7].dq_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq[7].dq_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[0].dq_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|wire_bidir_dq_0_output_ddio_out_inst_dataout ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|bidir_dq_0_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[8]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[0].dq_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[0].dq_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[1].dq_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|wire_bidir_dq_1_output_ddio_out_inst_dataout ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|bidir_dq_1_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[9]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[1].dq_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[1].dq_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[2].dq_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|wire_bidir_dq_2_output_ddio_out_inst_dataout ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|bidir_dq_2_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[10]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[2].dq_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[2].dq_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[3].dq_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|wire_bidir_dq_3_output_ddio_out_inst_dataout ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|bidir_dq_3_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[11]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[3].dq_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[3].dq_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[4].dq_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|wire_bidir_dq_4_output_ddio_out_inst_dataout ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|bidir_dq_4_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[12]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[4].dq_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[4].dq_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[5].dq_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|wire_bidir_dq_5_output_ddio_out_inst_dataout ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|bidir_dq_5_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[13]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[5].dq_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[5].dq_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[6].dq_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|wire_bidir_dq_6_output_ddio_out_inst_dataout ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|bidir_dq_6_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[14]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[6].dq_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[6].dq_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[7].dq_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|wire_bidir_dq_7_output_ddio_out_inst_dataout ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|bidir_dq_7_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[15]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[7].dq_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq[7].dq_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq[0].dq_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|wire_bidir_dq_0_output_ddio_out_inst_dataout ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|bidir_dq_0_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[16]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq[0].dq_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq[0].dq_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq[1].dq_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|wire_bidir_dq_1_output_ddio_out_inst_dataout ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|bidir_dq_1_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[17]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq[1].dq_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq[1].dq_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq[2].dq_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|wire_bidir_dq_2_output_ddio_out_inst_dataout ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|bidir_dq_2_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[18]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq[2].dq_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq[2].dq_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq[3].dq_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|wire_bidir_dq_3_output_ddio_out_inst_dataout ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|bidir_dq_3_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[19]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq[3].dq_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq[3].dq_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq[4].dq_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|wire_bidir_dq_4_output_ddio_out_inst_dataout ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|bidir_dq_4_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[20]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq[4].dq_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq[4].dq_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq[5].dq_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|wire_bidir_dq_5_output_ddio_out_inst_dataout ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|bidir_dq_5_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[21]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq[5].dq_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq[5].dq_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq[6].dq_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|wire_bidir_dq_6_output_ddio_out_inst_dataout ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|bidir_dq_6_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[22]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq[6].dq_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq[6].dq_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq[7].dq_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|wire_bidir_dq_7_output_ddio_out_inst_dataout ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|bidir_dq_7_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[23]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq[7].dq_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq[7].dq_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq[0].dq_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|wire_bidir_dq_0_output_ddio_out_inst_dataout ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|bidir_dq_0_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[24]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq[0].dq_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq[0].dq_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq[1].dq_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|wire_bidir_dq_1_output_ddio_out_inst_dataout ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|bidir_dq_1_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[25]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq[1].dq_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq[1].dq_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq[2].dq_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|wire_bidir_dq_2_output_ddio_out_inst_dataout ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|bidir_dq_2_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[26]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq[2].dq_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq[2].dq_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq[3].dq_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|wire_bidir_dq_3_output_ddio_out_inst_dataout ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|bidir_dq_3_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[27]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq[3].dq_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq[3].dq_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq[4].dq_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|wire_bidir_dq_4_output_ddio_out_inst_dataout ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|bidir_dq_4_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[28]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq[4].dq_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq[4].dq_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq[5].dq_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|wire_bidir_dq_5_output_ddio_out_inst_dataout ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|bidir_dq_5_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[29]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq[5].dq_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq[5].dq_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq[6].dq_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|wire_bidir_dq_6_output_ddio_out_inst_dataout ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|bidir_dq_6_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[30]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq[6].dq_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq[6].dq_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq[7].dq_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|wire_bidir_dq_7_output_ddio_out_inst_dataout ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|bidir_dq_7_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dq[31]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq[7].dq_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq[7].dq_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].ddr2_with_dqsn_buf_gen.dqs_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_pseudo_diff_out[0] ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|dqs_0_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dqs[0]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].ddr2_with_dqsn_buf_gen.dqs_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].ddr2_with_dqsn_buf_gen.dqs_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].ddr2_with_dqsn_buf_gen.dqs_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_pseudo_diff_out[1] ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|dqs_0_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dqs[1]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].ddr2_with_dqsn_buf_gen.dqs_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].ddr2_with_dqsn_buf_gen.dqs_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].ddr2_with_dqsn_buf_gen.dqs_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_pseudo_diff_out[2] ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|dqs_0_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dqs[2]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].ddr2_with_dqsn_buf_gen.dqs_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].ddr2_with_dqsn_buf_gen.dqs_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].ddr2_with_dqsn_buf_gen.dqs_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_pseudo_diff_out[3] ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|dqs_0_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dqs[3]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].ddr2_with_dqsn_buf_gen.dqs_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].ddr2_with_dqsn_buf_gen.dqs_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].ddr2_with_dqsn_buf_gen.dqsn_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqsn_pseudo_diff_out[0] ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].dq_dqs|dqsn_0_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dqsn[0]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].ddr2_with_dqsn_buf_gen.dqsn_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[0].ddr2_with_dqsn_buf_gen.dqsn_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].ddr2_with_dqsn_buf_gen.dqsn_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqsn_pseudo_diff_out[1] ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].dq_dqs|dqsn_0_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dqsn[1]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].ddr2_with_dqsn_buf_gen.dqsn_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[1].ddr2_with_dqsn_buf_gen.dqsn_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].ddr2_with_dqsn_buf_gen.dqsn_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqsn_pseudo_diff_out[2] ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].dq_dqs|dqsn_0_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dqsn[2]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].ddr2_with_dqsn_buf_gen.dqsn_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[2].ddr2_with_dqsn_buf_gen.dqsn_obuf .open_drain_output = "false";

arriaii_io_obuf \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].ddr2_with_dqsn_buf_gen.dqsn_obuf (
	.i(\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqsn_pseudo_diff_out[3] ),
	.oe(!\ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].dq_dqs|dqsn_0_oe_ff_inst~q ),
	.seriesterminationcontrol(16'b0000000000000000),
	.o(mem_dqsn[3]),
	.obar());
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].ddr2_with_dqsn_buf_gen.dqsn_obuf .bus_hold = "false";
defparam \ddr3_int_controller_phy_inst|ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|dpio|dqs_group[3].ddr2_with_dqsn_buf_gen.dqsn_obuf .open_drain_output = "false";

assign \mem_clk_n[0]~input_o  = mem_clk_n[0];

endmodule

module ddr3_int_ddr3_int_controller_phy (
	q_b_0,
	q_b_64,
	q_b_1,
	q_b_65,
	q_b_2,
	q_b_66,
	q_b_3,
	q_b_67,
	q_b_4,
	q_b_68,
	q_b_5,
	q_b_69,
	q_b_6,
	q_b_70,
	q_b_7,
	q_b_71,
	q_b_16,
	q_b_80,
	q_b_17,
	q_b_81,
	q_b_18,
	q_b_82,
	q_b_19,
	q_b_83,
	q_b_20,
	q_b_84,
	q_b_21,
	q_b_85,
	q_b_22,
	q_b_86,
	q_b_23,
	q_b_87,
	q_b_32,
	q_b_96,
	q_b_33,
	q_b_97,
	q_b_34,
	q_b_98,
	q_b_35,
	q_b_99,
	q_b_36,
	q_b_100,
	q_b_37,
	q_b_101,
	q_b_38,
	q_b_102,
	q_b_39,
	q_b_103,
	q_b_48,
	q_b_112,
	q_b_49,
	q_b_113,
	q_b_50,
	q_b_114,
	q_b_51,
	q_b_115,
	q_b_52,
	q_b_116,
	q_b_53,
	q_b_117,
	q_b_54,
	q_b_118,
	q_b_55,
	q_b_119,
	q_b_8,
	q_b_72,
	q_b_9,
	q_b_73,
	q_b_10,
	q_b_74,
	q_b_11,
	q_b_75,
	q_b_12,
	q_b_76,
	q_b_13,
	q_b_77,
	q_b_14,
	q_b_78,
	q_b_15,
	q_b_79,
	q_b_24,
	q_b_88,
	q_b_25,
	q_b_89,
	q_b_26,
	q_b_90,
	q_b_27,
	q_b_91,
	q_b_28,
	q_b_92,
	q_b_29,
	q_b_93,
	q_b_30,
	q_b_94,
	q_b_31,
	q_b_95,
	q_b_40,
	q_b_104,
	q_b_41,
	q_b_105,
	q_b_42,
	q_b_106,
	q_b_43,
	q_b_107,
	q_b_44,
	q_b_108,
	q_b_45,
	q_b_109,
	q_b_46,
	q_b_110,
	q_b_47,
	q_b_111,
	q_b_56,
	q_b_120,
	q_b_57,
	q_b_121,
	q_b_58,
	q_b_122,
	q_b_59,
	q_b_123,
	q_b_60,
	q_b_124,
	q_b_61,
	q_b_125,
	q_b_62,
	q_b_126,
	q_b_63,
	q_b_127,
	clk_0,
	clk_1,
	dataout_0,
	dataout_01,
	dataout_02,
	dataout_03,
	dataout_04,
	dataout_05,
	dataout_06,
	dataout_07,
	dataout_08,
	dataout_09,
	dataout_010,
	dataout_011,
	dataout_012,
	dataout_013,
	dataout_014,
	dataout_015,
	dataout_016,
	dataout_017,
	dataout_018,
	dataout_019,
	dataout_020,
	dataout_021,
	dataout_022,
	dataout_023,
	dqs_delay_ctrl_0,
	dqs_delay_ctrl_1,
	dqs_delay_ctrl_2,
	dqs_delay_ctrl_3,
	dqs_delay_ctrl_4,
	dqs_delay_ctrl_5,
	wire_output_dq_0_output_ddio_out_inst_dataout,
	wire_output_dq_0_output_ddio_out_inst_dataout1,
	wire_output_dq_0_output_ddio_out_inst_dataout2,
	wire_output_dq_0_output_ddio_out_inst_dataout3,
	mem_clk_buf_in_0,
	mem_clk_n_buf_in_0,
	wire_bidir_dq_0_output_ddio_out_inst_dataout,
	wire_bidir_dq_1_output_ddio_out_inst_dataout,
	wire_bidir_dq_2_output_ddio_out_inst_dataout,
	wire_bidir_dq_3_output_ddio_out_inst_dataout,
	wire_bidir_dq_4_output_ddio_out_inst_dataout,
	wire_bidir_dq_5_output_ddio_out_inst_dataout,
	wire_bidir_dq_6_output_ddio_out_inst_dataout,
	wire_bidir_dq_7_output_ddio_out_inst_dataout,
	wire_bidir_dq_0_output_ddio_out_inst_dataout1,
	wire_bidir_dq_1_output_ddio_out_inst_dataout1,
	wire_bidir_dq_2_output_ddio_out_inst_dataout1,
	wire_bidir_dq_3_output_ddio_out_inst_dataout1,
	wire_bidir_dq_4_output_ddio_out_inst_dataout1,
	wire_bidir_dq_5_output_ddio_out_inst_dataout1,
	wire_bidir_dq_6_output_ddio_out_inst_dataout1,
	wire_bidir_dq_7_output_ddio_out_inst_dataout1,
	wire_bidir_dq_0_output_ddio_out_inst_dataout2,
	wire_bidir_dq_1_output_ddio_out_inst_dataout2,
	wire_bidir_dq_2_output_ddio_out_inst_dataout2,
	wire_bidir_dq_3_output_ddio_out_inst_dataout2,
	wire_bidir_dq_4_output_ddio_out_inst_dataout2,
	wire_bidir_dq_5_output_ddio_out_inst_dataout2,
	wire_bidir_dq_6_output_ddio_out_inst_dataout2,
	wire_bidir_dq_7_output_ddio_out_inst_dataout2,
	wire_bidir_dq_0_output_ddio_out_inst_dataout3,
	wire_bidir_dq_1_output_ddio_out_inst_dataout3,
	wire_bidir_dq_2_output_ddio_out_inst_dataout3,
	wire_bidir_dq_3_output_ddio_out_inst_dataout3,
	wire_bidir_dq_4_output_ddio_out_inst_dataout3,
	wire_bidir_dq_5_output_ddio_out_inst_dataout3,
	wire_bidir_dq_6_output_ddio_out_inst_dataout3,
	wire_bidir_dq_7_output_ddio_out_inst_dataout3,
	dqs_pseudo_diff_out_0,
	dqsn_pseudo_diff_out_0,
	dqs_pseudo_diff_out_1,
	dqsn_pseudo_diff_out_1,
	dqs_pseudo_diff_out_2,
	dqsn_pseudo_diff_out_2,
	dqs_pseudo_diff_out_3,
	dqsn_pseudo_diff_out_3,
	dq_datain_0,
	dq_datain_1,
	dq_datain_2,
	dq_datain_3,
	dq_datain_4,
	dq_datain_5,
	dq_datain_6,
	dq_datain_7,
	dq_datain_8,
	dq_datain_9,
	dq_datain_10,
	dq_datain_11,
	dq_datain_12,
	dq_datain_13,
	dq_datain_14,
	dq_datain_15,
	dq_datain_16,
	dq_datain_17,
	dq_datain_18,
	dq_datain_19,
	dq_datain_20,
	dq_datain_21,
	dq_datain_22,
	dq_datain_23,
	dq_datain_24,
	dq_datain_25,
	dq_datain_26,
	dq_datain_27,
	dq_datain_28,
	dq_datain_29,
	dq_datain_30,
	dq_datain_31,
	dqs_buffered_0,
	dqs_buffered_1,
	dqs_buffered_2,
	dqs_buffered_3,
	fb_clk,
	ready_out,
	ctl_rdata_valid_0,
	reset_request_n,
	int_refresh_ack,
	local_init_done,
	reset_phy_clk_1x_n,
	bidir_dq_0_oe_ff_inst,
	bidir_dq_1_oe_ff_inst,
	bidir_dq_2_oe_ff_inst,
	bidir_dq_3_oe_ff_inst,
	bidir_dq_4_oe_ff_inst,
	bidir_dq_5_oe_ff_inst,
	bidir_dq_6_oe_ff_inst,
	bidir_dq_7_oe_ff_inst,
	bidir_dq_0_oe_ff_inst1,
	bidir_dq_1_oe_ff_inst1,
	bidir_dq_2_oe_ff_inst1,
	bidir_dq_3_oe_ff_inst1,
	bidir_dq_4_oe_ff_inst1,
	bidir_dq_5_oe_ff_inst1,
	bidir_dq_6_oe_ff_inst1,
	bidir_dq_7_oe_ff_inst1,
	bidir_dq_0_oe_ff_inst2,
	bidir_dq_1_oe_ff_inst2,
	bidir_dq_2_oe_ff_inst2,
	bidir_dq_3_oe_ff_inst2,
	bidir_dq_4_oe_ff_inst2,
	bidir_dq_5_oe_ff_inst2,
	bidir_dq_6_oe_ff_inst2,
	bidir_dq_7_oe_ff_inst2,
	bidir_dq_0_oe_ff_inst3,
	bidir_dq_1_oe_ff_inst3,
	bidir_dq_2_oe_ff_inst3,
	bidir_dq_3_oe_ff_inst3,
	bidir_dq_4_oe_ff_inst3,
	bidir_dq_5_oe_ff_inst3,
	bidir_dq_6_oe_ff_inst3,
	bidir_dq_7_oe_ff_inst3,
	dqs_0_oe_ff_inst,
	dqs_0_oe_ff_inst1,
	dqs_0_oe_ff_inst2,
	dqs_0_oe_ff_inst3,
	dqsn_0_oe_ff_inst,
	dqsn_0_oe_ff_inst1,
	dqsn_0_oe_ff_inst2,
	dqsn_0_oe_ff_inst3,
	GND_port,
	local_size_1,
	local_address_0,
	local_size_0,
	local_size_6,
	local_size_5,
	local_size_4,
	local_size_2,
	local_size_3,
	local_read_req,
	local_write_req,
	local_burstbegin,
	global_reset_n,
	pll_ref_clk,
	soft_reset_n,
	local_address_8,
	local_address_10,
	local_address_9,
	local_address_23,
	local_address_24,
	local_address_22,
	local_address_20,
	local_address_21,
	local_address_19,
	local_address_17,
	local_address_18,
	local_address_13,
	local_address_11,
	local_address_12,
	local_address_16,
	local_address_14,
	local_address_15,
	local_address_1,
	local_address_2,
	local_address_3,
	local_address_4,
	local_address_5,
	local_address_7,
	local_address_6,
	local_be_4,
	local_be_12,
	local_be_0,
	local_be_8,
	local_be_5,
	local_be_13,
	local_be_1,
	local_be_9,
	local_be_6,
	local_be_14,
	local_be_2,
	local_be_10,
	local_be_7,
	local_be_15,
	local_be_3,
	local_be_11,
	local_wdata_96,
	local_wdata_32,
	local_wdata_64,
	local_wdata_0,
	local_wdata_97,
	local_wdata_33,
	local_wdata_65,
	local_wdata_1,
	local_wdata_98,
	local_wdata_34,
	local_wdata_66,
	local_wdata_2,
	local_wdata_99,
	local_wdata_35,
	local_wdata_67,
	local_wdata_3,
	local_wdata_100,
	local_wdata_36,
	local_wdata_68,
	local_wdata_4,
	local_wdata_101,
	local_wdata_37,
	local_wdata_69,
	local_wdata_5,
	local_wdata_102,
	local_wdata_38,
	local_wdata_70,
	local_wdata_6,
	local_wdata_103,
	local_wdata_39,
	local_wdata_71,
	local_wdata_7,
	local_wdata_104,
	local_wdata_40,
	local_wdata_72,
	local_wdata_8,
	local_wdata_105,
	local_wdata_41,
	local_wdata_73,
	local_wdata_9,
	local_wdata_106,
	local_wdata_42,
	local_wdata_74,
	local_wdata_10,
	local_wdata_107,
	local_wdata_43,
	local_wdata_75,
	local_wdata_11,
	local_wdata_108,
	local_wdata_44,
	local_wdata_76,
	local_wdata_12,
	local_wdata_109,
	local_wdata_45,
	local_wdata_77,
	local_wdata_13,
	local_wdata_110,
	local_wdata_46,
	local_wdata_78,
	local_wdata_14,
	local_wdata_111,
	local_wdata_47,
	local_wdata_79,
	local_wdata_15,
	local_wdata_112,
	local_wdata_48,
	local_wdata_80,
	local_wdata_16,
	local_wdata_113,
	local_wdata_49,
	local_wdata_81,
	local_wdata_17,
	local_wdata_114,
	local_wdata_50,
	local_wdata_82,
	local_wdata_18,
	local_wdata_115,
	local_wdata_51,
	local_wdata_83,
	local_wdata_19,
	local_wdata_116,
	local_wdata_52,
	local_wdata_84,
	local_wdata_20,
	local_wdata_117,
	local_wdata_53,
	local_wdata_85,
	local_wdata_21,
	local_wdata_118,
	local_wdata_54,
	local_wdata_86,
	local_wdata_22,
	local_wdata_119,
	local_wdata_55,
	local_wdata_87,
	local_wdata_23,
	local_wdata_120,
	local_wdata_56,
	local_wdata_88,
	local_wdata_24,
	local_wdata_121,
	local_wdata_57,
	local_wdata_89,
	local_wdata_25,
	local_wdata_122,
	local_wdata_58,
	local_wdata_90,
	local_wdata_26,
	local_wdata_123,
	local_wdata_59,
	local_wdata_91,
	local_wdata_27,
	local_wdata_124,
	local_wdata_60,
	local_wdata_92,
	local_wdata_28,
	local_wdata_125,
	local_wdata_61,
	local_wdata_93,
	local_wdata_29,
	local_wdata_126,
	local_wdata_62,
	local_wdata_94,
	local_wdata_30,
	local_wdata_127,
	local_wdata_63,
	local_wdata_95,
	local_wdata_31)/* synthesis synthesis_greybox=0 */;
output 	q_b_0;
output 	q_b_64;
output 	q_b_1;
output 	q_b_65;
output 	q_b_2;
output 	q_b_66;
output 	q_b_3;
output 	q_b_67;
output 	q_b_4;
output 	q_b_68;
output 	q_b_5;
output 	q_b_69;
output 	q_b_6;
output 	q_b_70;
output 	q_b_7;
output 	q_b_71;
output 	q_b_16;
output 	q_b_80;
output 	q_b_17;
output 	q_b_81;
output 	q_b_18;
output 	q_b_82;
output 	q_b_19;
output 	q_b_83;
output 	q_b_20;
output 	q_b_84;
output 	q_b_21;
output 	q_b_85;
output 	q_b_22;
output 	q_b_86;
output 	q_b_23;
output 	q_b_87;
output 	q_b_32;
output 	q_b_96;
output 	q_b_33;
output 	q_b_97;
output 	q_b_34;
output 	q_b_98;
output 	q_b_35;
output 	q_b_99;
output 	q_b_36;
output 	q_b_100;
output 	q_b_37;
output 	q_b_101;
output 	q_b_38;
output 	q_b_102;
output 	q_b_39;
output 	q_b_103;
output 	q_b_48;
output 	q_b_112;
output 	q_b_49;
output 	q_b_113;
output 	q_b_50;
output 	q_b_114;
output 	q_b_51;
output 	q_b_115;
output 	q_b_52;
output 	q_b_116;
output 	q_b_53;
output 	q_b_117;
output 	q_b_54;
output 	q_b_118;
output 	q_b_55;
output 	q_b_119;
output 	q_b_8;
output 	q_b_72;
output 	q_b_9;
output 	q_b_73;
output 	q_b_10;
output 	q_b_74;
output 	q_b_11;
output 	q_b_75;
output 	q_b_12;
output 	q_b_76;
output 	q_b_13;
output 	q_b_77;
output 	q_b_14;
output 	q_b_78;
output 	q_b_15;
output 	q_b_79;
output 	q_b_24;
output 	q_b_88;
output 	q_b_25;
output 	q_b_89;
output 	q_b_26;
output 	q_b_90;
output 	q_b_27;
output 	q_b_91;
output 	q_b_28;
output 	q_b_92;
output 	q_b_29;
output 	q_b_93;
output 	q_b_30;
output 	q_b_94;
output 	q_b_31;
output 	q_b_95;
output 	q_b_40;
output 	q_b_104;
output 	q_b_41;
output 	q_b_105;
output 	q_b_42;
output 	q_b_106;
output 	q_b_43;
output 	q_b_107;
output 	q_b_44;
output 	q_b_108;
output 	q_b_45;
output 	q_b_109;
output 	q_b_46;
output 	q_b_110;
output 	q_b_47;
output 	q_b_111;
output 	q_b_56;
output 	q_b_120;
output 	q_b_57;
output 	q_b_121;
output 	q_b_58;
output 	q_b_122;
output 	q_b_59;
output 	q_b_123;
output 	q_b_60;
output 	q_b_124;
output 	q_b_61;
output 	q_b_125;
output 	q_b_62;
output 	q_b_126;
output 	q_b_63;
output 	q_b_127;
output 	clk_0;
output 	clk_1;
output 	dataout_0;
output 	dataout_01;
output 	dataout_02;
output 	dataout_03;
output 	dataout_04;
output 	dataout_05;
output 	dataout_06;
output 	dataout_07;
output 	dataout_08;
output 	dataout_09;
output 	dataout_010;
output 	dataout_011;
output 	dataout_012;
output 	dataout_013;
output 	dataout_014;
output 	dataout_015;
output 	dataout_016;
output 	dataout_017;
output 	dataout_018;
output 	dataout_019;
output 	dataout_020;
output 	dataout_021;
output 	dataout_022;
output 	dataout_023;
output 	dqs_delay_ctrl_0;
output 	dqs_delay_ctrl_1;
output 	dqs_delay_ctrl_2;
output 	dqs_delay_ctrl_3;
output 	dqs_delay_ctrl_4;
output 	dqs_delay_ctrl_5;
output 	wire_output_dq_0_output_ddio_out_inst_dataout;
output 	wire_output_dq_0_output_ddio_out_inst_dataout1;
output 	wire_output_dq_0_output_ddio_out_inst_dataout2;
output 	wire_output_dq_0_output_ddio_out_inst_dataout3;
output 	mem_clk_buf_in_0;
output 	mem_clk_n_buf_in_0;
output 	wire_bidir_dq_0_output_ddio_out_inst_dataout;
output 	wire_bidir_dq_1_output_ddio_out_inst_dataout;
output 	wire_bidir_dq_2_output_ddio_out_inst_dataout;
output 	wire_bidir_dq_3_output_ddio_out_inst_dataout;
output 	wire_bidir_dq_4_output_ddio_out_inst_dataout;
output 	wire_bidir_dq_5_output_ddio_out_inst_dataout;
output 	wire_bidir_dq_6_output_ddio_out_inst_dataout;
output 	wire_bidir_dq_7_output_ddio_out_inst_dataout;
output 	wire_bidir_dq_0_output_ddio_out_inst_dataout1;
output 	wire_bidir_dq_1_output_ddio_out_inst_dataout1;
output 	wire_bidir_dq_2_output_ddio_out_inst_dataout1;
output 	wire_bidir_dq_3_output_ddio_out_inst_dataout1;
output 	wire_bidir_dq_4_output_ddio_out_inst_dataout1;
output 	wire_bidir_dq_5_output_ddio_out_inst_dataout1;
output 	wire_bidir_dq_6_output_ddio_out_inst_dataout1;
output 	wire_bidir_dq_7_output_ddio_out_inst_dataout1;
output 	wire_bidir_dq_0_output_ddio_out_inst_dataout2;
output 	wire_bidir_dq_1_output_ddio_out_inst_dataout2;
output 	wire_bidir_dq_2_output_ddio_out_inst_dataout2;
output 	wire_bidir_dq_3_output_ddio_out_inst_dataout2;
output 	wire_bidir_dq_4_output_ddio_out_inst_dataout2;
output 	wire_bidir_dq_5_output_ddio_out_inst_dataout2;
output 	wire_bidir_dq_6_output_ddio_out_inst_dataout2;
output 	wire_bidir_dq_7_output_ddio_out_inst_dataout2;
output 	wire_bidir_dq_0_output_ddio_out_inst_dataout3;
output 	wire_bidir_dq_1_output_ddio_out_inst_dataout3;
output 	wire_bidir_dq_2_output_ddio_out_inst_dataout3;
output 	wire_bidir_dq_3_output_ddio_out_inst_dataout3;
output 	wire_bidir_dq_4_output_ddio_out_inst_dataout3;
output 	wire_bidir_dq_5_output_ddio_out_inst_dataout3;
output 	wire_bidir_dq_6_output_ddio_out_inst_dataout3;
output 	wire_bidir_dq_7_output_ddio_out_inst_dataout3;
output 	dqs_pseudo_diff_out_0;
output 	dqsn_pseudo_diff_out_0;
output 	dqs_pseudo_diff_out_1;
output 	dqsn_pseudo_diff_out_1;
output 	dqs_pseudo_diff_out_2;
output 	dqsn_pseudo_diff_out_2;
output 	dqs_pseudo_diff_out_3;
output 	dqsn_pseudo_diff_out_3;
input 	dq_datain_0;
input 	dq_datain_1;
input 	dq_datain_2;
input 	dq_datain_3;
input 	dq_datain_4;
input 	dq_datain_5;
input 	dq_datain_6;
input 	dq_datain_7;
input 	dq_datain_8;
input 	dq_datain_9;
input 	dq_datain_10;
input 	dq_datain_11;
input 	dq_datain_12;
input 	dq_datain_13;
input 	dq_datain_14;
input 	dq_datain_15;
input 	dq_datain_16;
input 	dq_datain_17;
input 	dq_datain_18;
input 	dq_datain_19;
input 	dq_datain_20;
input 	dq_datain_21;
input 	dq_datain_22;
input 	dq_datain_23;
input 	dq_datain_24;
input 	dq_datain_25;
input 	dq_datain_26;
input 	dq_datain_27;
input 	dq_datain_28;
input 	dq_datain_29;
input 	dq_datain_30;
input 	dq_datain_31;
input 	dqs_buffered_0;
input 	dqs_buffered_1;
input 	dqs_buffered_2;
input 	dqs_buffered_3;
input 	fb_clk;
output 	ready_out;
output 	ctl_rdata_valid_0;
output 	reset_request_n;
output 	int_refresh_ack;
output 	local_init_done;
output 	reset_phy_clk_1x_n;
output 	bidir_dq_0_oe_ff_inst;
output 	bidir_dq_1_oe_ff_inst;
output 	bidir_dq_2_oe_ff_inst;
output 	bidir_dq_3_oe_ff_inst;
output 	bidir_dq_4_oe_ff_inst;
output 	bidir_dq_5_oe_ff_inst;
output 	bidir_dq_6_oe_ff_inst;
output 	bidir_dq_7_oe_ff_inst;
output 	bidir_dq_0_oe_ff_inst1;
output 	bidir_dq_1_oe_ff_inst1;
output 	bidir_dq_2_oe_ff_inst1;
output 	bidir_dq_3_oe_ff_inst1;
output 	bidir_dq_4_oe_ff_inst1;
output 	bidir_dq_5_oe_ff_inst1;
output 	bidir_dq_6_oe_ff_inst1;
output 	bidir_dq_7_oe_ff_inst1;
output 	bidir_dq_0_oe_ff_inst2;
output 	bidir_dq_1_oe_ff_inst2;
output 	bidir_dq_2_oe_ff_inst2;
output 	bidir_dq_3_oe_ff_inst2;
output 	bidir_dq_4_oe_ff_inst2;
output 	bidir_dq_5_oe_ff_inst2;
output 	bidir_dq_6_oe_ff_inst2;
output 	bidir_dq_7_oe_ff_inst2;
output 	bidir_dq_0_oe_ff_inst3;
output 	bidir_dq_1_oe_ff_inst3;
output 	bidir_dq_2_oe_ff_inst3;
output 	bidir_dq_3_oe_ff_inst3;
output 	bidir_dq_4_oe_ff_inst3;
output 	bidir_dq_5_oe_ff_inst3;
output 	bidir_dq_6_oe_ff_inst3;
output 	bidir_dq_7_oe_ff_inst3;
output 	dqs_0_oe_ff_inst;
output 	dqs_0_oe_ff_inst1;
output 	dqs_0_oe_ff_inst2;
output 	dqs_0_oe_ff_inst3;
output 	dqsn_0_oe_ff_inst;
output 	dqsn_0_oe_ff_inst1;
output 	dqsn_0_oe_ff_inst2;
output 	dqsn_0_oe_ff_inst3;
input 	GND_port;
input 	local_size_1;
input 	local_address_0;
input 	local_size_0;
input 	local_size_6;
input 	local_size_5;
input 	local_size_4;
input 	local_size_2;
input 	local_size_3;
input 	local_read_req;
input 	local_write_req;
input 	local_burstbegin;
input 	global_reset_n;
input 	pll_ref_clk;
input 	soft_reset_n;
input 	local_address_8;
input 	local_address_10;
input 	local_address_9;
input 	local_address_23;
input 	local_address_24;
input 	local_address_22;
input 	local_address_20;
input 	local_address_21;
input 	local_address_19;
input 	local_address_17;
input 	local_address_18;
input 	local_address_13;
input 	local_address_11;
input 	local_address_12;
input 	local_address_16;
input 	local_address_14;
input 	local_address_15;
input 	local_address_1;
input 	local_address_2;
input 	local_address_3;
input 	local_address_4;
input 	local_address_5;
input 	local_address_7;
input 	local_address_6;
input 	local_be_4;
input 	local_be_12;
input 	local_be_0;
input 	local_be_8;
input 	local_be_5;
input 	local_be_13;
input 	local_be_1;
input 	local_be_9;
input 	local_be_6;
input 	local_be_14;
input 	local_be_2;
input 	local_be_10;
input 	local_be_7;
input 	local_be_15;
input 	local_be_3;
input 	local_be_11;
input 	local_wdata_96;
input 	local_wdata_32;
input 	local_wdata_64;
input 	local_wdata_0;
input 	local_wdata_97;
input 	local_wdata_33;
input 	local_wdata_65;
input 	local_wdata_1;
input 	local_wdata_98;
input 	local_wdata_34;
input 	local_wdata_66;
input 	local_wdata_2;
input 	local_wdata_99;
input 	local_wdata_35;
input 	local_wdata_67;
input 	local_wdata_3;
input 	local_wdata_100;
input 	local_wdata_36;
input 	local_wdata_68;
input 	local_wdata_4;
input 	local_wdata_101;
input 	local_wdata_37;
input 	local_wdata_69;
input 	local_wdata_5;
input 	local_wdata_102;
input 	local_wdata_38;
input 	local_wdata_70;
input 	local_wdata_6;
input 	local_wdata_103;
input 	local_wdata_39;
input 	local_wdata_71;
input 	local_wdata_7;
input 	local_wdata_104;
input 	local_wdata_40;
input 	local_wdata_72;
input 	local_wdata_8;
input 	local_wdata_105;
input 	local_wdata_41;
input 	local_wdata_73;
input 	local_wdata_9;
input 	local_wdata_106;
input 	local_wdata_42;
input 	local_wdata_74;
input 	local_wdata_10;
input 	local_wdata_107;
input 	local_wdata_43;
input 	local_wdata_75;
input 	local_wdata_11;
input 	local_wdata_108;
input 	local_wdata_44;
input 	local_wdata_76;
input 	local_wdata_12;
input 	local_wdata_109;
input 	local_wdata_45;
input 	local_wdata_77;
input 	local_wdata_13;
input 	local_wdata_110;
input 	local_wdata_46;
input 	local_wdata_78;
input 	local_wdata_14;
input 	local_wdata_111;
input 	local_wdata_47;
input 	local_wdata_79;
input 	local_wdata_15;
input 	local_wdata_112;
input 	local_wdata_48;
input 	local_wdata_80;
input 	local_wdata_16;
input 	local_wdata_113;
input 	local_wdata_49;
input 	local_wdata_81;
input 	local_wdata_17;
input 	local_wdata_114;
input 	local_wdata_50;
input 	local_wdata_82;
input 	local_wdata_18;
input 	local_wdata_115;
input 	local_wdata_51;
input 	local_wdata_83;
input 	local_wdata_19;
input 	local_wdata_116;
input 	local_wdata_52;
input 	local_wdata_84;
input 	local_wdata_20;
input 	local_wdata_117;
input 	local_wdata_53;
input 	local_wdata_85;
input 	local_wdata_21;
input 	local_wdata_118;
input 	local_wdata_54;
input 	local_wdata_86;
input 	local_wdata_22;
input 	local_wdata_119;
input 	local_wdata_55;
input 	local_wdata_87;
input 	local_wdata_23;
input 	local_wdata_120;
input 	local_wdata_56;
input 	local_wdata_88;
input 	local_wdata_24;
input 	local_wdata_121;
input 	local_wdata_57;
input 	local_wdata_89;
input 	local_wdata_25;
input 	local_wdata_122;
input 	local_wdata_58;
input 	local_wdata_90;
input 	local_wdata_26;
input 	local_wdata_123;
input 	local_wdata_59;
input 	local_wdata_91;
input 	local_wdata_27;
input 	local_wdata_124;
input 	local_wdata_60;
input 	local_wdata_92;
input 	local_wdata_28;
input 	local_wdata_125;
input 	local_wdata_61;
input 	local_wdata_93;
input 	local_wdata_29;
input 	local_wdata_126;
input 	local_wdata_62;
input 	local_wdata_94;
input 	local_wdata_30;
input 	local_wdata_127;
input 	local_wdata_63;
input 	local_wdata_95;
input 	local_wdata_31;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|state_machine_inst|do_read_r~q ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[96] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[32] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[64] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[97] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[33] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[65] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[98] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[34] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[66] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[99] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[35] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[67] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[100] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[36] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[68] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[101] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[37] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[69] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[102] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[38] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[70] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[103] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[39] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[71] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[104] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[40] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[72] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[8] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[105] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[41] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[73] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[9] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[106] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[42] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[74] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[10] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[107] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[43] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[75] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[11] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[108] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[44] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[76] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[12] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[109] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[45] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[77] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[13] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[110] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[46] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[78] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[14] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[111] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[47] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[79] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[15] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[112] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[48] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[80] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[16] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[113] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[49] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[81] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[17] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[114] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[50] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[82] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[18] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[115] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[51] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[83] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[19] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[116] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[52] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[84] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[20] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[117] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[53] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[85] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[21] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[118] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[54] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[86] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[22] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[119] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[55] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[87] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[23] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[120] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[56] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[88] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[24] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[121] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[57] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[89] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[25] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[122] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[58] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[90] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[26] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[123] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[59] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[91] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[27] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[124] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[60] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[92] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[28] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[125] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[61] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[93] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[29] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[126] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[62] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[94] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[30] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[127] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[63] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[95] ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[31] ;
wire \ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|ctl_init_fail~q ;
wire \ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|ctl_init_success~q ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|state_machine_inst|rdwr_data_valid_r~q ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|doing_read~q ;
wire \ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|dgrb|wd_lat[2]~q ;
wire \ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|dgrb|wd_lat[1]~q ;
wire \ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|dgrb|wd_lat[0]~q ;
wire \ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|dgrb|wd_lat[3]~q ;
wire \ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|dgrb|wd_lat[4]~q ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_cs_n[1]~0_combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|int_cke_r[0]~q ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[0]~0_combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[1]~1_combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[2]~2_combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[3]~3_combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[4]~4_combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[5]~5_combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[6]~6_combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[7]~7_combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[8]~8_combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[9]~9_combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[10]~10_combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[11]~11_combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[12]~12_combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[13]~13_combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_ba[0]~0_combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_ba[1]~1_combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_ba[2]~2_combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_ras_n[0]~0_combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_cas_n[0]~0_combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_we_n[0]~0_combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[4]~combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[12]~combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[0]~combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[8]~combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[5]~combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[13]~combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[1]~combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[9]~combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[6]~combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[14]~combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[2]~combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[10]~combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[7]~combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[15]~combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[3]~combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[11]~combout ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|int_wdata_valid~q ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|int_dqs_burst~q ;
wire \ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|int_dqs_burst_hr~q ;


ddr3_int_ddr3_int_alt_ddrx_controller_wrapper ddr3_int_alt_ddrx_controller_wrapper_inst(
	.clk_0(clk_0),
	.do_read_r(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|state_machine_inst|do_read_r~q ),
	.q_b_96(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[96] ),
	.q_b_32(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[32] ),
	.q_b_64(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[64] ),
	.q_b_0(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.q_b_97(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[97] ),
	.q_b_33(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[33] ),
	.q_b_65(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[65] ),
	.q_b_1(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_98(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[98] ),
	.q_b_34(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[34] ),
	.q_b_66(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[66] ),
	.q_b_2(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_99(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[99] ),
	.q_b_35(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[35] ),
	.q_b_67(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[67] ),
	.q_b_3(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_100(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[100] ),
	.q_b_36(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[36] ),
	.q_b_68(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[68] ),
	.q_b_4(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_101(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[101] ),
	.q_b_37(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[37] ),
	.q_b_69(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[69] ),
	.q_b_5(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_102(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[102] ),
	.q_b_38(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[38] ),
	.q_b_70(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[70] ),
	.q_b_6(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.q_b_103(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[103] ),
	.q_b_39(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[39] ),
	.q_b_71(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[71] ),
	.q_b_7(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.q_b_104(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[104] ),
	.q_b_40(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[40] ),
	.q_b_72(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[72] ),
	.q_b_8(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.q_b_105(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[105] ),
	.q_b_41(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[41] ),
	.q_b_73(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[73] ),
	.q_b_9(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.q_b_106(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[106] ),
	.q_b_42(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[42] ),
	.q_b_74(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[74] ),
	.q_b_10(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.q_b_107(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[107] ),
	.q_b_43(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[43] ),
	.q_b_75(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[75] ),
	.q_b_11(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.q_b_108(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[108] ),
	.q_b_44(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[44] ),
	.q_b_76(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[76] ),
	.q_b_12(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.q_b_109(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[109] ),
	.q_b_45(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[45] ),
	.q_b_77(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[77] ),
	.q_b_13(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.q_b_110(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[110] ),
	.q_b_46(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[46] ),
	.q_b_78(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[78] ),
	.q_b_14(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.q_b_111(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[111] ),
	.q_b_47(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[47] ),
	.q_b_79(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[79] ),
	.q_b_15(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.q_b_112(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[112] ),
	.q_b_48(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[48] ),
	.q_b_80(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[80] ),
	.q_b_16(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.q_b_113(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[113] ),
	.q_b_49(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[49] ),
	.q_b_81(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[81] ),
	.q_b_17(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.q_b_114(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[114] ),
	.q_b_50(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[50] ),
	.q_b_82(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[82] ),
	.q_b_18(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.q_b_115(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[115] ),
	.q_b_51(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[51] ),
	.q_b_83(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[83] ),
	.q_b_19(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.q_b_116(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[116] ),
	.q_b_52(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[52] ),
	.q_b_84(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[84] ),
	.q_b_20(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.q_b_117(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[117] ),
	.q_b_53(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[53] ),
	.q_b_85(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[85] ),
	.q_b_21(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.q_b_118(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[118] ),
	.q_b_54(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[54] ),
	.q_b_86(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[86] ),
	.q_b_22(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[22] ),
	.q_b_119(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[119] ),
	.q_b_55(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[55] ),
	.q_b_87(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[87] ),
	.q_b_23(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[23] ),
	.q_b_120(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[120] ),
	.q_b_56(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[56] ),
	.q_b_88(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[88] ),
	.q_b_24(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[24] ),
	.q_b_121(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[121] ),
	.q_b_57(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[57] ),
	.q_b_89(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[89] ),
	.q_b_25(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[25] ),
	.q_b_122(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[122] ),
	.q_b_58(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[58] ),
	.q_b_90(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[90] ),
	.q_b_26(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[26] ),
	.q_b_123(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[123] ),
	.q_b_59(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[59] ),
	.q_b_91(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[91] ),
	.q_b_27(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[27] ),
	.q_b_124(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[124] ),
	.q_b_60(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[60] ),
	.q_b_92(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[92] ),
	.q_b_28(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[28] ),
	.q_b_125(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[125] ),
	.q_b_61(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[61] ),
	.q_b_93(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[93] ),
	.q_b_29(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[29] ),
	.q_b_126(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[126] ),
	.q_b_62(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[62] ),
	.q_b_94(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[94] ),
	.q_b_30(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[30] ),
	.q_b_127(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[127] ),
	.q_b_63(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[63] ),
	.q_b_95(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[95] ),
	.q_b_31(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[31] ),
	.ready_out(ready_out),
	.int_refresh_ack(int_refresh_ack),
	.ctl_init_fail(\ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|ctl_init_fail~q ),
	.ctl_init_success(\ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|ctl_init_success~q ),
	.local_init_done(local_init_done),
	.reset_phy_clk_1x_n(reset_phy_clk_1x_n),
	.rdwr_data_valid_r(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|state_machine_inst|rdwr_data_valid_r~q ),
	.doing_read(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|doing_read~q ),
	.wd_lat_2(\ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|dgrb|wd_lat[2]~q ),
	.wd_lat_1(\ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|dgrb|wd_lat[1]~q ),
	.wd_lat_0(\ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|dgrb|wd_lat[0]~q ),
	.wd_lat_3(\ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|dgrb|wd_lat[3]~q ),
	.wd_lat_4(\ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|dgrb|wd_lat[4]~q ),
	.afi_cs_n_1(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_cs_n[1]~0_combout ),
	.int_cke_r_0(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|int_cke_r[0]~q ),
	.afi_addr_0(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[0]~0_combout ),
	.afi_addr_1(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[1]~1_combout ),
	.afi_addr_2(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[2]~2_combout ),
	.afi_addr_3(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[3]~3_combout ),
	.afi_addr_4(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[4]~4_combout ),
	.afi_addr_5(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[5]~5_combout ),
	.afi_addr_6(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[6]~6_combout ),
	.afi_addr_7(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[7]~7_combout ),
	.afi_addr_8(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[8]~8_combout ),
	.afi_addr_9(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[9]~9_combout ),
	.afi_addr_10(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[10]~10_combout ),
	.afi_addr_11(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[11]~11_combout ),
	.afi_addr_12(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[12]~12_combout ),
	.afi_addr_13(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[13]~13_combout ),
	.afi_ba_0(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_ba[0]~0_combout ),
	.afi_ba_1(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_ba[1]~1_combout ),
	.afi_ba_2(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_ba[2]~2_combout ),
	.afi_ras_n_0(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_ras_n[0]~0_combout ),
	.afi_cas_n_0(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_cas_n[0]~0_combout ),
	.afi_we_n_0(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_we_n[0]~0_combout ),
	.afi_dm_4(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[4]~combout ),
	.afi_dm_12(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[12]~combout ),
	.afi_dm_0(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[0]~combout ),
	.afi_dm_8(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[8]~combout ),
	.afi_dm_5(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[5]~combout ),
	.afi_dm_13(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[13]~combout ),
	.afi_dm_1(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[1]~combout ),
	.afi_dm_9(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[9]~combout ),
	.afi_dm_6(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[6]~combout ),
	.afi_dm_14(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[14]~combout ),
	.afi_dm_2(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[2]~combout ),
	.afi_dm_10(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[10]~combout ),
	.afi_dm_7(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[7]~combout ),
	.afi_dm_15(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[15]~combout ),
	.afi_dm_3(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[3]~combout ),
	.afi_dm_11(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[11]~combout ),
	.int_wdata_valid(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|int_wdata_valid~q ),
	.int_dqs_burst(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|int_dqs_burst~q ),
	.int_dqs_burst_hr(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|int_dqs_burst_hr~q ),
	.GND_port(GND_port),
	.local_size_1(local_size_1),
	.local_address_0(local_address_0),
	.local_size_0(local_size_0),
	.local_size_6(local_size_6),
	.local_size_5(local_size_5),
	.local_size_4(local_size_4),
	.local_size_2(local_size_2),
	.local_size_3(local_size_3),
	.local_read_req(local_read_req),
	.local_write_req(local_write_req),
	.local_burstbegin(local_burstbegin),
	.local_address_8(local_address_8),
	.local_address_10(local_address_10),
	.local_address_9(local_address_9),
	.local_address_23(local_address_23),
	.local_address_24(local_address_24),
	.local_address_22(local_address_22),
	.local_address_20(local_address_20),
	.local_address_21(local_address_21),
	.local_address_19(local_address_19),
	.local_address_17(local_address_17),
	.local_address_18(local_address_18),
	.local_address_13(local_address_13),
	.local_address_11(local_address_11),
	.local_address_12(local_address_12),
	.local_address_16(local_address_16),
	.local_address_14(local_address_14),
	.local_address_15(local_address_15),
	.local_address_1(local_address_1),
	.local_address_2(local_address_2),
	.local_address_3(local_address_3),
	.local_address_4(local_address_4),
	.local_address_5(local_address_5),
	.local_address_7(local_address_7),
	.local_address_6(local_address_6),
	.local_be_4(local_be_4),
	.local_be_12(local_be_12),
	.local_be_0(local_be_0),
	.local_be_8(local_be_8),
	.local_be_5(local_be_5),
	.local_be_13(local_be_13),
	.local_be_1(local_be_1),
	.local_be_9(local_be_9),
	.local_be_6(local_be_6),
	.local_be_14(local_be_14),
	.local_be_2(local_be_2),
	.local_be_10(local_be_10),
	.local_be_7(local_be_7),
	.local_be_15(local_be_15),
	.local_be_3(local_be_3),
	.local_be_11(local_be_11),
	.local_wdata_96(local_wdata_96),
	.local_wdata_32(local_wdata_32),
	.local_wdata_64(local_wdata_64),
	.local_wdata_0(local_wdata_0),
	.local_wdata_97(local_wdata_97),
	.local_wdata_33(local_wdata_33),
	.local_wdata_65(local_wdata_65),
	.local_wdata_1(local_wdata_1),
	.local_wdata_98(local_wdata_98),
	.local_wdata_34(local_wdata_34),
	.local_wdata_66(local_wdata_66),
	.local_wdata_2(local_wdata_2),
	.local_wdata_99(local_wdata_99),
	.local_wdata_35(local_wdata_35),
	.local_wdata_67(local_wdata_67),
	.local_wdata_3(local_wdata_3),
	.local_wdata_100(local_wdata_100),
	.local_wdata_36(local_wdata_36),
	.local_wdata_68(local_wdata_68),
	.local_wdata_4(local_wdata_4),
	.local_wdata_101(local_wdata_101),
	.local_wdata_37(local_wdata_37),
	.local_wdata_69(local_wdata_69),
	.local_wdata_5(local_wdata_5),
	.local_wdata_102(local_wdata_102),
	.local_wdata_38(local_wdata_38),
	.local_wdata_70(local_wdata_70),
	.local_wdata_6(local_wdata_6),
	.local_wdata_103(local_wdata_103),
	.local_wdata_39(local_wdata_39),
	.local_wdata_71(local_wdata_71),
	.local_wdata_7(local_wdata_7),
	.local_wdata_104(local_wdata_104),
	.local_wdata_40(local_wdata_40),
	.local_wdata_72(local_wdata_72),
	.local_wdata_8(local_wdata_8),
	.local_wdata_105(local_wdata_105),
	.local_wdata_41(local_wdata_41),
	.local_wdata_73(local_wdata_73),
	.local_wdata_9(local_wdata_9),
	.local_wdata_106(local_wdata_106),
	.local_wdata_42(local_wdata_42),
	.local_wdata_74(local_wdata_74),
	.local_wdata_10(local_wdata_10),
	.local_wdata_107(local_wdata_107),
	.local_wdata_43(local_wdata_43),
	.local_wdata_75(local_wdata_75),
	.local_wdata_11(local_wdata_11),
	.local_wdata_108(local_wdata_108),
	.local_wdata_44(local_wdata_44),
	.local_wdata_76(local_wdata_76),
	.local_wdata_12(local_wdata_12),
	.local_wdata_109(local_wdata_109),
	.local_wdata_45(local_wdata_45),
	.local_wdata_77(local_wdata_77),
	.local_wdata_13(local_wdata_13),
	.local_wdata_110(local_wdata_110),
	.local_wdata_46(local_wdata_46),
	.local_wdata_78(local_wdata_78),
	.local_wdata_14(local_wdata_14),
	.local_wdata_111(local_wdata_111),
	.local_wdata_47(local_wdata_47),
	.local_wdata_79(local_wdata_79),
	.local_wdata_15(local_wdata_15),
	.local_wdata_112(local_wdata_112),
	.local_wdata_48(local_wdata_48),
	.local_wdata_80(local_wdata_80),
	.local_wdata_16(local_wdata_16),
	.local_wdata_113(local_wdata_113),
	.local_wdata_49(local_wdata_49),
	.local_wdata_81(local_wdata_81),
	.local_wdata_17(local_wdata_17),
	.local_wdata_114(local_wdata_114),
	.local_wdata_50(local_wdata_50),
	.local_wdata_82(local_wdata_82),
	.local_wdata_18(local_wdata_18),
	.local_wdata_115(local_wdata_115),
	.local_wdata_51(local_wdata_51),
	.local_wdata_83(local_wdata_83),
	.local_wdata_19(local_wdata_19),
	.local_wdata_116(local_wdata_116),
	.local_wdata_52(local_wdata_52),
	.local_wdata_84(local_wdata_84),
	.local_wdata_20(local_wdata_20),
	.local_wdata_117(local_wdata_117),
	.local_wdata_53(local_wdata_53),
	.local_wdata_85(local_wdata_85),
	.local_wdata_21(local_wdata_21),
	.local_wdata_118(local_wdata_118),
	.local_wdata_54(local_wdata_54),
	.local_wdata_86(local_wdata_86),
	.local_wdata_22(local_wdata_22),
	.local_wdata_119(local_wdata_119),
	.local_wdata_55(local_wdata_55),
	.local_wdata_87(local_wdata_87),
	.local_wdata_23(local_wdata_23),
	.local_wdata_120(local_wdata_120),
	.local_wdata_56(local_wdata_56),
	.local_wdata_88(local_wdata_88),
	.local_wdata_24(local_wdata_24),
	.local_wdata_121(local_wdata_121),
	.local_wdata_57(local_wdata_57),
	.local_wdata_89(local_wdata_89),
	.local_wdata_25(local_wdata_25),
	.local_wdata_122(local_wdata_122),
	.local_wdata_58(local_wdata_58),
	.local_wdata_90(local_wdata_90),
	.local_wdata_26(local_wdata_26),
	.local_wdata_123(local_wdata_123),
	.local_wdata_59(local_wdata_59),
	.local_wdata_91(local_wdata_91),
	.local_wdata_27(local_wdata_27),
	.local_wdata_124(local_wdata_124),
	.local_wdata_60(local_wdata_60),
	.local_wdata_92(local_wdata_92),
	.local_wdata_28(local_wdata_28),
	.local_wdata_125(local_wdata_125),
	.local_wdata_61(local_wdata_61),
	.local_wdata_93(local_wdata_93),
	.local_wdata_29(local_wdata_29),
	.local_wdata_126(local_wdata_126),
	.local_wdata_62(local_wdata_62),
	.local_wdata_94(local_wdata_94),
	.local_wdata_30(local_wdata_30),
	.local_wdata_127(local_wdata_127),
	.local_wdata_63(local_wdata_63),
	.local_wdata_95(local_wdata_95),
	.local_wdata_31(local_wdata_31));

ddr3_int_ddr3_int_phy ddr3_int_phy_inst(
	.q_b_0(q_b_0),
	.q_b_64(q_b_64),
	.q_b_1(q_b_1),
	.q_b_65(q_b_65),
	.q_b_2(q_b_2),
	.q_b_66(q_b_66),
	.q_b_3(q_b_3),
	.q_b_67(q_b_67),
	.q_b_4(q_b_4),
	.q_b_68(q_b_68),
	.q_b_5(q_b_5),
	.q_b_69(q_b_69),
	.q_b_6(q_b_6),
	.q_b_70(q_b_70),
	.q_b_7(q_b_7),
	.q_b_71(q_b_71),
	.q_b_16(q_b_16),
	.q_b_80(q_b_80),
	.q_b_17(q_b_17),
	.q_b_81(q_b_81),
	.q_b_18(q_b_18),
	.q_b_82(q_b_82),
	.q_b_19(q_b_19),
	.q_b_83(q_b_83),
	.q_b_20(q_b_20),
	.q_b_84(q_b_84),
	.q_b_21(q_b_21),
	.q_b_85(q_b_85),
	.q_b_22(q_b_22),
	.q_b_86(q_b_86),
	.q_b_23(q_b_23),
	.q_b_87(q_b_87),
	.q_b_32(q_b_32),
	.q_b_96(q_b_96),
	.q_b_33(q_b_33),
	.q_b_97(q_b_97),
	.q_b_34(q_b_34),
	.q_b_98(q_b_98),
	.q_b_35(q_b_35),
	.q_b_99(q_b_99),
	.q_b_36(q_b_36),
	.q_b_100(q_b_100),
	.q_b_37(q_b_37),
	.q_b_101(q_b_101),
	.q_b_38(q_b_38),
	.q_b_102(q_b_102),
	.q_b_39(q_b_39),
	.q_b_103(q_b_103),
	.q_b_48(q_b_48),
	.q_b_112(q_b_112),
	.q_b_49(q_b_49),
	.q_b_113(q_b_113),
	.q_b_50(q_b_50),
	.q_b_114(q_b_114),
	.q_b_51(q_b_51),
	.q_b_115(q_b_115),
	.q_b_52(q_b_52),
	.q_b_116(q_b_116),
	.q_b_53(q_b_53),
	.q_b_117(q_b_117),
	.q_b_54(q_b_54),
	.q_b_118(q_b_118),
	.q_b_55(q_b_55),
	.q_b_119(q_b_119),
	.q_b_8(q_b_8),
	.q_b_72(q_b_72),
	.q_b_9(q_b_9),
	.q_b_73(q_b_73),
	.q_b_10(q_b_10),
	.q_b_74(q_b_74),
	.q_b_11(q_b_11),
	.q_b_75(q_b_75),
	.q_b_12(q_b_12),
	.q_b_76(q_b_76),
	.q_b_13(q_b_13),
	.q_b_77(q_b_77),
	.q_b_14(q_b_14),
	.q_b_78(q_b_78),
	.q_b_15(q_b_15),
	.q_b_79(q_b_79),
	.q_b_24(q_b_24),
	.q_b_88(q_b_88),
	.q_b_25(q_b_25),
	.q_b_89(q_b_89),
	.q_b_26(q_b_26),
	.q_b_90(q_b_90),
	.q_b_27(q_b_27),
	.q_b_91(q_b_91),
	.q_b_28(q_b_28),
	.q_b_92(q_b_92),
	.q_b_29(q_b_29),
	.q_b_93(q_b_93),
	.q_b_30(q_b_30),
	.q_b_94(q_b_94),
	.q_b_31(q_b_31),
	.q_b_95(q_b_95),
	.q_b_40(q_b_40),
	.q_b_104(q_b_104),
	.q_b_41(q_b_41),
	.q_b_105(q_b_105),
	.q_b_42(q_b_42),
	.q_b_106(q_b_106),
	.q_b_43(q_b_43),
	.q_b_107(q_b_107),
	.q_b_44(q_b_44),
	.q_b_108(q_b_108),
	.q_b_45(q_b_45),
	.q_b_109(q_b_109),
	.q_b_46(q_b_46),
	.q_b_110(q_b_110),
	.q_b_47(q_b_47),
	.q_b_111(q_b_111),
	.q_b_56(q_b_56),
	.q_b_120(q_b_120),
	.q_b_57(q_b_57),
	.q_b_121(q_b_121),
	.q_b_58(q_b_58),
	.q_b_122(q_b_122),
	.q_b_59(q_b_59),
	.q_b_123(q_b_123),
	.q_b_60(q_b_60),
	.q_b_124(q_b_124),
	.q_b_61(q_b_61),
	.q_b_125(q_b_125),
	.q_b_62(q_b_62),
	.q_b_126(q_b_126),
	.q_b_63(q_b_63),
	.q_b_127(q_b_127),
	.clk_0(clk_0),
	.clk_1(clk_1),
	.dataout_0(dataout_0),
	.dataout_01(dataout_01),
	.dataout_02(dataout_02),
	.dataout_03(dataout_03),
	.dataout_04(dataout_04),
	.dataout_05(dataout_05),
	.dataout_06(dataout_06),
	.dataout_07(dataout_07),
	.dataout_08(dataout_08),
	.dataout_09(dataout_09),
	.dataout_010(dataout_010),
	.dataout_011(dataout_011),
	.dataout_012(dataout_012),
	.dataout_013(dataout_013),
	.dataout_014(dataout_014),
	.dataout_015(dataout_015),
	.dataout_016(dataout_016),
	.dataout_017(dataout_017),
	.dataout_018(dataout_018),
	.dataout_019(dataout_019),
	.dataout_020(dataout_020),
	.dataout_021(dataout_021),
	.dataout_022(dataout_022),
	.dataout_023(dataout_023),
	.dqs_delay_ctrl_0(dqs_delay_ctrl_0),
	.dqs_delay_ctrl_1(dqs_delay_ctrl_1),
	.dqs_delay_ctrl_2(dqs_delay_ctrl_2),
	.dqs_delay_ctrl_3(dqs_delay_ctrl_3),
	.dqs_delay_ctrl_4(dqs_delay_ctrl_4),
	.dqs_delay_ctrl_5(dqs_delay_ctrl_5),
	.wire_output_dq_0_output_ddio_out_inst_dataout(wire_output_dq_0_output_ddio_out_inst_dataout),
	.wire_output_dq_0_output_ddio_out_inst_dataout1(wire_output_dq_0_output_ddio_out_inst_dataout1),
	.wire_output_dq_0_output_ddio_out_inst_dataout2(wire_output_dq_0_output_ddio_out_inst_dataout2),
	.wire_output_dq_0_output_ddio_out_inst_dataout3(wire_output_dq_0_output_ddio_out_inst_dataout3),
	.do_read_r(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|state_machine_inst|do_read_r~q ),
	.mem_clk_buf_in_0(mem_clk_buf_in_0),
	.mem_clk_n_buf_in_0(mem_clk_n_buf_in_0),
	.wire_bidir_dq_0_output_ddio_out_inst_dataout(wire_bidir_dq_0_output_ddio_out_inst_dataout),
	.wire_bidir_dq_1_output_ddio_out_inst_dataout(wire_bidir_dq_1_output_ddio_out_inst_dataout),
	.wire_bidir_dq_2_output_ddio_out_inst_dataout(wire_bidir_dq_2_output_ddio_out_inst_dataout),
	.wire_bidir_dq_3_output_ddio_out_inst_dataout(wire_bidir_dq_3_output_ddio_out_inst_dataout),
	.wire_bidir_dq_4_output_ddio_out_inst_dataout(wire_bidir_dq_4_output_ddio_out_inst_dataout),
	.wire_bidir_dq_5_output_ddio_out_inst_dataout(wire_bidir_dq_5_output_ddio_out_inst_dataout),
	.wire_bidir_dq_6_output_ddio_out_inst_dataout(wire_bidir_dq_6_output_ddio_out_inst_dataout),
	.wire_bidir_dq_7_output_ddio_out_inst_dataout(wire_bidir_dq_7_output_ddio_out_inst_dataout),
	.wire_bidir_dq_0_output_ddio_out_inst_dataout1(wire_bidir_dq_0_output_ddio_out_inst_dataout1),
	.wire_bidir_dq_1_output_ddio_out_inst_dataout1(wire_bidir_dq_1_output_ddio_out_inst_dataout1),
	.wire_bidir_dq_2_output_ddio_out_inst_dataout1(wire_bidir_dq_2_output_ddio_out_inst_dataout1),
	.wire_bidir_dq_3_output_ddio_out_inst_dataout1(wire_bidir_dq_3_output_ddio_out_inst_dataout1),
	.wire_bidir_dq_4_output_ddio_out_inst_dataout1(wire_bidir_dq_4_output_ddio_out_inst_dataout1),
	.wire_bidir_dq_5_output_ddio_out_inst_dataout1(wire_bidir_dq_5_output_ddio_out_inst_dataout1),
	.wire_bidir_dq_6_output_ddio_out_inst_dataout1(wire_bidir_dq_6_output_ddio_out_inst_dataout1),
	.wire_bidir_dq_7_output_ddio_out_inst_dataout1(wire_bidir_dq_7_output_ddio_out_inst_dataout1),
	.wire_bidir_dq_0_output_ddio_out_inst_dataout2(wire_bidir_dq_0_output_ddio_out_inst_dataout2),
	.wire_bidir_dq_1_output_ddio_out_inst_dataout2(wire_bidir_dq_1_output_ddio_out_inst_dataout2),
	.wire_bidir_dq_2_output_ddio_out_inst_dataout2(wire_bidir_dq_2_output_ddio_out_inst_dataout2),
	.wire_bidir_dq_3_output_ddio_out_inst_dataout2(wire_bidir_dq_3_output_ddio_out_inst_dataout2),
	.wire_bidir_dq_4_output_ddio_out_inst_dataout2(wire_bidir_dq_4_output_ddio_out_inst_dataout2),
	.wire_bidir_dq_5_output_ddio_out_inst_dataout2(wire_bidir_dq_5_output_ddio_out_inst_dataout2),
	.wire_bidir_dq_6_output_ddio_out_inst_dataout2(wire_bidir_dq_6_output_ddio_out_inst_dataout2),
	.wire_bidir_dq_7_output_ddio_out_inst_dataout2(wire_bidir_dq_7_output_ddio_out_inst_dataout2),
	.wire_bidir_dq_0_output_ddio_out_inst_dataout3(wire_bidir_dq_0_output_ddio_out_inst_dataout3),
	.wire_bidir_dq_1_output_ddio_out_inst_dataout3(wire_bidir_dq_1_output_ddio_out_inst_dataout3),
	.wire_bidir_dq_2_output_ddio_out_inst_dataout3(wire_bidir_dq_2_output_ddio_out_inst_dataout3),
	.wire_bidir_dq_3_output_ddio_out_inst_dataout3(wire_bidir_dq_3_output_ddio_out_inst_dataout3),
	.wire_bidir_dq_4_output_ddio_out_inst_dataout3(wire_bidir_dq_4_output_ddio_out_inst_dataout3),
	.wire_bidir_dq_5_output_ddio_out_inst_dataout3(wire_bidir_dq_5_output_ddio_out_inst_dataout3),
	.wire_bidir_dq_6_output_ddio_out_inst_dataout3(wire_bidir_dq_6_output_ddio_out_inst_dataout3),
	.wire_bidir_dq_7_output_ddio_out_inst_dataout3(wire_bidir_dq_7_output_ddio_out_inst_dataout3),
	.dqs_pseudo_diff_out_0(dqs_pseudo_diff_out_0),
	.dqsn_pseudo_diff_out_0(dqsn_pseudo_diff_out_0),
	.dqs_pseudo_diff_out_1(dqs_pseudo_diff_out_1),
	.dqsn_pseudo_diff_out_1(dqsn_pseudo_diff_out_1),
	.dqs_pseudo_diff_out_2(dqs_pseudo_diff_out_2),
	.dqsn_pseudo_diff_out_2(dqsn_pseudo_diff_out_2),
	.dqs_pseudo_diff_out_3(dqs_pseudo_diff_out_3),
	.dqsn_pseudo_diff_out_3(dqsn_pseudo_diff_out_3),
	.dq_datain_0(dq_datain_0),
	.dq_datain_1(dq_datain_1),
	.dq_datain_2(dq_datain_2),
	.dq_datain_3(dq_datain_3),
	.dq_datain_4(dq_datain_4),
	.dq_datain_5(dq_datain_5),
	.dq_datain_6(dq_datain_6),
	.dq_datain_7(dq_datain_7),
	.dq_datain_8(dq_datain_8),
	.dq_datain_9(dq_datain_9),
	.dq_datain_10(dq_datain_10),
	.dq_datain_11(dq_datain_11),
	.dq_datain_12(dq_datain_12),
	.dq_datain_13(dq_datain_13),
	.dq_datain_14(dq_datain_14),
	.dq_datain_15(dq_datain_15),
	.dq_datain_16(dq_datain_16),
	.dq_datain_17(dq_datain_17),
	.dq_datain_18(dq_datain_18),
	.dq_datain_19(dq_datain_19),
	.dq_datain_20(dq_datain_20),
	.dq_datain_21(dq_datain_21),
	.dq_datain_22(dq_datain_22),
	.dq_datain_23(dq_datain_23),
	.dq_datain_24(dq_datain_24),
	.dq_datain_25(dq_datain_25),
	.dq_datain_26(dq_datain_26),
	.dq_datain_27(dq_datain_27),
	.dq_datain_28(dq_datain_28),
	.dq_datain_29(dq_datain_29),
	.dq_datain_30(dq_datain_30),
	.dq_datain_31(dq_datain_31),
	.dqs_buffered_0(dqs_buffered_0),
	.dqs_buffered_1(dqs_buffered_1),
	.dqs_buffered_2(dqs_buffered_2),
	.dqs_buffered_3(dqs_buffered_3),
	.q_b_961(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[96] ),
	.q_b_321(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[32] ),
	.q_b_641(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[64] ),
	.q_b_01(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.q_b_971(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[97] ),
	.q_b_331(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[33] ),
	.q_b_651(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[65] ),
	.q_b_128(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_981(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[98] ),
	.q_b_341(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[34] ),
	.q_b_661(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[66] ),
	.q_b_210(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_991(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[99] ),
	.q_b_351(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[35] ),
	.q_b_671(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[67] ),
	.q_b_310(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_1001(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[100] ),
	.q_b_361(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[36] ),
	.q_b_681(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[68] ),
	.q_b_410(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.q_b_1011(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[101] ),
	.q_b_371(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[37] ),
	.q_b_691(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[69] ),
	.q_b_510(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_1021(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[102] ),
	.q_b_381(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[38] ),
	.q_b_701(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[70] ),
	.q_b_610(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.q_b_1031(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[103] ),
	.q_b_391(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[39] ),
	.q_b_711(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[71] ),
	.q_b_710(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.q_b_1041(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[104] ),
	.q_b_401(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[40] ),
	.q_b_721(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[72] ),
	.q_b_810(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[8] ),
	.q_b_1051(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[105] ),
	.q_b_411(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[41] ),
	.q_b_731(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[73] ),
	.q_b_910(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[9] ),
	.q_b_1061(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[106] ),
	.q_b_421(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[42] ),
	.q_b_741(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[74] ),
	.q_b_1010(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[10] ),
	.q_b_1071(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[107] ),
	.q_b_431(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[43] ),
	.q_b_751(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[75] ),
	.q_b_1110(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[11] ),
	.q_b_1081(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[108] ),
	.q_b_441(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[44] ),
	.q_b_761(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[76] ),
	.q_b_129(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[12] ),
	.q_b_1091(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[109] ),
	.q_b_451(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[45] ),
	.q_b_771(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[77] ),
	.q_b_131(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[13] ),
	.q_b_1101(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[110] ),
	.q_b_461(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[46] ),
	.q_b_781(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[78] ),
	.q_b_141(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[14] ),
	.q_b_1111(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[111] ),
	.q_b_471(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[47] ),
	.q_b_791(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[79] ),
	.q_b_151(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[15] ),
	.q_b_1121(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[112] ),
	.q_b_481(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[48] ),
	.q_b_801(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[80] ),
	.q_b_161(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[16] ),
	.q_b_1131(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[113] ),
	.q_b_491(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[49] ),
	.q_b_811(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[81] ),
	.q_b_171(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[17] ),
	.q_b_1141(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[114] ),
	.q_b_501(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[50] ),
	.q_b_821(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[82] ),
	.q_b_181(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[18] ),
	.q_b_1151(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[115] ),
	.q_b_511(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[51] ),
	.q_b_831(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[83] ),
	.q_b_191(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[19] ),
	.q_b_1161(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[116] ),
	.q_b_521(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[52] ),
	.q_b_841(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[84] ),
	.q_b_201(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[20] ),
	.q_b_1171(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[117] ),
	.q_b_531(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[53] ),
	.q_b_851(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[85] ),
	.q_b_211(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[21] ),
	.q_b_1181(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[118] ),
	.q_b_541(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[54] ),
	.q_b_861(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[86] ),
	.q_b_221(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[22] ),
	.q_b_1191(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[119] ),
	.q_b_551(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[55] ),
	.q_b_871(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[87] ),
	.q_b_231(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[23] ),
	.q_b_1201(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[120] ),
	.q_b_561(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[56] ),
	.q_b_881(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[88] ),
	.q_b_241(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[24] ),
	.q_b_1211(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[121] ),
	.q_b_571(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[57] ),
	.q_b_891(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[89] ),
	.q_b_251(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[25] ),
	.q_b_1221(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[122] ),
	.q_b_581(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[58] ),
	.q_b_901(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[90] ),
	.q_b_261(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[26] ),
	.q_b_1231(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[123] ),
	.q_b_591(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[59] ),
	.q_b_911(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[91] ),
	.q_b_271(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[27] ),
	.q_b_1241(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[124] ),
	.q_b_601(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[60] ),
	.q_b_921(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[92] ),
	.q_b_281(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[28] ),
	.q_b_1251(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[125] ),
	.q_b_611(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[61] ),
	.q_b_931(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[93] ),
	.q_b_291(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[29] ),
	.q_b_1261(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[126] ),
	.q_b_621(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[62] ),
	.q_b_941(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[94] ),
	.q_b_301(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[30] ),
	.q_b_1271(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[127] ),
	.q_b_631(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[63] ),
	.q_b_951(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[95] ),
	.q_b_311(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[31] ),
	.fb_clk(fb_clk),
	.ctl_rdata_valid_0(ctl_rdata_valid_0),
	.reset_request_n(reset_request_n),
	.ctl_init_fail(\ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|ctl_init_fail~q ),
	.ctl_init_success(\ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|ctl_init_success~q ),
	.reset_phy_clk_1x_n(reset_phy_clk_1x_n),
	.rdwr_data_valid_r(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|state_machine_inst|rdwr_data_valid_r~q ),
	.doing_read(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|doing_read~q ),
	.bidir_dq_0_oe_ff_inst(bidir_dq_0_oe_ff_inst),
	.bidir_dq_1_oe_ff_inst(bidir_dq_1_oe_ff_inst),
	.bidir_dq_2_oe_ff_inst(bidir_dq_2_oe_ff_inst),
	.bidir_dq_3_oe_ff_inst(bidir_dq_3_oe_ff_inst),
	.bidir_dq_4_oe_ff_inst(bidir_dq_4_oe_ff_inst),
	.bidir_dq_5_oe_ff_inst(bidir_dq_5_oe_ff_inst),
	.bidir_dq_6_oe_ff_inst(bidir_dq_6_oe_ff_inst),
	.bidir_dq_7_oe_ff_inst(bidir_dq_7_oe_ff_inst),
	.bidir_dq_0_oe_ff_inst1(bidir_dq_0_oe_ff_inst1),
	.bidir_dq_1_oe_ff_inst1(bidir_dq_1_oe_ff_inst1),
	.bidir_dq_2_oe_ff_inst1(bidir_dq_2_oe_ff_inst1),
	.bidir_dq_3_oe_ff_inst1(bidir_dq_3_oe_ff_inst1),
	.bidir_dq_4_oe_ff_inst1(bidir_dq_4_oe_ff_inst1),
	.bidir_dq_5_oe_ff_inst1(bidir_dq_5_oe_ff_inst1),
	.bidir_dq_6_oe_ff_inst1(bidir_dq_6_oe_ff_inst1),
	.bidir_dq_7_oe_ff_inst1(bidir_dq_7_oe_ff_inst1),
	.bidir_dq_0_oe_ff_inst2(bidir_dq_0_oe_ff_inst2),
	.bidir_dq_1_oe_ff_inst2(bidir_dq_1_oe_ff_inst2),
	.bidir_dq_2_oe_ff_inst2(bidir_dq_2_oe_ff_inst2),
	.bidir_dq_3_oe_ff_inst2(bidir_dq_3_oe_ff_inst2),
	.bidir_dq_4_oe_ff_inst2(bidir_dq_4_oe_ff_inst2),
	.bidir_dq_5_oe_ff_inst2(bidir_dq_5_oe_ff_inst2),
	.bidir_dq_6_oe_ff_inst2(bidir_dq_6_oe_ff_inst2),
	.bidir_dq_7_oe_ff_inst2(bidir_dq_7_oe_ff_inst2),
	.bidir_dq_0_oe_ff_inst3(bidir_dq_0_oe_ff_inst3),
	.bidir_dq_1_oe_ff_inst3(bidir_dq_1_oe_ff_inst3),
	.bidir_dq_2_oe_ff_inst3(bidir_dq_2_oe_ff_inst3),
	.bidir_dq_3_oe_ff_inst3(bidir_dq_3_oe_ff_inst3),
	.bidir_dq_4_oe_ff_inst3(bidir_dq_4_oe_ff_inst3),
	.bidir_dq_5_oe_ff_inst3(bidir_dq_5_oe_ff_inst3),
	.bidir_dq_6_oe_ff_inst3(bidir_dq_6_oe_ff_inst3),
	.bidir_dq_7_oe_ff_inst3(bidir_dq_7_oe_ff_inst3),
	.dqs_0_oe_ff_inst(dqs_0_oe_ff_inst),
	.dqs_0_oe_ff_inst1(dqs_0_oe_ff_inst1),
	.dqs_0_oe_ff_inst2(dqs_0_oe_ff_inst2),
	.dqs_0_oe_ff_inst3(dqs_0_oe_ff_inst3),
	.dqsn_0_oe_ff_inst(dqsn_0_oe_ff_inst),
	.dqsn_0_oe_ff_inst1(dqsn_0_oe_ff_inst1),
	.dqsn_0_oe_ff_inst2(dqsn_0_oe_ff_inst2),
	.dqsn_0_oe_ff_inst3(dqsn_0_oe_ff_inst3),
	.wd_lat_2(\ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|dgrb|wd_lat[2]~q ),
	.wd_lat_1(\ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|dgrb|wd_lat[1]~q ),
	.wd_lat_0(\ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|dgrb|wd_lat[0]~q ),
	.wd_lat_3(\ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|dgrb|wd_lat[3]~q ),
	.wd_lat_4(\ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy_inst|seq_wrapper|seq_inst|dgrb|wd_lat[4]~q ),
	.afi_cs_n_1(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_cs_n[1]~0_combout ),
	.int_cke_r_0(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|int_cke_r[0]~q ),
	.afi_addr_0(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[0]~0_combout ),
	.afi_addr_1(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[1]~1_combout ),
	.afi_addr_2(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[2]~2_combout ),
	.afi_addr_3(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[3]~3_combout ),
	.afi_addr_4(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[4]~4_combout ),
	.afi_addr_5(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[5]~5_combout ),
	.afi_addr_6(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[6]~6_combout ),
	.afi_addr_7(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[7]~7_combout ),
	.afi_addr_8(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[8]~8_combout ),
	.afi_addr_9(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[9]~9_combout ),
	.afi_addr_10(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[10]~10_combout ),
	.afi_addr_11(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[11]~11_combout ),
	.afi_addr_12(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[12]~12_combout ),
	.afi_addr_13(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_addr[13]~13_combout ),
	.afi_ba_0(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_ba[0]~0_combout ),
	.afi_ba_1(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_ba[1]~1_combout ),
	.afi_ba_2(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_ba[2]~2_combout ),
	.afi_ras_n_0(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_ras_n[0]~0_combout ),
	.afi_cas_n_0(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_cas_n[0]~0_combout ),
	.afi_we_n_0(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|addr_cmd_inst|afi_we_n[0]~0_combout ),
	.afi_dm_4(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[4]~combout ),
	.afi_dm_12(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[12]~combout ),
	.afi_dm_0(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[0]~combout ),
	.afi_dm_8(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[8]~combout ),
	.afi_dm_5(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[5]~combout ),
	.afi_dm_13(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[13]~combout ),
	.afi_dm_1(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[1]~combout ),
	.afi_dm_9(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[9]~combout ),
	.afi_dm_6(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[6]~combout ),
	.afi_dm_14(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[14]~combout ),
	.afi_dm_2(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[2]~combout ),
	.afi_dm_10(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[10]~combout ),
	.afi_dm_7(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[7]~combout ),
	.afi_dm_15(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[15]~combout ),
	.afi_dm_3(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[3]~combout ),
	.afi_dm_11(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|afi_dm[11]~combout ),
	.int_wdata_valid(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|int_wdata_valid~q ),
	.int_dqs_burst(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|int_dqs_burst~q ),
	.int_dqs_burst_hr(\ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller_inst|afi_block_inst|int_dqs_burst_hr~q ),
	.GND_port(GND_port),
	.global_reset_n(global_reset_n),
	.pll_ref_clk(pll_ref_clk),
	.soft_reset_n(soft_reset_n));

endmodule

module ddr3_int_ddr3_int_alt_ddrx_controller_wrapper (
	clk_0,
	do_read_r,
	q_b_96,
	q_b_32,
	q_b_64,
	q_b_0,
	q_b_97,
	q_b_33,
	q_b_65,
	q_b_1,
	q_b_98,
	q_b_34,
	q_b_66,
	q_b_2,
	q_b_99,
	q_b_35,
	q_b_67,
	q_b_3,
	q_b_100,
	q_b_36,
	q_b_68,
	q_b_4,
	q_b_101,
	q_b_37,
	q_b_69,
	q_b_5,
	q_b_102,
	q_b_38,
	q_b_70,
	q_b_6,
	q_b_103,
	q_b_39,
	q_b_71,
	q_b_7,
	q_b_104,
	q_b_40,
	q_b_72,
	q_b_8,
	q_b_105,
	q_b_41,
	q_b_73,
	q_b_9,
	q_b_106,
	q_b_42,
	q_b_74,
	q_b_10,
	q_b_107,
	q_b_43,
	q_b_75,
	q_b_11,
	q_b_108,
	q_b_44,
	q_b_76,
	q_b_12,
	q_b_109,
	q_b_45,
	q_b_77,
	q_b_13,
	q_b_110,
	q_b_46,
	q_b_78,
	q_b_14,
	q_b_111,
	q_b_47,
	q_b_79,
	q_b_15,
	q_b_112,
	q_b_48,
	q_b_80,
	q_b_16,
	q_b_113,
	q_b_49,
	q_b_81,
	q_b_17,
	q_b_114,
	q_b_50,
	q_b_82,
	q_b_18,
	q_b_115,
	q_b_51,
	q_b_83,
	q_b_19,
	q_b_116,
	q_b_52,
	q_b_84,
	q_b_20,
	q_b_117,
	q_b_53,
	q_b_85,
	q_b_21,
	q_b_118,
	q_b_54,
	q_b_86,
	q_b_22,
	q_b_119,
	q_b_55,
	q_b_87,
	q_b_23,
	q_b_120,
	q_b_56,
	q_b_88,
	q_b_24,
	q_b_121,
	q_b_57,
	q_b_89,
	q_b_25,
	q_b_122,
	q_b_58,
	q_b_90,
	q_b_26,
	q_b_123,
	q_b_59,
	q_b_91,
	q_b_27,
	q_b_124,
	q_b_60,
	q_b_92,
	q_b_28,
	q_b_125,
	q_b_61,
	q_b_93,
	q_b_29,
	q_b_126,
	q_b_62,
	q_b_94,
	q_b_30,
	q_b_127,
	q_b_63,
	q_b_95,
	q_b_31,
	ready_out,
	int_refresh_ack,
	ctl_init_fail,
	ctl_init_success,
	local_init_done,
	reset_phy_clk_1x_n,
	rdwr_data_valid_r,
	doing_read,
	wd_lat_2,
	wd_lat_1,
	wd_lat_0,
	wd_lat_3,
	wd_lat_4,
	afi_cs_n_1,
	int_cke_r_0,
	afi_addr_0,
	afi_addr_1,
	afi_addr_2,
	afi_addr_3,
	afi_addr_4,
	afi_addr_5,
	afi_addr_6,
	afi_addr_7,
	afi_addr_8,
	afi_addr_9,
	afi_addr_10,
	afi_addr_11,
	afi_addr_12,
	afi_addr_13,
	afi_ba_0,
	afi_ba_1,
	afi_ba_2,
	afi_ras_n_0,
	afi_cas_n_0,
	afi_we_n_0,
	afi_dm_4,
	afi_dm_12,
	afi_dm_0,
	afi_dm_8,
	afi_dm_5,
	afi_dm_13,
	afi_dm_1,
	afi_dm_9,
	afi_dm_6,
	afi_dm_14,
	afi_dm_2,
	afi_dm_10,
	afi_dm_7,
	afi_dm_15,
	afi_dm_3,
	afi_dm_11,
	int_wdata_valid,
	int_dqs_burst,
	int_dqs_burst_hr,
	GND_port,
	local_size_1,
	local_address_0,
	local_size_0,
	local_size_6,
	local_size_5,
	local_size_4,
	local_size_2,
	local_size_3,
	local_read_req,
	local_write_req,
	local_burstbegin,
	local_address_8,
	local_address_10,
	local_address_9,
	local_address_23,
	local_address_24,
	local_address_22,
	local_address_20,
	local_address_21,
	local_address_19,
	local_address_17,
	local_address_18,
	local_address_13,
	local_address_11,
	local_address_12,
	local_address_16,
	local_address_14,
	local_address_15,
	local_address_1,
	local_address_2,
	local_address_3,
	local_address_4,
	local_address_5,
	local_address_7,
	local_address_6,
	local_be_4,
	local_be_12,
	local_be_0,
	local_be_8,
	local_be_5,
	local_be_13,
	local_be_1,
	local_be_9,
	local_be_6,
	local_be_14,
	local_be_2,
	local_be_10,
	local_be_7,
	local_be_15,
	local_be_3,
	local_be_11,
	local_wdata_96,
	local_wdata_32,
	local_wdata_64,
	local_wdata_0,
	local_wdata_97,
	local_wdata_33,
	local_wdata_65,
	local_wdata_1,
	local_wdata_98,
	local_wdata_34,
	local_wdata_66,
	local_wdata_2,
	local_wdata_99,
	local_wdata_35,
	local_wdata_67,
	local_wdata_3,
	local_wdata_100,
	local_wdata_36,
	local_wdata_68,
	local_wdata_4,
	local_wdata_101,
	local_wdata_37,
	local_wdata_69,
	local_wdata_5,
	local_wdata_102,
	local_wdata_38,
	local_wdata_70,
	local_wdata_6,
	local_wdata_103,
	local_wdata_39,
	local_wdata_71,
	local_wdata_7,
	local_wdata_104,
	local_wdata_40,
	local_wdata_72,
	local_wdata_8,
	local_wdata_105,
	local_wdata_41,
	local_wdata_73,
	local_wdata_9,
	local_wdata_106,
	local_wdata_42,
	local_wdata_74,
	local_wdata_10,
	local_wdata_107,
	local_wdata_43,
	local_wdata_75,
	local_wdata_11,
	local_wdata_108,
	local_wdata_44,
	local_wdata_76,
	local_wdata_12,
	local_wdata_109,
	local_wdata_45,
	local_wdata_77,
	local_wdata_13,
	local_wdata_110,
	local_wdata_46,
	local_wdata_78,
	local_wdata_14,
	local_wdata_111,
	local_wdata_47,
	local_wdata_79,
	local_wdata_15,
	local_wdata_112,
	local_wdata_48,
	local_wdata_80,
	local_wdata_16,
	local_wdata_113,
	local_wdata_49,
	local_wdata_81,
	local_wdata_17,
	local_wdata_114,
	local_wdata_50,
	local_wdata_82,
	local_wdata_18,
	local_wdata_115,
	local_wdata_51,
	local_wdata_83,
	local_wdata_19,
	local_wdata_116,
	local_wdata_52,
	local_wdata_84,
	local_wdata_20,
	local_wdata_117,
	local_wdata_53,
	local_wdata_85,
	local_wdata_21,
	local_wdata_118,
	local_wdata_54,
	local_wdata_86,
	local_wdata_22,
	local_wdata_119,
	local_wdata_55,
	local_wdata_87,
	local_wdata_23,
	local_wdata_120,
	local_wdata_56,
	local_wdata_88,
	local_wdata_24,
	local_wdata_121,
	local_wdata_57,
	local_wdata_89,
	local_wdata_25,
	local_wdata_122,
	local_wdata_58,
	local_wdata_90,
	local_wdata_26,
	local_wdata_123,
	local_wdata_59,
	local_wdata_91,
	local_wdata_27,
	local_wdata_124,
	local_wdata_60,
	local_wdata_92,
	local_wdata_28,
	local_wdata_125,
	local_wdata_61,
	local_wdata_93,
	local_wdata_29,
	local_wdata_126,
	local_wdata_62,
	local_wdata_94,
	local_wdata_30,
	local_wdata_127,
	local_wdata_63,
	local_wdata_95,
	local_wdata_31)/* synthesis synthesis_greybox=0 */;
input 	clk_0;
output 	do_read_r;
output 	q_b_96;
output 	q_b_32;
output 	q_b_64;
output 	q_b_0;
output 	q_b_97;
output 	q_b_33;
output 	q_b_65;
output 	q_b_1;
output 	q_b_98;
output 	q_b_34;
output 	q_b_66;
output 	q_b_2;
output 	q_b_99;
output 	q_b_35;
output 	q_b_67;
output 	q_b_3;
output 	q_b_100;
output 	q_b_36;
output 	q_b_68;
output 	q_b_4;
output 	q_b_101;
output 	q_b_37;
output 	q_b_69;
output 	q_b_5;
output 	q_b_102;
output 	q_b_38;
output 	q_b_70;
output 	q_b_6;
output 	q_b_103;
output 	q_b_39;
output 	q_b_71;
output 	q_b_7;
output 	q_b_104;
output 	q_b_40;
output 	q_b_72;
output 	q_b_8;
output 	q_b_105;
output 	q_b_41;
output 	q_b_73;
output 	q_b_9;
output 	q_b_106;
output 	q_b_42;
output 	q_b_74;
output 	q_b_10;
output 	q_b_107;
output 	q_b_43;
output 	q_b_75;
output 	q_b_11;
output 	q_b_108;
output 	q_b_44;
output 	q_b_76;
output 	q_b_12;
output 	q_b_109;
output 	q_b_45;
output 	q_b_77;
output 	q_b_13;
output 	q_b_110;
output 	q_b_46;
output 	q_b_78;
output 	q_b_14;
output 	q_b_111;
output 	q_b_47;
output 	q_b_79;
output 	q_b_15;
output 	q_b_112;
output 	q_b_48;
output 	q_b_80;
output 	q_b_16;
output 	q_b_113;
output 	q_b_49;
output 	q_b_81;
output 	q_b_17;
output 	q_b_114;
output 	q_b_50;
output 	q_b_82;
output 	q_b_18;
output 	q_b_115;
output 	q_b_51;
output 	q_b_83;
output 	q_b_19;
output 	q_b_116;
output 	q_b_52;
output 	q_b_84;
output 	q_b_20;
output 	q_b_117;
output 	q_b_53;
output 	q_b_85;
output 	q_b_21;
output 	q_b_118;
output 	q_b_54;
output 	q_b_86;
output 	q_b_22;
output 	q_b_119;
output 	q_b_55;
output 	q_b_87;
output 	q_b_23;
output 	q_b_120;
output 	q_b_56;
output 	q_b_88;
output 	q_b_24;
output 	q_b_121;
output 	q_b_57;
output 	q_b_89;
output 	q_b_25;
output 	q_b_122;
output 	q_b_58;
output 	q_b_90;
output 	q_b_26;
output 	q_b_123;
output 	q_b_59;
output 	q_b_91;
output 	q_b_27;
output 	q_b_124;
output 	q_b_60;
output 	q_b_92;
output 	q_b_28;
output 	q_b_125;
output 	q_b_61;
output 	q_b_93;
output 	q_b_29;
output 	q_b_126;
output 	q_b_62;
output 	q_b_94;
output 	q_b_30;
output 	q_b_127;
output 	q_b_63;
output 	q_b_95;
output 	q_b_31;
output 	ready_out;
output 	int_refresh_ack;
input 	ctl_init_fail;
input 	ctl_init_success;
output 	local_init_done;
input 	reset_phy_clk_1x_n;
output 	rdwr_data_valid_r;
output 	doing_read;
input 	wd_lat_2;
input 	wd_lat_1;
input 	wd_lat_0;
input 	wd_lat_3;
input 	wd_lat_4;
output 	afi_cs_n_1;
output 	int_cke_r_0;
output 	afi_addr_0;
output 	afi_addr_1;
output 	afi_addr_2;
output 	afi_addr_3;
output 	afi_addr_4;
output 	afi_addr_5;
output 	afi_addr_6;
output 	afi_addr_7;
output 	afi_addr_8;
output 	afi_addr_9;
output 	afi_addr_10;
output 	afi_addr_11;
output 	afi_addr_12;
output 	afi_addr_13;
output 	afi_ba_0;
output 	afi_ba_1;
output 	afi_ba_2;
output 	afi_ras_n_0;
output 	afi_cas_n_0;
output 	afi_we_n_0;
output 	afi_dm_4;
output 	afi_dm_12;
output 	afi_dm_0;
output 	afi_dm_8;
output 	afi_dm_5;
output 	afi_dm_13;
output 	afi_dm_1;
output 	afi_dm_9;
output 	afi_dm_6;
output 	afi_dm_14;
output 	afi_dm_2;
output 	afi_dm_10;
output 	afi_dm_7;
output 	afi_dm_15;
output 	afi_dm_3;
output 	afi_dm_11;
output 	int_wdata_valid;
output 	int_dqs_burst;
output 	int_dqs_burst_hr;
input 	GND_port;
input 	local_size_1;
input 	local_address_0;
input 	local_size_0;
input 	local_size_6;
input 	local_size_5;
input 	local_size_4;
input 	local_size_2;
input 	local_size_3;
input 	local_read_req;
input 	local_write_req;
input 	local_burstbegin;
input 	local_address_8;
input 	local_address_10;
input 	local_address_9;
input 	local_address_23;
input 	local_address_24;
input 	local_address_22;
input 	local_address_20;
input 	local_address_21;
input 	local_address_19;
input 	local_address_17;
input 	local_address_18;
input 	local_address_13;
input 	local_address_11;
input 	local_address_12;
input 	local_address_16;
input 	local_address_14;
input 	local_address_15;
input 	local_address_1;
input 	local_address_2;
input 	local_address_3;
input 	local_address_4;
input 	local_address_5;
input 	local_address_7;
input 	local_address_6;
input 	local_be_4;
input 	local_be_12;
input 	local_be_0;
input 	local_be_8;
input 	local_be_5;
input 	local_be_13;
input 	local_be_1;
input 	local_be_9;
input 	local_be_6;
input 	local_be_14;
input 	local_be_2;
input 	local_be_10;
input 	local_be_7;
input 	local_be_15;
input 	local_be_3;
input 	local_be_11;
input 	local_wdata_96;
input 	local_wdata_32;
input 	local_wdata_64;
input 	local_wdata_0;
input 	local_wdata_97;
input 	local_wdata_33;
input 	local_wdata_65;
input 	local_wdata_1;
input 	local_wdata_98;
input 	local_wdata_34;
input 	local_wdata_66;
input 	local_wdata_2;
input 	local_wdata_99;
input 	local_wdata_35;
input 	local_wdata_67;
input 	local_wdata_3;
input 	local_wdata_100;
input 	local_wdata_36;
input 	local_wdata_68;
input 	local_wdata_4;
input 	local_wdata_101;
input 	local_wdata_37;
input 	local_wdata_69;
input 	local_wdata_5;
input 	local_wdata_102;
input 	local_wdata_38;
input 	local_wdata_70;
input 	local_wdata_6;
input 	local_wdata_103;
input 	local_wdata_39;
input 	local_wdata_71;
input 	local_wdata_7;
input 	local_wdata_104;
input 	local_wdata_40;
input 	local_wdata_72;
input 	local_wdata_8;
input 	local_wdata_105;
input 	local_wdata_41;
input 	local_wdata_73;
input 	local_wdata_9;
input 	local_wdata_106;
input 	local_wdata_42;
input 	local_wdata_74;
input 	local_wdata_10;
input 	local_wdata_107;
input 	local_wdata_43;
input 	local_wdata_75;
input 	local_wdata_11;
input 	local_wdata_108;
input 	local_wdata_44;
input 	local_wdata_76;
input 	local_wdata_12;
input 	local_wdata_109;
input 	local_wdata_45;
input 	local_wdata_77;
input 	local_wdata_13;
input 	local_wdata_110;
input 	local_wdata_46;
input 	local_wdata_78;
input 	local_wdata_14;
input 	local_wdata_111;
input 	local_wdata_47;
input 	local_wdata_79;
input 	local_wdata_15;
input 	local_wdata_112;
input 	local_wdata_48;
input 	local_wdata_80;
input 	local_wdata_16;
input 	local_wdata_113;
input 	local_wdata_49;
input 	local_wdata_81;
input 	local_wdata_17;
input 	local_wdata_114;
input 	local_wdata_50;
input 	local_wdata_82;
input 	local_wdata_18;
input 	local_wdata_115;
input 	local_wdata_51;
input 	local_wdata_83;
input 	local_wdata_19;
input 	local_wdata_116;
input 	local_wdata_52;
input 	local_wdata_84;
input 	local_wdata_20;
input 	local_wdata_117;
input 	local_wdata_53;
input 	local_wdata_85;
input 	local_wdata_21;
input 	local_wdata_118;
input 	local_wdata_54;
input 	local_wdata_86;
input 	local_wdata_22;
input 	local_wdata_119;
input 	local_wdata_55;
input 	local_wdata_87;
input 	local_wdata_23;
input 	local_wdata_120;
input 	local_wdata_56;
input 	local_wdata_88;
input 	local_wdata_24;
input 	local_wdata_121;
input 	local_wdata_57;
input 	local_wdata_89;
input 	local_wdata_25;
input 	local_wdata_122;
input 	local_wdata_58;
input 	local_wdata_90;
input 	local_wdata_26;
input 	local_wdata_123;
input 	local_wdata_59;
input 	local_wdata_91;
input 	local_wdata_27;
input 	local_wdata_124;
input 	local_wdata_60;
input 	local_wdata_92;
input 	local_wdata_28;
input 	local_wdata_125;
input 	local_wdata_61;
input 	local_wdata_93;
input 	local_wdata_29;
input 	local_wdata_126;
input 	local_wdata_62;
input 	local_wdata_94;
input 	local_wdata_30;
input 	local_wdata_127;
input 	local_wdata_63;
input 	local_wdata_95;
input 	local_wdata_31;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_alt_ddrx_controller alt_ddrx_controller_inst(
	.clk_0(clk_0),
	.do_read_r(do_read_r),
	.q_b_96(q_b_96),
	.q_b_32(q_b_32),
	.q_b_64(q_b_64),
	.q_b_0(q_b_0),
	.q_b_97(q_b_97),
	.q_b_33(q_b_33),
	.q_b_65(q_b_65),
	.q_b_1(q_b_1),
	.q_b_98(q_b_98),
	.q_b_34(q_b_34),
	.q_b_66(q_b_66),
	.q_b_2(q_b_2),
	.q_b_99(q_b_99),
	.q_b_35(q_b_35),
	.q_b_67(q_b_67),
	.q_b_3(q_b_3),
	.q_b_100(q_b_100),
	.q_b_36(q_b_36),
	.q_b_68(q_b_68),
	.q_b_4(q_b_4),
	.q_b_101(q_b_101),
	.q_b_37(q_b_37),
	.q_b_69(q_b_69),
	.q_b_5(q_b_5),
	.q_b_102(q_b_102),
	.q_b_38(q_b_38),
	.q_b_70(q_b_70),
	.q_b_6(q_b_6),
	.q_b_103(q_b_103),
	.q_b_39(q_b_39),
	.q_b_71(q_b_71),
	.q_b_7(q_b_7),
	.q_b_104(q_b_104),
	.q_b_40(q_b_40),
	.q_b_72(q_b_72),
	.q_b_8(q_b_8),
	.q_b_105(q_b_105),
	.q_b_41(q_b_41),
	.q_b_73(q_b_73),
	.q_b_9(q_b_9),
	.q_b_106(q_b_106),
	.q_b_42(q_b_42),
	.q_b_74(q_b_74),
	.q_b_10(q_b_10),
	.q_b_107(q_b_107),
	.q_b_43(q_b_43),
	.q_b_75(q_b_75),
	.q_b_11(q_b_11),
	.q_b_108(q_b_108),
	.q_b_44(q_b_44),
	.q_b_76(q_b_76),
	.q_b_12(q_b_12),
	.q_b_109(q_b_109),
	.q_b_45(q_b_45),
	.q_b_77(q_b_77),
	.q_b_13(q_b_13),
	.q_b_110(q_b_110),
	.q_b_46(q_b_46),
	.q_b_78(q_b_78),
	.q_b_14(q_b_14),
	.q_b_111(q_b_111),
	.q_b_47(q_b_47),
	.q_b_79(q_b_79),
	.q_b_15(q_b_15),
	.q_b_112(q_b_112),
	.q_b_48(q_b_48),
	.q_b_80(q_b_80),
	.q_b_16(q_b_16),
	.q_b_113(q_b_113),
	.q_b_49(q_b_49),
	.q_b_81(q_b_81),
	.q_b_17(q_b_17),
	.q_b_114(q_b_114),
	.q_b_50(q_b_50),
	.q_b_82(q_b_82),
	.q_b_18(q_b_18),
	.q_b_115(q_b_115),
	.q_b_51(q_b_51),
	.q_b_83(q_b_83),
	.q_b_19(q_b_19),
	.q_b_116(q_b_116),
	.q_b_52(q_b_52),
	.q_b_84(q_b_84),
	.q_b_20(q_b_20),
	.q_b_117(q_b_117),
	.q_b_53(q_b_53),
	.q_b_85(q_b_85),
	.q_b_21(q_b_21),
	.q_b_118(q_b_118),
	.q_b_54(q_b_54),
	.q_b_86(q_b_86),
	.q_b_22(q_b_22),
	.q_b_119(q_b_119),
	.q_b_55(q_b_55),
	.q_b_87(q_b_87),
	.q_b_23(q_b_23),
	.q_b_120(q_b_120),
	.q_b_56(q_b_56),
	.q_b_88(q_b_88),
	.q_b_24(q_b_24),
	.q_b_121(q_b_121),
	.q_b_57(q_b_57),
	.q_b_89(q_b_89),
	.q_b_25(q_b_25),
	.q_b_122(q_b_122),
	.q_b_58(q_b_58),
	.q_b_90(q_b_90),
	.q_b_26(q_b_26),
	.q_b_123(q_b_123),
	.q_b_59(q_b_59),
	.q_b_91(q_b_91),
	.q_b_27(q_b_27),
	.q_b_124(q_b_124),
	.q_b_60(q_b_60),
	.q_b_92(q_b_92),
	.q_b_28(q_b_28),
	.q_b_125(q_b_125),
	.q_b_61(q_b_61),
	.q_b_93(q_b_93),
	.q_b_29(q_b_29),
	.q_b_126(q_b_126),
	.q_b_62(q_b_62),
	.q_b_94(q_b_94),
	.q_b_30(q_b_30),
	.q_b_127(q_b_127),
	.q_b_63(q_b_63),
	.q_b_95(q_b_95),
	.q_b_31(q_b_31),
	.ready_out(ready_out),
	.int_refresh_ack(int_refresh_ack),
	.ctl_init_fail(ctl_init_fail),
	.ctl_init_success(ctl_init_success),
	.local_init_done(local_init_done),
	.reset_phy_clk_1x_n(reset_phy_clk_1x_n),
	.rdwr_data_valid_r(rdwr_data_valid_r),
	.doing_read(doing_read),
	.wd_lat_2(wd_lat_2),
	.wd_lat_1(wd_lat_1),
	.wd_lat_0(wd_lat_0),
	.wd_lat_3(wd_lat_3),
	.wd_lat_4(wd_lat_4),
	.afi_cs_n_1(afi_cs_n_1),
	.int_cke_r_0(int_cke_r_0),
	.afi_addr_0(afi_addr_0),
	.afi_addr_1(afi_addr_1),
	.afi_addr_2(afi_addr_2),
	.afi_addr_3(afi_addr_3),
	.afi_addr_4(afi_addr_4),
	.afi_addr_5(afi_addr_5),
	.afi_addr_6(afi_addr_6),
	.afi_addr_7(afi_addr_7),
	.afi_addr_8(afi_addr_8),
	.afi_addr_9(afi_addr_9),
	.afi_addr_10(afi_addr_10),
	.afi_addr_11(afi_addr_11),
	.afi_addr_12(afi_addr_12),
	.afi_addr_13(afi_addr_13),
	.afi_ba_0(afi_ba_0),
	.afi_ba_1(afi_ba_1),
	.afi_ba_2(afi_ba_2),
	.afi_ras_n_0(afi_ras_n_0),
	.afi_cas_n_0(afi_cas_n_0),
	.afi_we_n_0(afi_we_n_0),
	.afi_dm_4(afi_dm_4),
	.afi_dm_12(afi_dm_12),
	.afi_dm_0(afi_dm_0),
	.afi_dm_8(afi_dm_8),
	.afi_dm_5(afi_dm_5),
	.afi_dm_13(afi_dm_13),
	.afi_dm_1(afi_dm_1),
	.afi_dm_9(afi_dm_9),
	.afi_dm_6(afi_dm_6),
	.afi_dm_14(afi_dm_14),
	.afi_dm_2(afi_dm_2),
	.afi_dm_10(afi_dm_10),
	.afi_dm_7(afi_dm_7),
	.afi_dm_15(afi_dm_15),
	.afi_dm_3(afi_dm_3),
	.afi_dm_11(afi_dm_11),
	.int_wdata_valid(int_wdata_valid),
	.int_dqs_burst(int_dqs_burst),
	.int_dqs_burst_hr(int_dqs_burst_hr),
	.GND_port(GND_port),
	.local_size_1(local_size_1),
	.local_address_0(local_address_0),
	.local_size_0(local_size_0),
	.local_size_6(local_size_6),
	.local_size_5(local_size_5),
	.local_size_4(local_size_4),
	.local_size_2(local_size_2),
	.local_size_3(local_size_3),
	.local_read_req(local_read_req),
	.local_write_req(local_write_req),
	.local_burstbegin(local_burstbegin),
	.local_address_8(local_address_8),
	.local_address_10(local_address_10),
	.local_address_9(local_address_9),
	.local_address_23(local_address_23),
	.local_address_24(local_address_24),
	.local_address_22(local_address_22),
	.local_address_20(local_address_20),
	.local_address_21(local_address_21),
	.local_address_19(local_address_19),
	.local_address_17(local_address_17),
	.local_address_18(local_address_18),
	.local_address_13(local_address_13),
	.local_address_11(local_address_11),
	.local_address_12(local_address_12),
	.local_address_16(local_address_16),
	.local_address_14(local_address_14),
	.local_address_15(local_address_15),
	.local_address_1(local_address_1),
	.local_address_2(local_address_2),
	.local_address_3(local_address_3),
	.local_address_4(local_address_4),
	.local_address_5(local_address_5),
	.local_address_7(local_address_7),
	.local_address_6(local_address_6),
	.local_be_4(local_be_4),
	.local_be_12(local_be_12),
	.local_be_0(local_be_0),
	.local_be_8(local_be_8),
	.local_be_5(local_be_5),
	.local_be_13(local_be_13),
	.local_be_1(local_be_1),
	.local_be_9(local_be_9),
	.local_be_6(local_be_6),
	.local_be_14(local_be_14),
	.local_be_2(local_be_2),
	.local_be_10(local_be_10),
	.local_be_7(local_be_7),
	.local_be_15(local_be_15),
	.local_be_3(local_be_3),
	.local_be_11(local_be_11),
	.local_wdata_96(local_wdata_96),
	.local_wdata_32(local_wdata_32),
	.local_wdata_64(local_wdata_64),
	.local_wdata_0(local_wdata_0),
	.local_wdata_97(local_wdata_97),
	.local_wdata_33(local_wdata_33),
	.local_wdata_65(local_wdata_65),
	.local_wdata_1(local_wdata_1),
	.local_wdata_98(local_wdata_98),
	.local_wdata_34(local_wdata_34),
	.local_wdata_66(local_wdata_66),
	.local_wdata_2(local_wdata_2),
	.local_wdata_99(local_wdata_99),
	.local_wdata_35(local_wdata_35),
	.local_wdata_67(local_wdata_67),
	.local_wdata_3(local_wdata_3),
	.local_wdata_100(local_wdata_100),
	.local_wdata_36(local_wdata_36),
	.local_wdata_68(local_wdata_68),
	.local_wdata_4(local_wdata_4),
	.local_wdata_101(local_wdata_101),
	.local_wdata_37(local_wdata_37),
	.local_wdata_69(local_wdata_69),
	.local_wdata_5(local_wdata_5),
	.local_wdata_102(local_wdata_102),
	.local_wdata_38(local_wdata_38),
	.local_wdata_70(local_wdata_70),
	.local_wdata_6(local_wdata_6),
	.local_wdata_103(local_wdata_103),
	.local_wdata_39(local_wdata_39),
	.local_wdata_71(local_wdata_71),
	.local_wdata_7(local_wdata_7),
	.local_wdata_104(local_wdata_104),
	.local_wdata_40(local_wdata_40),
	.local_wdata_72(local_wdata_72),
	.local_wdata_8(local_wdata_8),
	.local_wdata_105(local_wdata_105),
	.local_wdata_41(local_wdata_41),
	.local_wdata_73(local_wdata_73),
	.local_wdata_9(local_wdata_9),
	.local_wdata_106(local_wdata_106),
	.local_wdata_42(local_wdata_42),
	.local_wdata_74(local_wdata_74),
	.local_wdata_10(local_wdata_10),
	.local_wdata_107(local_wdata_107),
	.local_wdata_43(local_wdata_43),
	.local_wdata_75(local_wdata_75),
	.local_wdata_11(local_wdata_11),
	.local_wdata_108(local_wdata_108),
	.local_wdata_44(local_wdata_44),
	.local_wdata_76(local_wdata_76),
	.local_wdata_12(local_wdata_12),
	.local_wdata_109(local_wdata_109),
	.local_wdata_45(local_wdata_45),
	.local_wdata_77(local_wdata_77),
	.local_wdata_13(local_wdata_13),
	.local_wdata_110(local_wdata_110),
	.local_wdata_46(local_wdata_46),
	.local_wdata_78(local_wdata_78),
	.local_wdata_14(local_wdata_14),
	.local_wdata_111(local_wdata_111),
	.local_wdata_47(local_wdata_47),
	.local_wdata_79(local_wdata_79),
	.local_wdata_15(local_wdata_15),
	.local_wdata_112(local_wdata_112),
	.local_wdata_48(local_wdata_48),
	.local_wdata_80(local_wdata_80),
	.local_wdata_16(local_wdata_16),
	.local_wdata_113(local_wdata_113),
	.local_wdata_49(local_wdata_49),
	.local_wdata_81(local_wdata_81),
	.local_wdata_17(local_wdata_17),
	.local_wdata_114(local_wdata_114),
	.local_wdata_50(local_wdata_50),
	.local_wdata_82(local_wdata_82),
	.local_wdata_18(local_wdata_18),
	.local_wdata_115(local_wdata_115),
	.local_wdata_51(local_wdata_51),
	.local_wdata_83(local_wdata_83),
	.local_wdata_19(local_wdata_19),
	.local_wdata_116(local_wdata_116),
	.local_wdata_52(local_wdata_52),
	.local_wdata_84(local_wdata_84),
	.local_wdata_20(local_wdata_20),
	.local_wdata_117(local_wdata_117),
	.local_wdata_53(local_wdata_53),
	.local_wdata_85(local_wdata_85),
	.local_wdata_21(local_wdata_21),
	.local_wdata_118(local_wdata_118),
	.local_wdata_54(local_wdata_54),
	.local_wdata_86(local_wdata_86),
	.local_wdata_22(local_wdata_22),
	.local_wdata_119(local_wdata_119),
	.local_wdata_55(local_wdata_55),
	.local_wdata_87(local_wdata_87),
	.local_wdata_23(local_wdata_23),
	.local_wdata_120(local_wdata_120),
	.local_wdata_56(local_wdata_56),
	.local_wdata_88(local_wdata_88),
	.local_wdata_24(local_wdata_24),
	.local_wdata_121(local_wdata_121),
	.local_wdata_57(local_wdata_57),
	.local_wdata_89(local_wdata_89),
	.local_wdata_25(local_wdata_25),
	.local_wdata_122(local_wdata_122),
	.local_wdata_58(local_wdata_58),
	.local_wdata_90(local_wdata_90),
	.local_wdata_26(local_wdata_26),
	.local_wdata_123(local_wdata_123),
	.local_wdata_59(local_wdata_59),
	.local_wdata_91(local_wdata_91),
	.local_wdata_27(local_wdata_27),
	.local_wdata_124(local_wdata_124),
	.local_wdata_60(local_wdata_60),
	.local_wdata_92(local_wdata_92),
	.local_wdata_28(local_wdata_28),
	.local_wdata_125(local_wdata_125),
	.local_wdata_61(local_wdata_61),
	.local_wdata_93(local_wdata_93),
	.local_wdata_29(local_wdata_29),
	.local_wdata_126(local_wdata_126),
	.local_wdata_62(local_wdata_62),
	.local_wdata_94(local_wdata_94),
	.local_wdata_30(local_wdata_30),
	.local_wdata_127(local_wdata_127),
	.local_wdata_63(local_wdata_63),
	.local_wdata_95(local_wdata_95),
	.local_wdata_31(local_wdata_31));

endmodule

module ddr3_int_alt_ddrx_controller (
	clk_0,
	do_read_r,
	q_b_96,
	q_b_32,
	q_b_64,
	q_b_0,
	q_b_97,
	q_b_33,
	q_b_65,
	q_b_1,
	q_b_98,
	q_b_34,
	q_b_66,
	q_b_2,
	q_b_99,
	q_b_35,
	q_b_67,
	q_b_3,
	q_b_100,
	q_b_36,
	q_b_68,
	q_b_4,
	q_b_101,
	q_b_37,
	q_b_69,
	q_b_5,
	q_b_102,
	q_b_38,
	q_b_70,
	q_b_6,
	q_b_103,
	q_b_39,
	q_b_71,
	q_b_7,
	q_b_104,
	q_b_40,
	q_b_72,
	q_b_8,
	q_b_105,
	q_b_41,
	q_b_73,
	q_b_9,
	q_b_106,
	q_b_42,
	q_b_74,
	q_b_10,
	q_b_107,
	q_b_43,
	q_b_75,
	q_b_11,
	q_b_108,
	q_b_44,
	q_b_76,
	q_b_12,
	q_b_109,
	q_b_45,
	q_b_77,
	q_b_13,
	q_b_110,
	q_b_46,
	q_b_78,
	q_b_14,
	q_b_111,
	q_b_47,
	q_b_79,
	q_b_15,
	q_b_112,
	q_b_48,
	q_b_80,
	q_b_16,
	q_b_113,
	q_b_49,
	q_b_81,
	q_b_17,
	q_b_114,
	q_b_50,
	q_b_82,
	q_b_18,
	q_b_115,
	q_b_51,
	q_b_83,
	q_b_19,
	q_b_116,
	q_b_52,
	q_b_84,
	q_b_20,
	q_b_117,
	q_b_53,
	q_b_85,
	q_b_21,
	q_b_118,
	q_b_54,
	q_b_86,
	q_b_22,
	q_b_119,
	q_b_55,
	q_b_87,
	q_b_23,
	q_b_120,
	q_b_56,
	q_b_88,
	q_b_24,
	q_b_121,
	q_b_57,
	q_b_89,
	q_b_25,
	q_b_122,
	q_b_58,
	q_b_90,
	q_b_26,
	q_b_123,
	q_b_59,
	q_b_91,
	q_b_27,
	q_b_124,
	q_b_60,
	q_b_92,
	q_b_28,
	q_b_125,
	q_b_61,
	q_b_93,
	q_b_29,
	q_b_126,
	q_b_62,
	q_b_94,
	q_b_30,
	q_b_127,
	q_b_63,
	q_b_95,
	q_b_31,
	ready_out,
	int_refresh_ack,
	ctl_init_fail,
	ctl_init_success,
	local_init_done,
	reset_phy_clk_1x_n,
	rdwr_data_valid_r,
	doing_read,
	wd_lat_2,
	wd_lat_1,
	wd_lat_0,
	wd_lat_3,
	wd_lat_4,
	afi_cs_n_1,
	int_cke_r_0,
	afi_addr_0,
	afi_addr_1,
	afi_addr_2,
	afi_addr_3,
	afi_addr_4,
	afi_addr_5,
	afi_addr_6,
	afi_addr_7,
	afi_addr_8,
	afi_addr_9,
	afi_addr_10,
	afi_addr_11,
	afi_addr_12,
	afi_addr_13,
	afi_ba_0,
	afi_ba_1,
	afi_ba_2,
	afi_ras_n_0,
	afi_cas_n_0,
	afi_we_n_0,
	afi_dm_4,
	afi_dm_12,
	afi_dm_0,
	afi_dm_8,
	afi_dm_5,
	afi_dm_13,
	afi_dm_1,
	afi_dm_9,
	afi_dm_6,
	afi_dm_14,
	afi_dm_2,
	afi_dm_10,
	afi_dm_7,
	afi_dm_15,
	afi_dm_3,
	afi_dm_11,
	int_wdata_valid,
	int_dqs_burst,
	int_dqs_burst_hr,
	GND_port,
	local_size_1,
	local_address_0,
	local_size_0,
	local_size_6,
	local_size_5,
	local_size_4,
	local_size_2,
	local_size_3,
	local_read_req,
	local_write_req,
	local_burstbegin,
	local_address_8,
	local_address_10,
	local_address_9,
	local_address_23,
	local_address_24,
	local_address_22,
	local_address_20,
	local_address_21,
	local_address_19,
	local_address_17,
	local_address_18,
	local_address_13,
	local_address_11,
	local_address_12,
	local_address_16,
	local_address_14,
	local_address_15,
	local_address_1,
	local_address_2,
	local_address_3,
	local_address_4,
	local_address_5,
	local_address_7,
	local_address_6,
	local_be_4,
	local_be_12,
	local_be_0,
	local_be_8,
	local_be_5,
	local_be_13,
	local_be_1,
	local_be_9,
	local_be_6,
	local_be_14,
	local_be_2,
	local_be_10,
	local_be_7,
	local_be_15,
	local_be_3,
	local_be_11,
	local_wdata_96,
	local_wdata_32,
	local_wdata_64,
	local_wdata_0,
	local_wdata_97,
	local_wdata_33,
	local_wdata_65,
	local_wdata_1,
	local_wdata_98,
	local_wdata_34,
	local_wdata_66,
	local_wdata_2,
	local_wdata_99,
	local_wdata_35,
	local_wdata_67,
	local_wdata_3,
	local_wdata_100,
	local_wdata_36,
	local_wdata_68,
	local_wdata_4,
	local_wdata_101,
	local_wdata_37,
	local_wdata_69,
	local_wdata_5,
	local_wdata_102,
	local_wdata_38,
	local_wdata_70,
	local_wdata_6,
	local_wdata_103,
	local_wdata_39,
	local_wdata_71,
	local_wdata_7,
	local_wdata_104,
	local_wdata_40,
	local_wdata_72,
	local_wdata_8,
	local_wdata_105,
	local_wdata_41,
	local_wdata_73,
	local_wdata_9,
	local_wdata_106,
	local_wdata_42,
	local_wdata_74,
	local_wdata_10,
	local_wdata_107,
	local_wdata_43,
	local_wdata_75,
	local_wdata_11,
	local_wdata_108,
	local_wdata_44,
	local_wdata_76,
	local_wdata_12,
	local_wdata_109,
	local_wdata_45,
	local_wdata_77,
	local_wdata_13,
	local_wdata_110,
	local_wdata_46,
	local_wdata_78,
	local_wdata_14,
	local_wdata_111,
	local_wdata_47,
	local_wdata_79,
	local_wdata_15,
	local_wdata_112,
	local_wdata_48,
	local_wdata_80,
	local_wdata_16,
	local_wdata_113,
	local_wdata_49,
	local_wdata_81,
	local_wdata_17,
	local_wdata_114,
	local_wdata_50,
	local_wdata_82,
	local_wdata_18,
	local_wdata_115,
	local_wdata_51,
	local_wdata_83,
	local_wdata_19,
	local_wdata_116,
	local_wdata_52,
	local_wdata_84,
	local_wdata_20,
	local_wdata_117,
	local_wdata_53,
	local_wdata_85,
	local_wdata_21,
	local_wdata_118,
	local_wdata_54,
	local_wdata_86,
	local_wdata_22,
	local_wdata_119,
	local_wdata_55,
	local_wdata_87,
	local_wdata_23,
	local_wdata_120,
	local_wdata_56,
	local_wdata_88,
	local_wdata_24,
	local_wdata_121,
	local_wdata_57,
	local_wdata_89,
	local_wdata_25,
	local_wdata_122,
	local_wdata_58,
	local_wdata_90,
	local_wdata_26,
	local_wdata_123,
	local_wdata_59,
	local_wdata_91,
	local_wdata_27,
	local_wdata_124,
	local_wdata_60,
	local_wdata_92,
	local_wdata_28,
	local_wdata_125,
	local_wdata_61,
	local_wdata_93,
	local_wdata_29,
	local_wdata_126,
	local_wdata_62,
	local_wdata_94,
	local_wdata_30,
	local_wdata_127,
	local_wdata_63,
	local_wdata_95,
	local_wdata_31)/* synthesis synthesis_greybox=0 */;
input 	clk_0;
output 	do_read_r;
output 	q_b_96;
output 	q_b_32;
output 	q_b_64;
output 	q_b_0;
output 	q_b_97;
output 	q_b_33;
output 	q_b_65;
output 	q_b_1;
output 	q_b_98;
output 	q_b_34;
output 	q_b_66;
output 	q_b_2;
output 	q_b_99;
output 	q_b_35;
output 	q_b_67;
output 	q_b_3;
output 	q_b_100;
output 	q_b_36;
output 	q_b_68;
output 	q_b_4;
output 	q_b_101;
output 	q_b_37;
output 	q_b_69;
output 	q_b_5;
output 	q_b_102;
output 	q_b_38;
output 	q_b_70;
output 	q_b_6;
output 	q_b_103;
output 	q_b_39;
output 	q_b_71;
output 	q_b_7;
output 	q_b_104;
output 	q_b_40;
output 	q_b_72;
output 	q_b_8;
output 	q_b_105;
output 	q_b_41;
output 	q_b_73;
output 	q_b_9;
output 	q_b_106;
output 	q_b_42;
output 	q_b_74;
output 	q_b_10;
output 	q_b_107;
output 	q_b_43;
output 	q_b_75;
output 	q_b_11;
output 	q_b_108;
output 	q_b_44;
output 	q_b_76;
output 	q_b_12;
output 	q_b_109;
output 	q_b_45;
output 	q_b_77;
output 	q_b_13;
output 	q_b_110;
output 	q_b_46;
output 	q_b_78;
output 	q_b_14;
output 	q_b_111;
output 	q_b_47;
output 	q_b_79;
output 	q_b_15;
output 	q_b_112;
output 	q_b_48;
output 	q_b_80;
output 	q_b_16;
output 	q_b_113;
output 	q_b_49;
output 	q_b_81;
output 	q_b_17;
output 	q_b_114;
output 	q_b_50;
output 	q_b_82;
output 	q_b_18;
output 	q_b_115;
output 	q_b_51;
output 	q_b_83;
output 	q_b_19;
output 	q_b_116;
output 	q_b_52;
output 	q_b_84;
output 	q_b_20;
output 	q_b_117;
output 	q_b_53;
output 	q_b_85;
output 	q_b_21;
output 	q_b_118;
output 	q_b_54;
output 	q_b_86;
output 	q_b_22;
output 	q_b_119;
output 	q_b_55;
output 	q_b_87;
output 	q_b_23;
output 	q_b_120;
output 	q_b_56;
output 	q_b_88;
output 	q_b_24;
output 	q_b_121;
output 	q_b_57;
output 	q_b_89;
output 	q_b_25;
output 	q_b_122;
output 	q_b_58;
output 	q_b_90;
output 	q_b_26;
output 	q_b_123;
output 	q_b_59;
output 	q_b_91;
output 	q_b_27;
output 	q_b_124;
output 	q_b_60;
output 	q_b_92;
output 	q_b_28;
output 	q_b_125;
output 	q_b_61;
output 	q_b_93;
output 	q_b_29;
output 	q_b_126;
output 	q_b_62;
output 	q_b_94;
output 	q_b_30;
output 	q_b_127;
output 	q_b_63;
output 	q_b_95;
output 	q_b_31;
output 	ready_out;
output 	int_refresh_ack;
input 	ctl_init_fail;
input 	ctl_init_success;
output 	local_init_done;
input 	reset_phy_clk_1x_n;
output 	rdwr_data_valid_r;
output 	doing_read;
input 	wd_lat_2;
input 	wd_lat_1;
input 	wd_lat_0;
input 	wd_lat_3;
input 	wd_lat_4;
output 	afi_cs_n_1;
output 	int_cke_r_0;
output 	afi_addr_0;
output 	afi_addr_1;
output 	afi_addr_2;
output 	afi_addr_3;
output 	afi_addr_4;
output 	afi_addr_5;
output 	afi_addr_6;
output 	afi_addr_7;
output 	afi_addr_8;
output 	afi_addr_9;
output 	afi_addr_10;
output 	afi_addr_11;
output 	afi_addr_12;
output 	afi_addr_13;
output 	afi_ba_0;
output 	afi_ba_1;
output 	afi_ba_2;
output 	afi_ras_n_0;
output 	afi_cas_n_0;
output 	afi_we_n_0;
output 	afi_dm_4;
output 	afi_dm_12;
output 	afi_dm_0;
output 	afi_dm_8;
output 	afi_dm_5;
output 	afi_dm_13;
output 	afi_dm_1;
output 	afi_dm_9;
output 	afi_dm_6;
output 	afi_dm_14;
output 	afi_dm_2;
output 	afi_dm_10;
output 	afi_dm_7;
output 	afi_dm_15;
output 	afi_dm_3;
output 	afi_dm_11;
output 	int_wdata_valid;
output 	int_dqs_burst;
output 	int_dqs_burst_hr;
input 	GND_port;
input 	local_size_1;
input 	local_address_0;
input 	local_size_0;
input 	local_size_6;
input 	local_size_5;
input 	local_size_4;
input 	local_size_2;
input 	local_size_3;
input 	local_read_req;
input 	local_write_req;
input 	local_burstbegin;
input 	local_address_8;
input 	local_address_10;
input 	local_address_9;
input 	local_address_23;
input 	local_address_24;
input 	local_address_22;
input 	local_address_20;
input 	local_address_21;
input 	local_address_19;
input 	local_address_17;
input 	local_address_18;
input 	local_address_13;
input 	local_address_11;
input 	local_address_12;
input 	local_address_16;
input 	local_address_14;
input 	local_address_15;
input 	local_address_1;
input 	local_address_2;
input 	local_address_3;
input 	local_address_4;
input 	local_address_5;
input 	local_address_7;
input 	local_address_6;
input 	local_be_4;
input 	local_be_12;
input 	local_be_0;
input 	local_be_8;
input 	local_be_5;
input 	local_be_13;
input 	local_be_1;
input 	local_be_9;
input 	local_be_6;
input 	local_be_14;
input 	local_be_2;
input 	local_be_10;
input 	local_be_7;
input 	local_be_15;
input 	local_be_3;
input 	local_be_11;
input 	local_wdata_96;
input 	local_wdata_32;
input 	local_wdata_64;
input 	local_wdata_0;
input 	local_wdata_97;
input 	local_wdata_33;
input 	local_wdata_65;
input 	local_wdata_1;
input 	local_wdata_98;
input 	local_wdata_34;
input 	local_wdata_66;
input 	local_wdata_2;
input 	local_wdata_99;
input 	local_wdata_35;
input 	local_wdata_67;
input 	local_wdata_3;
input 	local_wdata_100;
input 	local_wdata_36;
input 	local_wdata_68;
input 	local_wdata_4;
input 	local_wdata_101;
input 	local_wdata_37;
input 	local_wdata_69;
input 	local_wdata_5;
input 	local_wdata_102;
input 	local_wdata_38;
input 	local_wdata_70;
input 	local_wdata_6;
input 	local_wdata_103;
input 	local_wdata_39;
input 	local_wdata_71;
input 	local_wdata_7;
input 	local_wdata_104;
input 	local_wdata_40;
input 	local_wdata_72;
input 	local_wdata_8;
input 	local_wdata_105;
input 	local_wdata_41;
input 	local_wdata_73;
input 	local_wdata_9;
input 	local_wdata_106;
input 	local_wdata_42;
input 	local_wdata_74;
input 	local_wdata_10;
input 	local_wdata_107;
input 	local_wdata_43;
input 	local_wdata_75;
input 	local_wdata_11;
input 	local_wdata_108;
input 	local_wdata_44;
input 	local_wdata_76;
input 	local_wdata_12;
input 	local_wdata_109;
input 	local_wdata_45;
input 	local_wdata_77;
input 	local_wdata_13;
input 	local_wdata_110;
input 	local_wdata_46;
input 	local_wdata_78;
input 	local_wdata_14;
input 	local_wdata_111;
input 	local_wdata_47;
input 	local_wdata_79;
input 	local_wdata_15;
input 	local_wdata_112;
input 	local_wdata_48;
input 	local_wdata_80;
input 	local_wdata_16;
input 	local_wdata_113;
input 	local_wdata_49;
input 	local_wdata_81;
input 	local_wdata_17;
input 	local_wdata_114;
input 	local_wdata_50;
input 	local_wdata_82;
input 	local_wdata_18;
input 	local_wdata_115;
input 	local_wdata_51;
input 	local_wdata_83;
input 	local_wdata_19;
input 	local_wdata_116;
input 	local_wdata_52;
input 	local_wdata_84;
input 	local_wdata_20;
input 	local_wdata_117;
input 	local_wdata_53;
input 	local_wdata_85;
input 	local_wdata_21;
input 	local_wdata_118;
input 	local_wdata_54;
input 	local_wdata_86;
input 	local_wdata_22;
input 	local_wdata_119;
input 	local_wdata_55;
input 	local_wdata_87;
input 	local_wdata_23;
input 	local_wdata_120;
input 	local_wdata_56;
input 	local_wdata_88;
input 	local_wdata_24;
input 	local_wdata_121;
input 	local_wdata_57;
input 	local_wdata_89;
input 	local_wdata_25;
input 	local_wdata_122;
input 	local_wdata_58;
input 	local_wdata_90;
input 	local_wdata_26;
input 	local_wdata_123;
input 	local_wdata_59;
input 	local_wdata_91;
input 	local_wdata_27;
input 	local_wdata_124;
input 	local_wdata_60;
input 	local_wdata_92;
input 	local_wdata_28;
input 	local_wdata_125;
input 	local_wdata_61;
input 	local_wdata_93;
input 	local_wdata_29;
input 	local_wdata_126;
input 	local_wdata_62;
input 	local_wdata_94;
input 	local_wdata_30;
input 	local_wdata_127;
input 	local_wdata_63;
input 	local_wdata_95;
input 	local_wdata_31;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \bank_timer_wrapper_inst|rank_monitor_inst|auto_refresh_logic_per_chip[0].int_refresh_req~q ;
wire \bank_timer_wrapper_inst|bypass_inst|out_cmd_info_valid[0]~q ;
wire \state_machine_inst|do_auto_precharge_r~q ;
wire \state_machine_inst|do_write_r~q ;
wire \bank_timer_wrapper_inst|bypass_inst|out_cmd_info_valid[2]~q ;
wire \bank_timer_wrapper_inst|bypass_inst|out_cmd_info_valid[3]~q ;
wire \bank_timer_wrapper_inst|bypass_inst|out_cmd_info_valid[4]~q ;
wire \bank_timer_wrapper_inst|bypass_inst|out_cmd_info_valid[1]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[0][10]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[0][12]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[0][11]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[0][32]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[2][12]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[3][12]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[1][12]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[2][10]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[3][10]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[1][10]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[2][11]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[3][11]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[1][11]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[0][29]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[0][28]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[0][33]~q ;
wire \state_machine_inst|do_burst_chop_r~q ;
wire \input_if_inst|cmd_queue_inst|pipe[4][12]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[4][11]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[4][10]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[5][25]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[0][25]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[5][26]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[0][26]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[5][24]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[0][24]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[5][22]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[0][22]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[5][23]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[0][23]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[5][21]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[0][21]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[5][19]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[0][19]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[5][20]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[0][20]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[5][15]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[0][15]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[5][13]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[0][13]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[5][14]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[0][14]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[5][18]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[0][18]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[5][16]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[0][16]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[5][17]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[0][17]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[5][12]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[5][11]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[5][10]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[3][25]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[3][26]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[3][24]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[3][22]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[3][23]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[3][21]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[3][19]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[3][20]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[3][15]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[3][13]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[3][14]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[3][18]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[3][16]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[3][17]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[4][25]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[4][26]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[4][24]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[4][22]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[4][23]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[4][21]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[4][19]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[4][20]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[4][15]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[4][13]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[4][14]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[4][18]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[4][16]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[4][17]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[6][12]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[6][11]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[6][10]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[6][25]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[6][26]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[6][24]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[6][22]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[6][23]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[6][21]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[6][19]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[6][20]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[6][15]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[6][13]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[6][14]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[6][18]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[6][16]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[6][17]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[7][26]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[7][24]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[7][25]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[7][23]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[7][21]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[7][22]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[7][20]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[7][18]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[7][19]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[7][17]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[7][15]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[7][16]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[7][11]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[7][10]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[7][14]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[7][12]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[7][13]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[2][25]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[2][26]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[2][24]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[2][22]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[2][23]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[2][21]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[2][19]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[2][20]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[2][15]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[2][13]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[2][14]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[2][18]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[2][16]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[2][17]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[1][25]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[1][26]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[1][24]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[1][22]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[1][23]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[1][21]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[1][19]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[1][20]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[1][15]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[1][13]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[1][14]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[1][18]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[1][16]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[1][17]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[0][2]~q ;
wire \state_machine_inst|to_row_addr_r[0]~q ;
wire \state_machine_inst|to_row_addr_r[1]~q ;
wire \state_machine_inst|to_col_addr_r[2]~q ;
wire \state_machine_inst|to_row_addr_r[2]~q ;
wire \state_machine_inst|to_col_addr_r[3]~q ;
wire \state_machine_inst|to_row_addr_r[3]~q ;
wire \state_machine_inst|to_col_addr_r[4]~q ;
wire \state_machine_inst|to_row_addr_r[4]~q ;
wire \state_machine_inst|to_col_addr_r[5]~q ;
wire \state_machine_inst|to_row_addr_r[5]~q ;
wire \state_machine_inst|to_col_addr_r[6]~q ;
wire \state_machine_inst|to_row_addr_r[6]~q ;
wire \state_machine_inst|to_col_addr_r[7]~q ;
wire \state_machine_inst|to_row_addr_r[7]~q ;
wire \state_machine_inst|to_col_addr_r[8]~q ;
wire \state_machine_inst|to_row_addr_r[8]~q ;
wire \state_machine_inst|to_col_addr_r[9]~q ;
wire \state_machine_inst|to_row_addr_r[9]~q ;
wire \state_machine_inst|to_row_addr_r[10]~q ;
wire \state_machine_inst|to_row_addr_r[11]~q ;
wire \state_machine_inst|to_row_addr_r[12]~q ;
wire \state_machine_inst|to_row_addr_r[13]~q ;
wire \input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[132] ;
wire \input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[140] ;
wire \input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[128] ;
wire \input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[136] ;
wire \input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[133] ;
wire \input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[141] ;
wire \input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[129] ;
wire \input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[137] ;
wire \input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[134] ;
wire \input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[142] ;
wire \input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[130] ;
wire \input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[138] ;
wire \input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[135] ;
wire \input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[143] ;
wire \input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[131] ;
wire \input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[139] ;
wire \input_if_inst|cmd_queue_inst|pipe[0][3]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[0][4]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[0][5]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[0][6]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[0][7]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[0][8]~q ;
wire \input_if_inst|cmd_queue_inst|pipe[0][9]~q ;
wire \input_if_inst|cmd_gen_inst|hold_ready~q ;
wire \input_if_inst|cmd_queue_inst|pipefull[7]~q ;
wire \input_if_inst|internal_ready~0_combout ;
wire \input_if_inst|avalon_if_inst|avalon_write_req~combout ;
wire \clock_and_reset_inst|reset_sync_inst|reset_reg[4]~q ;
wire \state_machine_inst|fetch~q ;
wire \input_if_inst|cmd_gen_inst|read_req~0_combout ;
wire \input_if_inst|cmd_gen_inst|write_req~1_combout ;
wire \input_if_inst|cmd_queue_inst|pipefull[6]~q ;
wire \clock_and_reset_inst|reset_sync_inst|reset_reg[5]~q ;
wire \clock_and_reset_inst|reset_sync_inst|reset_reg[7]~q ;
wire \afi_block_inst|ecc_wdata_fifo_read~q ;
wire \clock_and_reset_inst|reset_sync_inst|reset_reg[3]~q ;
wire \state_machine_inst|do_precharge_all_r~q ;
wire \bank_timer_wrapper_inst|bypass_inst|out_cs_can_refresh[0]~q ;
wire \clock_and_reset_inst|reset_sync_inst|reset_reg[14]~q ;
wire \state_machine_inst|always38~0_combout ;
wire \input_if_inst|cmd_queue_inst|pipefull[0]~q ;
wire \state_machine_inst|do_refresh_r~q ;
wire \bank_timer_wrapper_inst|timing_param_inst|add_lat_on~q ;
wire \bank_timer_wrapper_inst|bypass_inst|out_cmd_can_activate[0]~q ;
wire \bank_timer_wrapper_inst|bypass_inst|out_cmd_bank_is_open[0]~q ;
wire \bank_timer_wrapper_inst|bank_timer_inst|can_al_activate_write~q ;
wire \state_machine_inst|to_chip_r[0]~q ;
wire \state_machine_inst|always38~3_combout ;
wire \state_machine_inst|to_bank_addr_r[2]~q ;
wire \state_machine_inst|current_bank[2]~q ;
wire \state_machine_inst|to_bank_addr_r[0]~q ;
wire \state_machine_inst|current_bank[0]~q ;
wire \state_machine_inst|to_bank_addr_r[1]~q ;
wire \state_machine_inst|current_bank[1]~q ;
wire \state_machine_inst|always38~4_combout ;
wire \bank_timer_wrapper_inst|bypass_inst|out_cmd_can_write[0]~q ;
wire \bank_timer_wrapper_inst|bank_timer_inst|can_al_activate_read~q ;
wire \bank_timer_wrapper_inst|bypass_inst|out_cmd_can_read[0]~q ;
wire \input_if_inst|cmd_queue_inst|pipefull[5]~q ;
wire \clock_and_reset_inst|reset_sync_inst|reset_reg[16]~q ;
wire \bank_timer_wrapper_inst|bypass_inst|out_cs_all_banks_closed[0]~q ;
wire \bank_timer_wrapper_inst|bypass_inst|out_cs_can_precharge_all[0]~q ;
wire \state_machine_inst|do_activate_r~q ;
wire \clock_and_reset_inst|reset_sync_inst|reset_reg[11]~q ;
wire \input_if_inst|cmd_queue_inst|pipefull[1]~q ;
wire \clock_and_reset_inst|reset_sync_inst|reset_reg[9]~q ;
wire \clock_and_reset_inst|reset_sync_inst|reset_reg[12]~q ;
wire \bank_timer_wrapper_inst|bypass_inst|out_cmd_can_activate[2]~q ;
wire \bank_timer_wrapper_inst|bypass_inst|out_cmd_bank_is_open[2]~q ;
wire \bank_timer_wrapper_inst|bypass_inst|out_cmd_can_activate[3]~q ;
wire \bank_timer_wrapper_inst|bypass_inst|out_cmd_bank_is_open[3]~q ;
wire \bank_timer_wrapper_inst|bypass_inst|out_cmd_can_activate[4]~q ;
wire \bank_timer_wrapper_inst|bypass_inst|out_cmd_bank_is_open[4]~q ;
wire \bank_timer_wrapper_inst|bypass_inst|out_cmd_can_activate[1]~q ;
wire \bank_timer_wrapper_inst|bypass_inst|out_cmd_bank_is_open[1]~q ;
wire \clock_and_reset_inst|reset_sync_inst|reset_reg[8]~q ;
wire \input_if_inst|cmd_queue_inst|pipefull[4]~q ;
wire \input_if_inst|cmd_queue_inst|pipefull[2]~q ;
wire \clock_and_reset_inst|reset_sync_inst|reset_reg[10]~q ;
wire \input_if_inst|cmd_queue_inst|pipefull[3]~q ;
wire \bank_timer_wrapper_inst|bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[2].bank_timer_info_inst|always1~0_combout ;
wire \clock_and_reset_inst|reset_sync_inst|reset_reg[15]~q ;


ddr3_int_alt_ddrx_state_machine state_machine_inst(
	.ctl_clk(clk_0),
	.auto_refresh_logic_per_chip0int_refresh_req(\bank_timer_wrapper_inst|rank_monitor_inst|auto_refresh_logic_per_chip[0].int_refresh_req~q ),
	.out_cmd_info_valid_0(\bank_timer_wrapper_inst|bypass_inst|out_cmd_info_valid[0]~q ),
	.do_read_r1(do_read_r),
	.do_auto_precharge_r1(\state_machine_inst|do_auto_precharge_r~q ),
	.do_write_r1(\state_machine_inst|do_write_r~q ),
	.out_cmd_info_valid_2(\bank_timer_wrapper_inst|bypass_inst|out_cmd_info_valid[2]~q ),
	.out_cmd_info_valid_3(\bank_timer_wrapper_inst|bypass_inst|out_cmd_info_valid[3]~q ),
	.out_cmd_info_valid_4(\bank_timer_wrapper_inst|bypass_inst|out_cmd_info_valid[4]~q ),
	.out_cmd_info_valid_1(\bank_timer_wrapper_inst|bypass_inst|out_cmd_info_valid[1]~q ),
	.pipe_10_0(\input_if_inst|cmd_queue_inst|pipe[0][10]~q ),
	.pipe_12_0(\input_if_inst|cmd_queue_inst|pipe[0][12]~q ),
	.pipe_11_0(\input_if_inst|cmd_queue_inst|pipe[0][11]~q ),
	.pipe_32_0(\input_if_inst|cmd_queue_inst|pipe[0][32]~q ),
	.pipe_12_2(\input_if_inst|cmd_queue_inst|pipe[2][12]~q ),
	.pipe_12_3(\input_if_inst|cmd_queue_inst|pipe[3][12]~q ),
	.pipe_12_1(\input_if_inst|cmd_queue_inst|pipe[1][12]~q ),
	.pipe_10_2(\input_if_inst|cmd_queue_inst|pipe[2][10]~q ),
	.pipe_10_3(\input_if_inst|cmd_queue_inst|pipe[3][10]~q ),
	.pipe_10_1(\input_if_inst|cmd_queue_inst|pipe[1][10]~q ),
	.pipe_11_2(\input_if_inst|cmd_queue_inst|pipe[2][11]~q ),
	.pipe_11_3(\input_if_inst|cmd_queue_inst|pipe[3][11]~q ),
	.pipe_11_1(\input_if_inst|cmd_queue_inst|pipe[1][11]~q ),
	.pipe_29_0(\input_if_inst|cmd_queue_inst|pipe[0][29]~q ),
	.pipe_28_0(\input_if_inst|cmd_queue_inst|pipe[0][28]~q ),
	.pipe_33_0(\input_if_inst|cmd_queue_inst|pipe[0][33]~q ),
	.do_burst_chop_r1(\state_machine_inst|do_burst_chop_r~q ),
	.pipe_12_4(\input_if_inst|cmd_queue_inst|pipe[4][12]~q ),
	.pipe_11_4(\input_if_inst|cmd_queue_inst|pipe[4][11]~q ),
	.pipe_10_4(\input_if_inst|cmd_queue_inst|pipe[4][10]~q ),
	.pipe_25_5(\input_if_inst|cmd_queue_inst|pipe[5][25]~q ),
	.pipe_25_0(\input_if_inst|cmd_queue_inst|pipe[0][25]~q ),
	.pipe_26_5(\input_if_inst|cmd_queue_inst|pipe[5][26]~q ),
	.pipe_26_0(\input_if_inst|cmd_queue_inst|pipe[0][26]~q ),
	.pipe_24_5(\input_if_inst|cmd_queue_inst|pipe[5][24]~q ),
	.pipe_24_0(\input_if_inst|cmd_queue_inst|pipe[0][24]~q ),
	.pipe_22_5(\input_if_inst|cmd_queue_inst|pipe[5][22]~q ),
	.pipe_22_0(\input_if_inst|cmd_queue_inst|pipe[0][22]~q ),
	.pipe_23_5(\input_if_inst|cmd_queue_inst|pipe[5][23]~q ),
	.pipe_23_0(\input_if_inst|cmd_queue_inst|pipe[0][23]~q ),
	.pipe_21_5(\input_if_inst|cmd_queue_inst|pipe[5][21]~q ),
	.pipe_21_0(\input_if_inst|cmd_queue_inst|pipe[0][21]~q ),
	.pipe_19_5(\input_if_inst|cmd_queue_inst|pipe[5][19]~q ),
	.pipe_19_0(\input_if_inst|cmd_queue_inst|pipe[0][19]~q ),
	.pipe_20_5(\input_if_inst|cmd_queue_inst|pipe[5][20]~q ),
	.pipe_20_0(\input_if_inst|cmd_queue_inst|pipe[0][20]~q ),
	.pipe_15_5(\input_if_inst|cmd_queue_inst|pipe[5][15]~q ),
	.pipe_15_0(\input_if_inst|cmd_queue_inst|pipe[0][15]~q ),
	.pipe_13_5(\input_if_inst|cmd_queue_inst|pipe[5][13]~q ),
	.pipe_13_0(\input_if_inst|cmd_queue_inst|pipe[0][13]~q ),
	.pipe_14_5(\input_if_inst|cmd_queue_inst|pipe[5][14]~q ),
	.pipe_14_0(\input_if_inst|cmd_queue_inst|pipe[0][14]~q ),
	.pipe_18_5(\input_if_inst|cmd_queue_inst|pipe[5][18]~q ),
	.pipe_18_0(\input_if_inst|cmd_queue_inst|pipe[0][18]~q ),
	.pipe_16_5(\input_if_inst|cmd_queue_inst|pipe[5][16]~q ),
	.pipe_16_0(\input_if_inst|cmd_queue_inst|pipe[0][16]~q ),
	.pipe_17_5(\input_if_inst|cmd_queue_inst|pipe[5][17]~q ),
	.pipe_17_0(\input_if_inst|cmd_queue_inst|pipe[0][17]~q ),
	.pipe_12_5(\input_if_inst|cmd_queue_inst|pipe[5][12]~q ),
	.pipe_11_5(\input_if_inst|cmd_queue_inst|pipe[5][11]~q ),
	.pipe_10_5(\input_if_inst|cmd_queue_inst|pipe[5][10]~q ),
	.pipe_25_3(\input_if_inst|cmd_queue_inst|pipe[3][25]~q ),
	.pipe_26_3(\input_if_inst|cmd_queue_inst|pipe[3][26]~q ),
	.pipe_24_3(\input_if_inst|cmd_queue_inst|pipe[3][24]~q ),
	.pipe_22_3(\input_if_inst|cmd_queue_inst|pipe[3][22]~q ),
	.pipe_23_3(\input_if_inst|cmd_queue_inst|pipe[3][23]~q ),
	.pipe_21_3(\input_if_inst|cmd_queue_inst|pipe[3][21]~q ),
	.pipe_19_3(\input_if_inst|cmd_queue_inst|pipe[3][19]~q ),
	.pipe_20_3(\input_if_inst|cmd_queue_inst|pipe[3][20]~q ),
	.pipe_15_3(\input_if_inst|cmd_queue_inst|pipe[3][15]~q ),
	.pipe_13_3(\input_if_inst|cmd_queue_inst|pipe[3][13]~q ),
	.pipe_14_3(\input_if_inst|cmd_queue_inst|pipe[3][14]~q ),
	.pipe_18_3(\input_if_inst|cmd_queue_inst|pipe[3][18]~q ),
	.pipe_16_3(\input_if_inst|cmd_queue_inst|pipe[3][16]~q ),
	.pipe_17_3(\input_if_inst|cmd_queue_inst|pipe[3][17]~q ),
	.pipe_25_4(\input_if_inst|cmd_queue_inst|pipe[4][25]~q ),
	.pipe_26_4(\input_if_inst|cmd_queue_inst|pipe[4][26]~q ),
	.pipe_24_4(\input_if_inst|cmd_queue_inst|pipe[4][24]~q ),
	.pipe_22_4(\input_if_inst|cmd_queue_inst|pipe[4][22]~q ),
	.pipe_23_4(\input_if_inst|cmd_queue_inst|pipe[4][23]~q ),
	.pipe_21_4(\input_if_inst|cmd_queue_inst|pipe[4][21]~q ),
	.pipe_19_4(\input_if_inst|cmd_queue_inst|pipe[4][19]~q ),
	.pipe_20_4(\input_if_inst|cmd_queue_inst|pipe[4][20]~q ),
	.pipe_15_4(\input_if_inst|cmd_queue_inst|pipe[4][15]~q ),
	.pipe_13_4(\input_if_inst|cmd_queue_inst|pipe[4][13]~q ),
	.pipe_14_4(\input_if_inst|cmd_queue_inst|pipe[4][14]~q ),
	.pipe_18_4(\input_if_inst|cmd_queue_inst|pipe[4][18]~q ),
	.pipe_16_4(\input_if_inst|cmd_queue_inst|pipe[4][16]~q ),
	.pipe_17_4(\input_if_inst|cmd_queue_inst|pipe[4][17]~q ),
	.pipe_12_6(\input_if_inst|cmd_queue_inst|pipe[6][12]~q ),
	.pipe_11_6(\input_if_inst|cmd_queue_inst|pipe[6][11]~q ),
	.pipe_10_6(\input_if_inst|cmd_queue_inst|pipe[6][10]~q ),
	.pipe_25_6(\input_if_inst|cmd_queue_inst|pipe[6][25]~q ),
	.pipe_26_6(\input_if_inst|cmd_queue_inst|pipe[6][26]~q ),
	.pipe_24_6(\input_if_inst|cmd_queue_inst|pipe[6][24]~q ),
	.pipe_22_6(\input_if_inst|cmd_queue_inst|pipe[6][22]~q ),
	.pipe_23_6(\input_if_inst|cmd_queue_inst|pipe[6][23]~q ),
	.pipe_21_6(\input_if_inst|cmd_queue_inst|pipe[6][21]~q ),
	.pipe_19_6(\input_if_inst|cmd_queue_inst|pipe[6][19]~q ),
	.pipe_20_6(\input_if_inst|cmd_queue_inst|pipe[6][20]~q ),
	.pipe_15_6(\input_if_inst|cmd_queue_inst|pipe[6][15]~q ),
	.pipe_13_6(\input_if_inst|cmd_queue_inst|pipe[6][13]~q ),
	.pipe_14_6(\input_if_inst|cmd_queue_inst|pipe[6][14]~q ),
	.pipe_18_6(\input_if_inst|cmd_queue_inst|pipe[6][18]~q ),
	.pipe_16_6(\input_if_inst|cmd_queue_inst|pipe[6][16]~q ),
	.pipe_17_6(\input_if_inst|cmd_queue_inst|pipe[6][17]~q ),
	.pipe_26_7(\input_if_inst|cmd_queue_inst|pipe[7][26]~q ),
	.pipe_24_7(\input_if_inst|cmd_queue_inst|pipe[7][24]~q ),
	.pipe_25_7(\input_if_inst|cmd_queue_inst|pipe[7][25]~q ),
	.pipe_23_7(\input_if_inst|cmd_queue_inst|pipe[7][23]~q ),
	.pipe_21_7(\input_if_inst|cmd_queue_inst|pipe[7][21]~q ),
	.pipe_22_7(\input_if_inst|cmd_queue_inst|pipe[7][22]~q ),
	.pipe_20_7(\input_if_inst|cmd_queue_inst|pipe[7][20]~q ),
	.pipe_18_7(\input_if_inst|cmd_queue_inst|pipe[7][18]~q ),
	.pipe_19_7(\input_if_inst|cmd_queue_inst|pipe[7][19]~q ),
	.pipe_17_7(\input_if_inst|cmd_queue_inst|pipe[7][17]~q ),
	.pipe_15_7(\input_if_inst|cmd_queue_inst|pipe[7][15]~q ),
	.pipe_16_7(\input_if_inst|cmd_queue_inst|pipe[7][16]~q ),
	.pipe_11_7(\input_if_inst|cmd_queue_inst|pipe[7][11]~q ),
	.pipe_10_7(\input_if_inst|cmd_queue_inst|pipe[7][10]~q ),
	.pipe_14_7(\input_if_inst|cmd_queue_inst|pipe[7][14]~q ),
	.pipe_12_7(\input_if_inst|cmd_queue_inst|pipe[7][12]~q ),
	.pipe_13_7(\input_if_inst|cmd_queue_inst|pipe[7][13]~q ),
	.pipe_25_2(\input_if_inst|cmd_queue_inst|pipe[2][25]~q ),
	.pipe_26_2(\input_if_inst|cmd_queue_inst|pipe[2][26]~q ),
	.pipe_24_2(\input_if_inst|cmd_queue_inst|pipe[2][24]~q ),
	.pipe_22_2(\input_if_inst|cmd_queue_inst|pipe[2][22]~q ),
	.pipe_23_2(\input_if_inst|cmd_queue_inst|pipe[2][23]~q ),
	.pipe_21_2(\input_if_inst|cmd_queue_inst|pipe[2][21]~q ),
	.pipe_19_2(\input_if_inst|cmd_queue_inst|pipe[2][19]~q ),
	.pipe_20_2(\input_if_inst|cmd_queue_inst|pipe[2][20]~q ),
	.pipe_15_2(\input_if_inst|cmd_queue_inst|pipe[2][15]~q ),
	.pipe_13_2(\input_if_inst|cmd_queue_inst|pipe[2][13]~q ),
	.pipe_14_2(\input_if_inst|cmd_queue_inst|pipe[2][14]~q ),
	.pipe_18_2(\input_if_inst|cmd_queue_inst|pipe[2][18]~q ),
	.pipe_16_2(\input_if_inst|cmd_queue_inst|pipe[2][16]~q ),
	.pipe_17_2(\input_if_inst|cmd_queue_inst|pipe[2][17]~q ),
	.pipe_25_1(\input_if_inst|cmd_queue_inst|pipe[1][25]~q ),
	.pipe_26_1(\input_if_inst|cmd_queue_inst|pipe[1][26]~q ),
	.pipe_24_1(\input_if_inst|cmd_queue_inst|pipe[1][24]~q ),
	.pipe_22_1(\input_if_inst|cmd_queue_inst|pipe[1][22]~q ),
	.pipe_23_1(\input_if_inst|cmd_queue_inst|pipe[1][23]~q ),
	.pipe_21_1(\input_if_inst|cmd_queue_inst|pipe[1][21]~q ),
	.pipe_19_1(\input_if_inst|cmd_queue_inst|pipe[1][19]~q ),
	.pipe_20_1(\input_if_inst|cmd_queue_inst|pipe[1][20]~q ),
	.pipe_15_1(\input_if_inst|cmd_queue_inst|pipe[1][15]~q ),
	.pipe_13_1(\input_if_inst|cmd_queue_inst|pipe[1][13]~q ),
	.pipe_14_1(\input_if_inst|cmd_queue_inst|pipe[1][14]~q ),
	.pipe_18_1(\input_if_inst|cmd_queue_inst|pipe[1][18]~q ),
	.pipe_16_1(\input_if_inst|cmd_queue_inst|pipe[1][16]~q ),
	.pipe_17_1(\input_if_inst|cmd_queue_inst|pipe[1][17]~q ),
	.pipe_2_0(\input_if_inst|cmd_queue_inst|pipe[0][2]~q ),
	.to_row_addr_r_0(\state_machine_inst|to_row_addr_r[0]~q ),
	.to_row_addr_r_1(\state_machine_inst|to_row_addr_r[1]~q ),
	.to_col_addr_r_2(\state_machine_inst|to_col_addr_r[2]~q ),
	.to_row_addr_r_2(\state_machine_inst|to_row_addr_r[2]~q ),
	.to_col_addr_r_3(\state_machine_inst|to_col_addr_r[3]~q ),
	.to_row_addr_r_3(\state_machine_inst|to_row_addr_r[3]~q ),
	.to_col_addr_r_4(\state_machine_inst|to_col_addr_r[4]~q ),
	.to_row_addr_r_4(\state_machine_inst|to_row_addr_r[4]~q ),
	.to_col_addr_r_5(\state_machine_inst|to_col_addr_r[5]~q ),
	.to_row_addr_r_5(\state_machine_inst|to_row_addr_r[5]~q ),
	.to_col_addr_r_6(\state_machine_inst|to_col_addr_r[6]~q ),
	.to_row_addr_r_6(\state_machine_inst|to_row_addr_r[6]~q ),
	.to_col_addr_r_7(\state_machine_inst|to_col_addr_r[7]~q ),
	.to_row_addr_r_7(\state_machine_inst|to_row_addr_r[7]~q ),
	.to_col_addr_r_8(\state_machine_inst|to_col_addr_r[8]~q ),
	.to_row_addr_r_8(\state_machine_inst|to_row_addr_r[8]~q ),
	.to_col_addr_r_9(\state_machine_inst|to_col_addr_r[9]~q ),
	.to_row_addr_r_9(\state_machine_inst|to_row_addr_r[9]~q ),
	.to_row_addr_r_10(\state_machine_inst|to_row_addr_r[10]~q ),
	.to_row_addr_r_11(\state_machine_inst|to_row_addr_r[11]~q ),
	.to_row_addr_r_12(\state_machine_inst|to_row_addr_r[12]~q ),
	.to_row_addr_r_13(\state_machine_inst|to_row_addr_r[13]~q ),
	.pipe_3_0(\input_if_inst|cmd_queue_inst|pipe[0][3]~q ),
	.pipe_4_0(\input_if_inst|cmd_queue_inst|pipe[0][4]~q ),
	.pipe_5_0(\input_if_inst|cmd_queue_inst|pipe[0][5]~q ),
	.pipe_6_0(\input_if_inst|cmd_queue_inst|pipe[0][6]~q ),
	.pipe_7_0(\input_if_inst|cmd_queue_inst|pipe[0][7]~q ),
	.pipe_8_0(\input_if_inst|cmd_queue_inst|pipe[0][8]~q ),
	.pipe_9_0(\input_if_inst|cmd_queue_inst|pipe[0][9]~q ),
	.hold_ready(\input_if_inst|cmd_gen_inst|hold_ready~q ),
	.pipefull_7(\input_if_inst|cmd_queue_inst|pipefull[7]~q ),
	.int_refresh_ack1(int_refresh_ack),
	.ctl_init_success(ctl_init_success),
	.internal_ready(\input_if_inst|internal_ready~0_combout ),
	.avalon_write_req(\input_if_inst|avalon_if_inst|avalon_write_req~combout ),
	.fetch1(\state_machine_inst|fetch~q ),
	.read_req(\input_if_inst|cmd_gen_inst|read_req~0_combout ),
	.write_req(\input_if_inst|cmd_gen_inst|write_req~1_combout ),
	.pipefull_6(\input_if_inst|cmd_queue_inst|pipefull[6]~q ),
	.do_precharge_all_r1(\state_machine_inst|do_precharge_all_r~q ),
	.out_cs_can_refresh_0(\bank_timer_wrapper_inst|bypass_inst|out_cs_can_refresh[0]~q ),
	.ctl_reset_n(\clock_and_reset_inst|reset_sync_inst|reset_reg[14]~q ),
	.always38(\state_machine_inst|always38~0_combout ),
	.pipefull_0(\input_if_inst|cmd_queue_inst|pipefull[0]~q ),
	.do_refresh_r1(\state_machine_inst|do_refresh_r~q ),
	.add_lat_on(\bank_timer_wrapper_inst|timing_param_inst|add_lat_on~q ),
	.out_cmd_can_activate_0(\bank_timer_wrapper_inst|bypass_inst|out_cmd_can_activate[0]~q ),
	.out_cmd_bank_is_open_0(\bank_timer_wrapper_inst|bypass_inst|out_cmd_bank_is_open[0]~q ),
	.can_al_activate_write(\bank_timer_wrapper_inst|bank_timer_inst|can_al_activate_write~q ),
	.to_chip_r_0(\state_machine_inst|to_chip_r[0]~q ),
	.always381(\state_machine_inst|always38~3_combout ),
	.to_bank_addr_r_2(\state_machine_inst|to_bank_addr_r[2]~q ),
	.current_bank_2(\state_machine_inst|current_bank[2]~q ),
	.to_bank_addr_r_0(\state_machine_inst|to_bank_addr_r[0]~q ),
	.current_bank_0(\state_machine_inst|current_bank[0]~q ),
	.to_bank_addr_r_1(\state_machine_inst|to_bank_addr_r[1]~q ),
	.current_bank_1(\state_machine_inst|current_bank[1]~q ),
	.always382(\state_machine_inst|always38~4_combout ),
	.out_cmd_can_write_0(\bank_timer_wrapper_inst|bypass_inst|out_cmd_can_write[0]~q ),
	.can_al_activate_read(\bank_timer_wrapper_inst|bank_timer_inst|can_al_activate_read~q ),
	.out_cmd_can_read_0(\bank_timer_wrapper_inst|bypass_inst|out_cmd_can_read[0]~q ),
	.pipefull_5(\input_if_inst|cmd_queue_inst|pipefull[5]~q ),
	.rdwr_data_valid_r1(rdwr_data_valid_r),
	.out_cs_all_banks_closed_0(\bank_timer_wrapper_inst|bypass_inst|out_cs_all_banks_closed[0]~q ),
	.out_cs_can_precharge_all_0(\bank_timer_wrapper_inst|bypass_inst|out_cs_can_precharge_all[0]~q ),
	.do_activate_r1(\state_machine_inst|do_activate_r~q ),
	.pipefull_1(\input_if_inst|cmd_queue_inst|pipefull[1]~q ),
	.out_cmd_can_activate_2(\bank_timer_wrapper_inst|bypass_inst|out_cmd_can_activate[2]~q ),
	.out_cmd_bank_is_open_2(\bank_timer_wrapper_inst|bypass_inst|out_cmd_bank_is_open[2]~q ),
	.out_cmd_can_activate_3(\bank_timer_wrapper_inst|bypass_inst|out_cmd_can_activate[3]~q ),
	.out_cmd_bank_is_open_3(\bank_timer_wrapper_inst|bypass_inst|out_cmd_bank_is_open[3]~q ),
	.out_cmd_can_activate_4(\bank_timer_wrapper_inst|bypass_inst|out_cmd_can_activate[4]~q ),
	.out_cmd_bank_is_open_4(\bank_timer_wrapper_inst|bypass_inst|out_cmd_bank_is_open[4]~q ),
	.out_cmd_can_activate_1(\bank_timer_wrapper_inst|bypass_inst|out_cmd_can_activate[1]~q ),
	.out_cmd_bank_is_open_1(\bank_timer_wrapper_inst|bypass_inst|out_cmd_bank_is_open[1]~q ),
	.pipefull_4(\input_if_inst|cmd_queue_inst|pipefull[4]~q ),
	.pipefull_2(\input_if_inst|cmd_queue_inst|pipefull[2]~q ),
	.pipefull_3(\input_if_inst|cmd_queue_inst|pipefull[3]~q ),
	.local_write_req(local_write_req));

ddr3_int_alt_ddrx_addr_cmd addr_cmd_inst(
	.ctl_clk(clk_0),
	.do_read_r(do_read_r),
	.do_auto_precharge_r(\state_machine_inst|do_auto_precharge_r~q ),
	.do_write_r(\state_machine_inst|do_write_r~q ),
	.do_burst_chop_r(\state_machine_inst|do_burst_chop_r~q ),
	.to_row_addr_r_0(\state_machine_inst|to_row_addr_r[0]~q ),
	.to_row_addr_r_1(\state_machine_inst|to_row_addr_r[1]~q ),
	.to_col_addr_r_2(\state_machine_inst|to_col_addr_r[2]~q ),
	.to_row_addr_r_2(\state_machine_inst|to_row_addr_r[2]~q ),
	.to_col_addr_r_3(\state_machine_inst|to_col_addr_r[3]~q ),
	.to_row_addr_r_3(\state_machine_inst|to_row_addr_r[3]~q ),
	.to_col_addr_r_4(\state_machine_inst|to_col_addr_r[4]~q ),
	.to_row_addr_r_4(\state_machine_inst|to_row_addr_r[4]~q ),
	.to_col_addr_r_5(\state_machine_inst|to_col_addr_r[5]~q ),
	.to_row_addr_r_5(\state_machine_inst|to_row_addr_r[5]~q ),
	.to_col_addr_r_6(\state_machine_inst|to_col_addr_r[6]~q ),
	.to_row_addr_r_6(\state_machine_inst|to_row_addr_r[6]~q ),
	.to_col_addr_r_7(\state_machine_inst|to_col_addr_r[7]~q ),
	.to_row_addr_r_7(\state_machine_inst|to_row_addr_r[7]~q ),
	.to_col_addr_r_8(\state_machine_inst|to_col_addr_r[8]~q ),
	.to_row_addr_r_8(\state_machine_inst|to_row_addr_r[8]~q ),
	.to_col_addr_r_9(\state_machine_inst|to_col_addr_r[9]~q ),
	.to_row_addr_r_9(\state_machine_inst|to_row_addr_r[9]~q ),
	.to_row_addr_r_10(\state_machine_inst|to_row_addr_r[10]~q ),
	.to_row_addr_r_11(\state_machine_inst|to_row_addr_r[11]~q ),
	.to_row_addr_r_12(\state_machine_inst|to_row_addr_r[12]~q ),
	.to_row_addr_r_13(\state_machine_inst|to_row_addr_r[13]~q ),
	.ctl_init_success(ctl_init_success),
	.do_precharge_all_r(\state_machine_inst|do_precharge_all_r~q ),
	.do_refresh_r(\state_machine_inst|do_refresh_r~q ),
	.to_chip_r_0(\state_machine_inst|to_chip_r[0]~q ),
	.to_bank_addr_r_2(\state_machine_inst|to_bank_addr_r[2]~q ),
	.to_bank_addr_r_0(\state_machine_inst|to_bank_addr_r[0]~q ),
	.to_bank_addr_r_1(\state_machine_inst|to_bank_addr_r[1]~q ),
	.do_activate_r(\state_machine_inst|do_activate_r~q ),
	.always1(\bank_timer_wrapper_inst|bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[2].bank_timer_info_inst|always1~0_combout ),
	.afi_cs_n_1(afi_cs_n_1),
	.int_cke_r_0(int_cke_r_0),
	.afi_addr_0(afi_addr_0),
	.afi_addr_1(afi_addr_1),
	.afi_addr_2(afi_addr_2),
	.afi_addr_3(afi_addr_3),
	.afi_addr_4(afi_addr_4),
	.afi_addr_5(afi_addr_5),
	.afi_addr_6(afi_addr_6),
	.afi_addr_7(afi_addr_7),
	.afi_addr_8(afi_addr_8),
	.afi_addr_9(afi_addr_9),
	.afi_addr_10(afi_addr_10),
	.afi_addr_11(afi_addr_11),
	.afi_addr_12(afi_addr_12),
	.afi_addr_13(afi_addr_13),
	.afi_ba_0(afi_ba_0),
	.afi_ba_1(afi_ba_1),
	.afi_ba_2(afi_ba_2),
	.afi_ras_n_0(afi_ras_n_0),
	.afi_cas_n_0(afi_cas_n_0),
	.afi_we_n_0(afi_we_n_0),
	.ctl_reset_n(\clock_and_reset_inst|reset_sync_inst|reset_reg[15]~q ));

ddr3_int_alt_ddrx_afi_block afi_block_inst(
	.ctl_clk(clk_0),
	.do_read_r(do_read_r),
	.do_write_r(\state_machine_inst|do_write_r~q ),
	.do_burst_chop_r(\state_machine_inst|do_burst_chop_r~q ),
	.q_b_132(\input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[132] ),
	.q_b_140(\input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[140] ),
	.q_b_128(\input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[128] ),
	.q_b_136(\input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[136] ),
	.q_b_133(\input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[133] ),
	.q_b_141(\input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[141] ),
	.q_b_129(\input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[129] ),
	.q_b_137(\input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[137] ),
	.q_b_134(\input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[134] ),
	.q_b_142(\input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[142] ),
	.q_b_130(\input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[130] ),
	.q_b_138(\input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[138] ),
	.q_b_135(\input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[135] ),
	.q_b_143(\input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[143] ),
	.q_b_131(\input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[131] ),
	.q_b_139(\input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[139] ),
	.ecc_wdata_fifo_read1(\afi_block_inst|ecc_wdata_fifo_read~q ),
	.rdwr_data_valid(rdwr_data_valid_r),
	.ctl_reset_n(\clock_and_reset_inst|reset_sync_inst|reset_reg[16]~q ),
	.doing_read1(doing_read),
	.wd_lat_2(wd_lat_2),
	.afi_wlat({wd_lat_4,wd_lat_3,gnd,wd_lat_1,gnd}),
	.wd_lat_0(wd_lat_0),
	.afi_dm_4(afi_dm_4),
	.afi_dm_12(afi_dm_12),
	.afi_dm_0(afi_dm_0),
	.afi_dm_8(afi_dm_8),
	.afi_dm_5(afi_dm_5),
	.afi_dm_13(afi_dm_13),
	.afi_dm_1(afi_dm_1),
	.afi_dm_9(afi_dm_9),
	.afi_dm_6(afi_dm_6),
	.afi_dm_14(afi_dm_14),
	.afi_dm_2(afi_dm_2),
	.afi_dm_10(afi_dm_10),
	.afi_dm_7(afi_dm_7),
	.afi_dm_15(afi_dm_15),
	.afi_dm_3(afi_dm_3),
	.afi_dm_11(afi_dm_11),
	.int_wdata_valid1(int_wdata_valid),
	.int_dqs_burst1(int_dqs_burst),
	.int_dqs_burst_hr1(int_dqs_burst_hr));

ddr3_int_alt_ddrx_bank_timer_wrapper bank_timer_wrapper_inst(
	.clk_0(clk_0),
	.auto_refresh_logic_per_chip0int_refresh_req(\bank_timer_wrapper_inst|rank_monitor_inst|auto_refresh_logic_per_chip[0].int_refresh_req~q ),
	.out_cmd_info_valid_0(\bank_timer_wrapper_inst|bypass_inst|out_cmd_info_valid[0]~q ),
	.do_read_r(do_read_r),
	.do_auto_precharge_r(\state_machine_inst|do_auto_precharge_r~q ),
	.do_write_r(\state_machine_inst|do_write_r~q ),
	.out_cmd_info_valid_2(\bank_timer_wrapper_inst|bypass_inst|out_cmd_info_valid[2]~q ),
	.out_cmd_info_valid_3(\bank_timer_wrapper_inst|bypass_inst|out_cmd_info_valid[3]~q ),
	.out_cmd_info_valid_4(\bank_timer_wrapper_inst|bypass_inst|out_cmd_info_valid[4]~q ),
	.out_cmd_info_valid_1(\bank_timer_wrapper_inst|bypass_inst|out_cmd_info_valid[1]~q ),
	.pipe_10_0(\input_if_inst|cmd_queue_inst|pipe[0][10]~q ),
	.pipe_12_0(\input_if_inst|cmd_queue_inst|pipe[0][12]~q ),
	.pipe_11_0(\input_if_inst|cmd_queue_inst|pipe[0][11]~q ),
	.pipe_12_2(\input_if_inst|cmd_queue_inst|pipe[2][12]~q ),
	.pipe_12_3(\input_if_inst|cmd_queue_inst|pipe[3][12]~q ),
	.pipe_12_1(\input_if_inst|cmd_queue_inst|pipe[1][12]~q ),
	.pipe_10_2(\input_if_inst|cmd_queue_inst|pipe[2][10]~q ),
	.pipe_10_3(\input_if_inst|cmd_queue_inst|pipe[3][10]~q ),
	.pipe_10_1(\input_if_inst|cmd_queue_inst|pipe[1][10]~q ),
	.pipe_11_2(\input_if_inst|cmd_queue_inst|pipe[2][11]~q ),
	.pipe_11_3(\input_if_inst|cmd_queue_inst|pipe[3][11]~q ),
	.pipe_11_1(\input_if_inst|cmd_queue_inst|pipe[1][11]~q ),
	.do_burst_chop_r(\state_machine_inst|do_burst_chop_r~q ),
	.pipe_12_4(\input_if_inst|cmd_queue_inst|pipe[4][12]~q ),
	.pipe_11_4(\input_if_inst|cmd_queue_inst|pipe[4][11]~q ),
	.pipe_10_4(\input_if_inst|cmd_queue_inst|pipe[4][10]~q ),
	.fetch(\state_machine_inst|fetch~q ),
	.do_precharge_all_r(\state_machine_inst|do_precharge_all_r~q ),
	.out_cs_can_refresh_0(\bank_timer_wrapper_inst|bypass_inst|out_cs_can_refresh[0]~q ),
	.pipefull_0(\input_if_inst|cmd_queue_inst|pipefull[0]~q ),
	.do_refresh_r(\state_machine_inst|do_refresh_r~q ),
	.add_lat_on(\bank_timer_wrapper_inst|timing_param_inst|add_lat_on~q ),
	.out_cmd_can_activate_0(\bank_timer_wrapper_inst|bypass_inst|out_cmd_can_activate[0]~q ),
	.out_cmd_bank_is_open_0(\bank_timer_wrapper_inst|bypass_inst|out_cmd_bank_is_open[0]~q ),
	.can_al_activate_write(\bank_timer_wrapper_inst|bank_timer_inst|can_al_activate_write~q ),
	.to_chip_r_0(\state_machine_inst|to_chip_r[0]~q ),
	.always38(\state_machine_inst|always38~3_combout ),
	.to_bank_addr_r_2(\state_machine_inst|to_bank_addr_r[2]~q ),
	.current_bank_2(\state_machine_inst|current_bank[2]~q ),
	.to_bank_addr_r_0(\state_machine_inst|to_bank_addr_r[0]~q ),
	.current_bank_0(\state_machine_inst|current_bank[0]~q ),
	.to_bank_addr_r_1(\state_machine_inst|to_bank_addr_r[1]~q ),
	.current_bank_1(\state_machine_inst|current_bank[1]~q ),
	.always381(\state_machine_inst|always38~4_combout ),
	.out_cmd_can_write_0(\bank_timer_wrapper_inst|bypass_inst|out_cmd_can_write[0]~q ),
	.can_al_activate_read(\bank_timer_wrapper_inst|bank_timer_inst|can_al_activate_read~q ),
	.out_cmd_can_read_0(\bank_timer_wrapper_inst|bypass_inst|out_cmd_can_read[0]~q ),
	.out_cs_all_banks_closed_0(\bank_timer_wrapper_inst|bypass_inst|out_cs_all_banks_closed[0]~q ),
	.out_cs_can_precharge_all_0(\bank_timer_wrapper_inst|bypass_inst|out_cs_can_precharge_all[0]~q ),
	.do_activate_r(\state_machine_inst|do_activate_r~q ),
	.reset_reg_11(\clock_and_reset_inst|reset_sync_inst|reset_reg[11]~q ),
	.pipefull_1(\input_if_inst|cmd_queue_inst|pipefull[1]~q ),
	.reset_reg_9(\clock_and_reset_inst|reset_sync_inst|reset_reg[9]~q ),
	.reset_reg_12(\clock_and_reset_inst|reset_sync_inst|reset_reg[12]~q ),
	.out_cmd_can_activate_2(\bank_timer_wrapper_inst|bypass_inst|out_cmd_can_activate[2]~q ),
	.out_cmd_bank_is_open_2(\bank_timer_wrapper_inst|bypass_inst|out_cmd_bank_is_open[2]~q ),
	.out_cmd_can_activate_3(\bank_timer_wrapper_inst|bypass_inst|out_cmd_can_activate[3]~q ),
	.out_cmd_bank_is_open_3(\bank_timer_wrapper_inst|bypass_inst|out_cmd_bank_is_open[3]~q ),
	.out_cmd_can_activate_4(\bank_timer_wrapper_inst|bypass_inst|out_cmd_can_activate[4]~q ),
	.out_cmd_bank_is_open_4(\bank_timer_wrapper_inst|bypass_inst|out_cmd_bank_is_open[4]~q ),
	.out_cmd_can_activate_1(\bank_timer_wrapper_inst|bypass_inst|out_cmd_can_activate[1]~q ),
	.out_cmd_bank_is_open_1(\bank_timer_wrapper_inst|bypass_inst|out_cmd_bank_is_open[1]~q ),
	.reset_reg_8(\clock_and_reset_inst|reset_sync_inst|reset_reg[8]~q ),
	.pipefull_4(\input_if_inst|cmd_queue_inst|pipefull[4]~q ),
	.pipefull_2(\input_if_inst|cmd_queue_inst|pipefull[2]~q ),
	.reset_reg_10(\clock_and_reset_inst|reset_sync_inst|reset_reg[10]~q ),
	.pipefull_3(\input_if_inst|cmd_queue_inst|pipefull[3]~q ),
	.always1(\bank_timer_wrapper_inst|bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[2].bank_timer_info_inst|always1~0_combout ),
	.GND_port(GND_port));

ddr3_int_alt_ddrx_clock_and_reset clock_and_reset_inst(
	.clk_0(clk_0),
	.reset_phy_clk_1x_n(reset_phy_clk_1x_n),
	.reset_reg_4(\clock_and_reset_inst|reset_sync_inst|reset_reg[4]~q ),
	.reset_reg_5(\clock_and_reset_inst|reset_sync_inst|reset_reg[5]~q ),
	.reset_reg_7(\clock_and_reset_inst|reset_sync_inst|reset_reg[7]~q ),
	.reset_reg_3(\clock_and_reset_inst|reset_sync_inst|reset_reg[3]~q ),
	.reset_reg_14(\clock_and_reset_inst|reset_sync_inst|reset_reg[14]~q ),
	.reset_reg_16(\clock_and_reset_inst|reset_sync_inst|reset_reg[16]~q ),
	.reset_reg_11(\clock_and_reset_inst|reset_sync_inst|reset_reg[11]~q ),
	.reset_reg_9(\clock_and_reset_inst|reset_sync_inst|reset_reg[9]~q ),
	.reset_reg_12(\clock_and_reset_inst|reset_sync_inst|reset_reg[12]~q ),
	.reset_reg_8(\clock_and_reset_inst|reset_sync_inst|reset_reg[8]~q ),
	.reset_reg_10(\clock_and_reset_inst|reset_sync_inst|reset_reg[10]~q ),
	.reset_reg_15(\clock_and_reset_inst|reset_sync_inst|reset_reg[15]~q ));

ddr3_int_alt_ddrx_input_if input_if_inst(
	.clk_0(clk_0),
	.pipe_10_0(\input_if_inst|cmd_queue_inst|pipe[0][10]~q ),
	.pipe_12_0(\input_if_inst|cmd_queue_inst|pipe[0][12]~q ),
	.pipe_11_0(\input_if_inst|cmd_queue_inst|pipe[0][11]~q ),
	.pipe_32_0(\input_if_inst|cmd_queue_inst|pipe[0][32]~q ),
	.pipe_12_2(\input_if_inst|cmd_queue_inst|pipe[2][12]~q ),
	.pipe_12_3(\input_if_inst|cmd_queue_inst|pipe[3][12]~q ),
	.pipe_12_1(\input_if_inst|cmd_queue_inst|pipe[1][12]~q ),
	.pipe_10_2(\input_if_inst|cmd_queue_inst|pipe[2][10]~q ),
	.pipe_10_3(\input_if_inst|cmd_queue_inst|pipe[3][10]~q ),
	.pipe_10_1(\input_if_inst|cmd_queue_inst|pipe[1][10]~q ),
	.pipe_11_2(\input_if_inst|cmd_queue_inst|pipe[2][11]~q ),
	.pipe_11_3(\input_if_inst|cmd_queue_inst|pipe[3][11]~q ),
	.pipe_11_1(\input_if_inst|cmd_queue_inst|pipe[1][11]~q ),
	.pipe_29_0(\input_if_inst|cmd_queue_inst|pipe[0][29]~q ),
	.pipe_28_0(\input_if_inst|cmd_queue_inst|pipe[0][28]~q ),
	.pipe_33_0(\input_if_inst|cmd_queue_inst|pipe[0][33]~q ),
	.pipe_12_4(\input_if_inst|cmd_queue_inst|pipe[4][12]~q ),
	.pipe_11_4(\input_if_inst|cmd_queue_inst|pipe[4][11]~q ),
	.pipe_10_4(\input_if_inst|cmd_queue_inst|pipe[4][10]~q ),
	.pipe_25_5(\input_if_inst|cmd_queue_inst|pipe[5][25]~q ),
	.pipe_25_0(\input_if_inst|cmd_queue_inst|pipe[0][25]~q ),
	.pipe_26_5(\input_if_inst|cmd_queue_inst|pipe[5][26]~q ),
	.pipe_26_0(\input_if_inst|cmd_queue_inst|pipe[0][26]~q ),
	.pipe_24_5(\input_if_inst|cmd_queue_inst|pipe[5][24]~q ),
	.pipe_24_0(\input_if_inst|cmd_queue_inst|pipe[0][24]~q ),
	.pipe_22_5(\input_if_inst|cmd_queue_inst|pipe[5][22]~q ),
	.pipe_22_0(\input_if_inst|cmd_queue_inst|pipe[0][22]~q ),
	.pipe_23_5(\input_if_inst|cmd_queue_inst|pipe[5][23]~q ),
	.pipe_23_0(\input_if_inst|cmd_queue_inst|pipe[0][23]~q ),
	.pipe_21_5(\input_if_inst|cmd_queue_inst|pipe[5][21]~q ),
	.pipe_21_0(\input_if_inst|cmd_queue_inst|pipe[0][21]~q ),
	.pipe_19_5(\input_if_inst|cmd_queue_inst|pipe[5][19]~q ),
	.pipe_19_0(\input_if_inst|cmd_queue_inst|pipe[0][19]~q ),
	.pipe_20_5(\input_if_inst|cmd_queue_inst|pipe[5][20]~q ),
	.pipe_20_0(\input_if_inst|cmd_queue_inst|pipe[0][20]~q ),
	.pipe_15_5(\input_if_inst|cmd_queue_inst|pipe[5][15]~q ),
	.pipe_15_0(\input_if_inst|cmd_queue_inst|pipe[0][15]~q ),
	.pipe_13_5(\input_if_inst|cmd_queue_inst|pipe[5][13]~q ),
	.pipe_13_0(\input_if_inst|cmd_queue_inst|pipe[0][13]~q ),
	.pipe_14_5(\input_if_inst|cmd_queue_inst|pipe[5][14]~q ),
	.pipe_14_0(\input_if_inst|cmd_queue_inst|pipe[0][14]~q ),
	.pipe_18_5(\input_if_inst|cmd_queue_inst|pipe[5][18]~q ),
	.pipe_18_0(\input_if_inst|cmd_queue_inst|pipe[0][18]~q ),
	.pipe_16_5(\input_if_inst|cmd_queue_inst|pipe[5][16]~q ),
	.pipe_16_0(\input_if_inst|cmd_queue_inst|pipe[0][16]~q ),
	.pipe_17_5(\input_if_inst|cmd_queue_inst|pipe[5][17]~q ),
	.pipe_17_0(\input_if_inst|cmd_queue_inst|pipe[0][17]~q ),
	.pipe_12_5(\input_if_inst|cmd_queue_inst|pipe[5][12]~q ),
	.pipe_11_5(\input_if_inst|cmd_queue_inst|pipe[5][11]~q ),
	.pipe_10_5(\input_if_inst|cmd_queue_inst|pipe[5][10]~q ),
	.pipe_25_3(\input_if_inst|cmd_queue_inst|pipe[3][25]~q ),
	.pipe_26_3(\input_if_inst|cmd_queue_inst|pipe[3][26]~q ),
	.pipe_24_3(\input_if_inst|cmd_queue_inst|pipe[3][24]~q ),
	.pipe_22_3(\input_if_inst|cmd_queue_inst|pipe[3][22]~q ),
	.pipe_23_3(\input_if_inst|cmd_queue_inst|pipe[3][23]~q ),
	.pipe_21_3(\input_if_inst|cmd_queue_inst|pipe[3][21]~q ),
	.pipe_19_3(\input_if_inst|cmd_queue_inst|pipe[3][19]~q ),
	.pipe_20_3(\input_if_inst|cmd_queue_inst|pipe[3][20]~q ),
	.pipe_15_3(\input_if_inst|cmd_queue_inst|pipe[3][15]~q ),
	.pipe_13_3(\input_if_inst|cmd_queue_inst|pipe[3][13]~q ),
	.pipe_14_3(\input_if_inst|cmd_queue_inst|pipe[3][14]~q ),
	.pipe_18_3(\input_if_inst|cmd_queue_inst|pipe[3][18]~q ),
	.pipe_16_3(\input_if_inst|cmd_queue_inst|pipe[3][16]~q ),
	.pipe_17_3(\input_if_inst|cmd_queue_inst|pipe[3][17]~q ),
	.pipe_25_4(\input_if_inst|cmd_queue_inst|pipe[4][25]~q ),
	.pipe_26_4(\input_if_inst|cmd_queue_inst|pipe[4][26]~q ),
	.pipe_24_4(\input_if_inst|cmd_queue_inst|pipe[4][24]~q ),
	.pipe_22_4(\input_if_inst|cmd_queue_inst|pipe[4][22]~q ),
	.pipe_23_4(\input_if_inst|cmd_queue_inst|pipe[4][23]~q ),
	.pipe_21_4(\input_if_inst|cmd_queue_inst|pipe[4][21]~q ),
	.pipe_19_4(\input_if_inst|cmd_queue_inst|pipe[4][19]~q ),
	.pipe_20_4(\input_if_inst|cmd_queue_inst|pipe[4][20]~q ),
	.pipe_15_4(\input_if_inst|cmd_queue_inst|pipe[4][15]~q ),
	.pipe_13_4(\input_if_inst|cmd_queue_inst|pipe[4][13]~q ),
	.pipe_14_4(\input_if_inst|cmd_queue_inst|pipe[4][14]~q ),
	.pipe_18_4(\input_if_inst|cmd_queue_inst|pipe[4][18]~q ),
	.pipe_16_4(\input_if_inst|cmd_queue_inst|pipe[4][16]~q ),
	.pipe_17_4(\input_if_inst|cmd_queue_inst|pipe[4][17]~q ),
	.pipe_12_6(\input_if_inst|cmd_queue_inst|pipe[6][12]~q ),
	.pipe_11_6(\input_if_inst|cmd_queue_inst|pipe[6][11]~q ),
	.pipe_10_6(\input_if_inst|cmd_queue_inst|pipe[6][10]~q ),
	.pipe_25_6(\input_if_inst|cmd_queue_inst|pipe[6][25]~q ),
	.pipe_26_6(\input_if_inst|cmd_queue_inst|pipe[6][26]~q ),
	.pipe_24_6(\input_if_inst|cmd_queue_inst|pipe[6][24]~q ),
	.pipe_22_6(\input_if_inst|cmd_queue_inst|pipe[6][22]~q ),
	.pipe_23_6(\input_if_inst|cmd_queue_inst|pipe[6][23]~q ),
	.pipe_21_6(\input_if_inst|cmd_queue_inst|pipe[6][21]~q ),
	.pipe_19_6(\input_if_inst|cmd_queue_inst|pipe[6][19]~q ),
	.pipe_20_6(\input_if_inst|cmd_queue_inst|pipe[6][20]~q ),
	.pipe_15_6(\input_if_inst|cmd_queue_inst|pipe[6][15]~q ),
	.pipe_13_6(\input_if_inst|cmd_queue_inst|pipe[6][13]~q ),
	.pipe_14_6(\input_if_inst|cmd_queue_inst|pipe[6][14]~q ),
	.pipe_18_6(\input_if_inst|cmd_queue_inst|pipe[6][18]~q ),
	.pipe_16_6(\input_if_inst|cmd_queue_inst|pipe[6][16]~q ),
	.pipe_17_6(\input_if_inst|cmd_queue_inst|pipe[6][17]~q ),
	.pipe_26_7(\input_if_inst|cmd_queue_inst|pipe[7][26]~q ),
	.pipe_24_7(\input_if_inst|cmd_queue_inst|pipe[7][24]~q ),
	.pipe_25_7(\input_if_inst|cmd_queue_inst|pipe[7][25]~q ),
	.pipe_23_7(\input_if_inst|cmd_queue_inst|pipe[7][23]~q ),
	.pipe_21_7(\input_if_inst|cmd_queue_inst|pipe[7][21]~q ),
	.pipe_22_7(\input_if_inst|cmd_queue_inst|pipe[7][22]~q ),
	.pipe_20_7(\input_if_inst|cmd_queue_inst|pipe[7][20]~q ),
	.pipe_18_7(\input_if_inst|cmd_queue_inst|pipe[7][18]~q ),
	.pipe_19_7(\input_if_inst|cmd_queue_inst|pipe[7][19]~q ),
	.pipe_17_7(\input_if_inst|cmd_queue_inst|pipe[7][17]~q ),
	.pipe_15_7(\input_if_inst|cmd_queue_inst|pipe[7][15]~q ),
	.pipe_16_7(\input_if_inst|cmd_queue_inst|pipe[7][16]~q ),
	.pipe_11_7(\input_if_inst|cmd_queue_inst|pipe[7][11]~q ),
	.pipe_10_7(\input_if_inst|cmd_queue_inst|pipe[7][10]~q ),
	.pipe_14_7(\input_if_inst|cmd_queue_inst|pipe[7][14]~q ),
	.pipe_12_7(\input_if_inst|cmd_queue_inst|pipe[7][12]~q ),
	.pipe_13_7(\input_if_inst|cmd_queue_inst|pipe[7][13]~q ),
	.pipe_25_2(\input_if_inst|cmd_queue_inst|pipe[2][25]~q ),
	.pipe_26_2(\input_if_inst|cmd_queue_inst|pipe[2][26]~q ),
	.pipe_24_2(\input_if_inst|cmd_queue_inst|pipe[2][24]~q ),
	.pipe_22_2(\input_if_inst|cmd_queue_inst|pipe[2][22]~q ),
	.pipe_23_2(\input_if_inst|cmd_queue_inst|pipe[2][23]~q ),
	.pipe_21_2(\input_if_inst|cmd_queue_inst|pipe[2][21]~q ),
	.pipe_19_2(\input_if_inst|cmd_queue_inst|pipe[2][19]~q ),
	.pipe_20_2(\input_if_inst|cmd_queue_inst|pipe[2][20]~q ),
	.pipe_15_2(\input_if_inst|cmd_queue_inst|pipe[2][15]~q ),
	.pipe_13_2(\input_if_inst|cmd_queue_inst|pipe[2][13]~q ),
	.pipe_14_2(\input_if_inst|cmd_queue_inst|pipe[2][14]~q ),
	.pipe_18_2(\input_if_inst|cmd_queue_inst|pipe[2][18]~q ),
	.pipe_16_2(\input_if_inst|cmd_queue_inst|pipe[2][16]~q ),
	.pipe_17_2(\input_if_inst|cmd_queue_inst|pipe[2][17]~q ),
	.pipe_25_1(\input_if_inst|cmd_queue_inst|pipe[1][25]~q ),
	.pipe_26_1(\input_if_inst|cmd_queue_inst|pipe[1][26]~q ),
	.pipe_24_1(\input_if_inst|cmd_queue_inst|pipe[1][24]~q ),
	.pipe_22_1(\input_if_inst|cmd_queue_inst|pipe[1][22]~q ),
	.pipe_23_1(\input_if_inst|cmd_queue_inst|pipe[1][23]~q ),
	.pipe_21_1(\input_if_inst|cmd_queue_inst|pipe[1][21]~q ),
	.pipe_19_1(\input_if_inst|cmd_queue_inst|pipe[1][19]~q ),
	.pipe_20_1(\input_if_inst|cmd_queue_inst|pipe[1][20]~q ),
	.pipe_15_1(\input_if_inst|cmd_queue_inst|pipe[1][15]~q ),
	.pipe_13_1(\input_if_inst|cmd_queue_inst|pipe[1][13]~q ),
	.pipe_14_1(\input_if_inst|cmd_queue_inst|pipe[1][14]~q ),
	.pipe_18_1(\input_if_inst|cmd_queue_inst|pipe[1][18]~q ),
	.pipe_16_1(\input_if_inst|cmd_queue_inst|pipe[1][16]~q ),
	.pipe_17_1(\input_if_inst|cmd_queue_inst|pipe[1][17]~q ),
	.pipe_2_0(\input_if_inst|cmd_queue_inst|pipe[0][2]~q ),
	.q_b_132(\input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[132] ),
	.q_b_140(\input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[140] ),
	.q_b_128(\input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[128] ),
	.q_b_136(\input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[136] ),
	.q_b_133(\input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[133] ),
	.q_b_141(\input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[141] ),
	.q_b_129(\input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[129] ),
	.q_b_137(\input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[137] ),
	.q_b_134(\input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[134] ),
	.q_b_142(\input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[142] ),
	.q_b_130(\input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[130] ),
	.q_b_138(\input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[138] ),
	.q_b_135(\input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[135] ),
	.q_b_143(\input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[143] ),
	.q_b_131(\input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[131] ),
	.q_b_139(\input_if_inst|wdata_fifo_inst|wdata_fifo|auto_generated|dpfifo|FIFOram|q_b[139] ),
	.q_b_96(q_b_96),
	.q_b_32(q_b_32),
	.q_b_64(q_b_64),
	.q_b_0(q_b_0),
	.q_b_97(q_b_97),
	.q_b_33(q_b_33),
	.q_b_65(q_b_65),
	.q_b_1(q_b_1),
	.q_b_98(q_b_98),
	.q_b_34(q_b_34),
	.q_b_66(q_b_66),
	.q_b_2(q_b_2),
	.q_b_99(q_b_99),
	.q_b_35(q_b_35),
	.q_b_67(q_b_67),
	.q_b_3(q_b_3),
	.q_b_100(q_b_100),
	.q_b_36(q_b_36),
	.q_b_68(q_b_68),
	.q_b_4(q_b_4),
	.q_b_101(q_b_101),
	.q_b_37(q_b_37),
	.q_b_69(q_b_69),
	.q_b_5(q_b_5),
	.q_b_102(q_b_102),
	.q_b_38(q_b_38),
	.q_b_70(q_b_70),
	.q_b_6(q_b_6),
	.q_b_103(q_b_103),
	.q_b_39(q_b_39),
	.q_b_71(q_b_71),
	.q_b_7(q_b_7),
	.q_b_104(q_b_104),
	.q_b_40(q_b_40),
	.q_b_72(q_b_72),
	.q_b_8(q_b_8),
	.q_b_105(q_b_105),
	.q_b_41(q_b_41),
	.q_b_73(q_b_73),
	.q_b_9(q_b_9),
	.q_b_106(q_b_106),
	.q_b_42(q_b_42),
	.q_b_74(q_b_74),
	.q_b_10(q_b_10),
	.q_b_107(q_b_107),
	.q_b_43(q_b_43),
	.q_b_75(q_b_75),
	.q_b_11(q_b_11),
	.q_b_108(q_b_108),
	.q_b_44(q_b_44),
	.q_b_76(q_b_76),
	.q_b_12(q_b_12),
	.q_b_109(q_b_109),
	.q_b_45(q_b_45),
	.q_b_77(q_b_77),
	.q_b_13(q_b_13),
	.q_b_110(q_b_110),
	.q_b_46(q_b_46),
	.q_b_78(q_b_78),
	.q_b_14(q_b_14),
	.q_b_111(q_b_111),
	.q_b_47(q_b_47),
	.q_b_79(q_b_79),
	.q_b_15(q_b_15),
	.q_b_112(q_b_112),
	.q_b_48(q_b_48),
	.q_b_80(q_b_80),
	.q_b_16(q_b_16),
	.q_b_113(q_b_113),
	.q_b_49(q_b_49),
	.q_b_81(q_b_81),
	.q_b_17(q_b_17),
	.q_b_114(q_b_114),
	.q_b_50(q_b_50),
	.q_b_82(q_b_82),
	.q_b_18(q_b_18),
	.q_b_115(q_b_115),
	.q_b_51(q_b_51),
	.q_b_83(q_b_83),
	.q_b_19(q_b_19),
	.q_b_116(q_b_116),
	.q_b_52(q_b_52),
	.q_b_84(q_b_84),
	.q_b_20(q_b_20),
	.q_b_117(q_b_117),
	.q_b_53(q_b_53),
	.q_b_85(q_b_85),
	.q_b_21(q_b_21),
	.q_b_118(q_b_118),
	.q_b_54(q_b_54),
	.q_b_86(q_b_86),
	.q_b_22(q_b_22),
	.q_b_119(q_b_119),
	.q_b_55(q_b_55),
	.q_b_87(q_b_87),
	.q_b_23(q_b_23),
	.q_b_120(q_b_120),
	.q_b_56(q_b_56),
	.q_b_88(q_b_88),
	.q_b_24(q_b_24),
	.q_b_121(q_b_121),
	.q_b_57(q_b_57),
	.q_b_89(q_b_89),
	.q_b_25(q_b_25),
	.q_b_122(q_b_122),
	.q_b_58(q_b_58),
	.q_b_90(q_b_90),
	.q_b_26(q_b_26),
	.q_b_123(q_b_123),
	.q_b_59(q_b_59),
	.q_b_91(q_b_91),
	.q_b_27(q_b_27),
	.q_b_124(q_b_124),
	.q_b_60(q_b_60),
	.q_b_92(q_b_92),
	.q_b_28(q_b_28),
	.q_b_125(q_b_125),
	.q_b_61(q_b_61),
	.q_b_93(q_b_93),
	.q_b_29(q_b_29),
	.q_b_126(q_b_126),
	.q_b_62(q_b_62),
	.q_b_94(q_b_94),
	.q_b_30(q_b_30),
	.q_b_127(q_b_127),
	.q_b_63(q_b_63),
	.q_b_95(q_b_95),
	.q_b_31(q_b_31),
	.pipe_3_0(\input_if_inst|cmd_queue_inst|pipe[0][3]~q ),
	.pipe_4_0(\input_if_inst|cmd_queue_inst|pipe[0][4]~q ),
	.pipe_5_0(\input_if_inst|cmd_queue_inst|pipe[0][5]~q ),
	.pipe_6_0(\input_if_inst|cmd_queue_inst|pipe[0][6]~q ),
	.pipe_7_0(\input_if_inst|cmd_queue_inst|pipe[0][7]~q ),
	.pipe_8_0(\input_if_inst|cmd_queue_inst|pipe[0][8]~q ),
	.pipe_9_0(\input_if_inst|cmd_queue_inst|pipe[0][9]~q ),
	.hold_ready(\input_if_inst|cmd_gen_inst|hold_ready~q ),
	.pipefull_7(\input_if_inst|cmd_queue_inst|pipefull[7]~q ),
	.ready_out(ready_out),
	.ctl_init_fail(ctl_init_fail),
	.ctl_init_success(ctl_init_success),
	.local_init_done1(local_init_done),
	.internal_ready(\input_if_inst|internal_ready~0_combout ),
	.avalon_write_req(\input_if_inst|avalon_if_inst|avalon_write_req~combout ),
	.reset_reg_4(\clock_and_reset_inst|reset_sync_inst|reset_reg[4]~q ),
	.fetch(\state_machine_inst|fetch~q ),
	.read_req(\input_if_inst|cmd_gen_inst|read_req~0_combout ),
	.write_req(\input_if_inst|cmd_gen_inst|write_req~1_combout ),
	.pipefull_6(\input_if_inst|cmd_queue_inst|pipefull[6]~q ),
	.reset_reg_5(\clock_and_reset_inst|reset_sync_inst|reset_reg[5]~q ),
	.ctl_reset_n({\clock_and_reset_inst|reset_sync_inst|reset_reg[7]~q ,gnd,gnd,gnd,gnd}),
	.ecc_wdata_fifo_read(\afi_block_inst|ecc_wdata_fifo_read~q ),
	.reset_reg_3(\clock_and_reset_inst|reset_sync_inst|reset_reg[3]~q ),
	.always38(\state_machine_inst|always38~0_combout ),
	.pipefull_0(\input_if_inst|cmd_queue_inst|pipefull[0]~q ),
	.pipefull_5(\input_if_inst|cmd_queue_inst|pipefull[5]~q ),
	.pipefull_1(\input_if_inst|cmd_queue_inst|pipefull[1]~q ),
	.pipefull_4(\input_if_inst|cmd_queue_inst|pipefull[4]~q ),
	.pipefull_2(\input_if_inst|cmd_queue_inst|pipefull[2]~q ),
	.pipefull_3(\input_if_inst|cmd_queue_inst|pipefull[3]~q ),
	.GND_port(GND_port),
	.local_size_1(local_size_1),
	.local_address_0(local_address_0),
	.local_size_0(local_size_0),
	.local_size_6(local_size_6),
	.local_size_5(local_size_5),
	.local_size_4(local_size_4),
	.local_size_2(local_size_2),
	.local_size_3(local_size_3),
	.local_read_req(local_read_req),
	.local_write_req(local_write_req),
	.local_burstbegin(local_burstbegin),
	.local_address_8(local_address_8),
	.local_address_10(local_address_10),
	.local_address_9(local_address_9),
	.local_address_23(local_address_23),
	.local_address_24(local_address_24),
	.local_address_22(local_address_22),
	.local_address_20(local_address_20),
	.local_address_21(local_address_21),
	.local_address_19(local_address_19),
	.local_address_17(local_address_17),
	.local_address_18(local_address_18),
	.local_address_13(local_address_13),
	.local_address_11(local_address_11),
	.local_address_12(local_address_12),
	.local_address_16(local_address_16),
	.local_address_14(local_address_14),
	.local_address_15(local_address_15),
	.local_address_1(local_address_1),
	.local_address_2(local_address_2),
	.local_address_3(local_address_3),
	.local_address_4(local_address_4),
	.local_address_5(local_address_5),
	.local_address_7(local_address_7),
	.local_address_6(local_address_6),
	.local_be_4(local_be_4),
	.local_be_12(local_be_12),
	.local_be_0(local_be_0),
	.local_be_8(local_be_8),
	.local_be_5(local_be_5),
	.local_be_13(local_be_13),
	.local_be_1(local_be_1),
	.local_be_9(local_be_9),
	.local_be_6(local_be_6),
	.local_be_14(local_be_14),
	.local_be_2(local_be_2),
	.local_be_10(local_be_10),
	.local_be_7(local_be_7),
	.local_be_15(local_be_15),
	.local_be_3(local_be_3),
	.local_be_11(local_be_11),
	.local_wdata_96(local_wdata_96),
	.local_wdata_32(local_wdata_32),
	.local_wdata_64(local_wdata_64),
	.local_wdata_0(local_wdata_0),
	.local_wdata_97(local_wdata_97),
	.local_wdata_33(local_wdata_33),
	.local_wdata_65(local_wdata_65),
	.local_wdata_1(local_wdata_1),
	.local_wdata_98(local_wdata_98),
	.local_wdata_34(local_wdata_34),
	.local_wdata_66(local_wdata_66),
	.local_wdata_2(local_wdata_2),
	.local_wdata_99(local_wdata_99),
	.local_wdata_35(local_wdata_35),
	.local_wdata_67(local_wdata_67),
	.local_wdata_3(local_wdata_3),
	.local_wdata_100(local_wdata_100),
	.local_wdata_36(local_wdata_36),
	.local_wdata_68(local_wdata_68),
	.local_wdata_4(local_wdata_4),
	.local_wdata_101(local_wdata_101),
	.local_wdata_37(local_wdata_37),
	.local_wdata_69(local_wdata_69),
	.local_wdata_5(local_wdata_5),
	.local_wdata_102(local_wdata_102),
	.local_wdata_38(local_wdata_38),
	.local_wdata_70(local_wdata_70),
	.local_wdata_6(local_wdata_6),
	.local_wdata_103(local_wdata_103),
	.local_wdata_39(local_wdata_39),
	.local_wdata_71(local_wdata_71),
	.local_wdata_7(local_wdata_7),
	.local_wdata_104(local_wdata_104),
	.local_wdata_40(local_wdata_40),
	.local_wdata_72(local_wdata_72),
	.local_wdata_8(local_wdata_8),
	.local_wdata_105(local_wdata_105),
	.local_wdata_41(local_wdata_41),
	.local_wdata_73(local_wdata_73),
	.local_wdata_9(local_wdata_9),
	.local_wdata_106(local_wdata_106),
	.local_wdata_42(local_wdata_42),
	.local_wdata_74(local_wdata_74),
	.local_wdata_10(local_wdata_10),
	.local_wdata_107(local_wdata_107),
	.local_wdata_43(local_wdata_43),
	.local_wdata_75(local_wdata_75),
	.local_wdata_11(local_wdata_11),
	.local_wdata_108(local_wdata_108),
	.local_wdata_44(local_wdata_44),
	.local_wdata_76(local_wdata_76),
	.local_wdata_12(local_wdata_12),
	.local_wdata_109(local_wdata_109),
	.local_wdata_45(local_wdata_45),
	.local_wdata_77(local_wdata_77),
	.local_wdata_13(local_wdata_13),
	.local_wdata_110(local_wdata_110),
	.local_wdata_46(local_wdata_46),
	.local_wdata_78(local_wdata_78),
	.local_wdata_14(local_wdata_14),
	.local_wdata_111(local_wdata_111),
	.local_wdata_47(local_wdata_47),
	.local_wdata_79(local_wdata_79),
	.local_wdata_15(local_wdata_15),
	.local_wdata_112(local_wdata_112),
	.local_wdata_48(local_wdata_48),
	.local_wdata_80(local_wdata_80),
	.local_wdata_16(local_wdata_16),
	.local_wdata_113(local_wdata_113),
	.local_wdata_49(local_wdata_49),
	.local_wdata_81(local_wdata_81),
	.local_wdata_17(local_wdata_17),
	.local_wdata_114(local_wdata_114),
	.local_wdata_50(local_wdata_50),
	.local_wdata_82(local_wdata_82),
	.local_wdata_18(local_wdata_18),
	.local_wdata_115(local_wdata_115),
	.local_wdata_51(local_wdata_51),
	.local_wdata_83(local_wdata_83),
	.local_wdata_19(local_wdata_19),
	.local_wdata_116(local_wdata_116),
	.local_wdata_52(local_wdata_52),
	.local_wdata_84(local_wdata_84),
	.local_wdata_20(local_wdata_20),
	.local_wdata_117(local_wdata_117),
	.local_wdata_53(local_wdata_53),
	.local_wdata_85(local_wdata_85),
	.local_wdata_21(local_wdata_21),
	.local_wdata_118(local_wdata_118),
	.local_wdata_54(local_wdata_54),
	.local_wdata_86(local_wdata_86),
	.local_wdata_22(local_wdata_22),
	.local_wdata_119(local_wdata_119),
	.local_wdata_55(local_wdata_55),
	.local_wdata_87(local_wdata_87),
	.local_wdata_23(local_wdata_23),
	.local_wdata_120(local_wdata_120),
	.local_wdata_56(local_wdata_56),
	.local_wdata_88(local_wdata_88),
	.local_wdata_24(local_wdata_24),
	.local_wdata_121(local_wdata_121),
	.local_wdata_57(local_wdata_57),
	.local_wdata_89(local_wdata_89),
	.local_wdata_25(local_wdata_25),
	.local_wdata_122(local_wdata_122),
	.local_wdata_58(local_wdata_58),
	.local_wdata_90(local_wdata_90),
	.local_wdata_26(local_wdata_26),
	.local_wdata_123(local_wdata_123),
	.local_wdata_59(local_wdata_59),
	.local_wdata_91(local_wdata_91),
	.local_wdata_27(local_wdata_27),
	.local_wdata_124(local_wdata_124),
	.local_wdata_60(local_wdata_60),
	.local_wdata_92(local_wdata_92),
	.local_wdata_28(local_wdata_28),
	.local_wdata_125(local_wdata_125),
	.local_wdata_61(local_wdata_61),
	.local_wdata_93(local_wdata_93),
	.local_wdata_29(local_wdata_29),
	.local_wdata_126(local_wdata_126),
	.local_wdata_62(local_wdata_62),
	.local_wdata_94(local_wdata_94),
	.local_wdata_30(local_wdata_30),
	.local_wdata_127(local_wdata_127),
	.local_wdata_63(local_wdata_63),
	.local_wdata_95(local_wdata_95),
	.local_wdata_31(local_wdata_31));

endmodule

module ddr3_int_alt_ddrx_addr_cmd (
	ctl_clk,
	do_read_r,
	do_auto_precharge_r,
	do_write_r,
	do_burst_chop_r,
	to_row_addr_r_0,
	to_row_addr_r_1,
	to_col_addr_r_2,
	to_row_addr_r_2,
	to_col_addr_r_3,
	to_row_addr_r_3,
	to_col_addr_r_4,
	to_row_addr_r_4,
	to_col_addr_r_5,
	to_row_addr_r_5,
	to_col_addr_r_6,
	to_row_addr_r_6,
	to_col_addr_r_7,
	to_row_addr_r_7,
	to_col_addr_r_8,
	to_row_addr_r_8,
	to_col_addr_r_9,
	to_row_addr_r_9,
	to_row_addr_r_10,
	to_row_addr_r_11,
	to_row_addr_r_12,
	to_row_addr_r_13,
	ctl_init_success,
	do_precharge_all_r,
	do_refresh_r,
	to_chip_r_0,
	to_bank_addr_r_2,
	to_bank_addr_r_0,
	to_bank_addr_r_1,
	do_activate_r,
	always1,
	afi_cs_n_1,
	int_cke_r_0,
	afi_addr_0,
	afi_addr_1,
	afi_addr_2,
	afi_addr_3,
	afi_addr_4,
	afi_addr_5,
	afi_addr_6,
	afi_addr_7,
	afi_addr_8,
	afi_addr_9,
	afi_addr_10,
	afi_addr_11,
	afi_addr_12,
	afi_addr_13,
	afi_ba_0,
	afi_ba_1,
	afi_ba_2,
	afi_ras_n_0,
	afi_cas_n_0,
	afi_we_n_0,
	ctl_reset_n)/* synthesis synthesis_greybox=0 */;
input 	ctl_clk;
input 	do_read_r;
input 	do_auto_precharge_r;
input 	do_write_r;
input 	do_burst_chop_r;
input 	to_row_addr_r_0;
input 	to_row_addr_r_1;
input 	to_col_addr_r_2;
input 	to_row_addr_r_2;
input 	to_col_addr_r_3;
input 	to_row_addr_r_3;
input 	to_col_addr_r_4;
input 	to_row_addr_r_4;
input 	to_col_addr_r_5;
input 	to_row_addr_r_5;
input 	to_col_addr_r_6;
input 	to_row_addr_r_6;
input 	to_col_addr_r_7;
input 	to_row_addr_r_7;
input 	to_col_addr_r_8;
input 	to_row_addr_r_8;
input 	to_col_addr_r_9;
input 	to_row_addr_r_9;
input 	to_row_addr_r_10;
input 	to_row_addr_r_11;
input 	to_row_addr_r_12;
input 	to_row_addr_r_13;
input 	ctl_init_success;
input 	do_precharge_all_r;
input 	do_refresh_r;
input 	to_chip_r_0;
input 	to_bank_addr_r_2;
input 	to_bank_addr_r_0;
input 	to_bank_addr_r_1;
input 	do_activate_r;
input 	always1;
output 	afi_cs_n_1;
output 	int_cke_r_0;
output 	afi_addr_0;
output 	afi_addr_1;
output 	afi_addr_2;
output 	afi_addr_3;
output 	afi_addr_4;
output 	afi_addr_5;
output 	afi_addr_6;
output 	afi_addr_7;
output 	afi_addr_8;
output 	afi_addr_9;
output 	afi_addr_10;
output 	afi_addr_11;
output 	afi_addr_12;
output 	afi_addr_13;
output 	afi_ba_0;
output 	afi_ba_1;
output 	afi_ba_2;
output 	afi_ras_n_0;
output 	afi_cas_n_0;
output 	afi_we_n_0;
input 	ctl_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



arriaii_lcell_comb \afi_cs_n[1]~0 (
	.dataa(!ctl_init_success),
	.datab(!do_precharge_all_r),
	.datac(!do_refresh_r),
	.datad(!to_chip_r_0),
	.datae(!do_activate_r),
	.dataf(!always1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_cs_n_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_cs_n[1]~0 .extended_lut = "off";
defparam \afi_cs_n[1]~0 .lut_mask = 64'hFFEAFFAAFFAAFFAA;
defparam \afi_cs_n[1]~0 .shared_arith = "off";

dffeas \int_cke_r[0] (
	.clk(ctl_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(int_cke_r_0),
	.prn(vcc));
defparam \int_cke_r[0] .is_wysiwyg = "true";
defparam \int_cke_r[0] .power_up = "low";

arriaii_lcell_comb \afi_addr[0]~0 (
	.dataa(!ctl_init_success),
	.datab(!do_activate_r),
	.datac(!always1),
	.datad(!to_row_addr_r_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_addr_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_addr[0]~0 .extended_lut = "off";
defparam \afi_addr[0]~0 .lut_mask = 64'h0010001000100010;
defparam \afi_addr[0]~0 .shared_arith = "off";

arriaii_lcell_comb \afi_addr[1]~1 (
	.dataa(!ctl_init_success),
	.datab(!do_activate_r),
	.datac(!always1),
	.datad(!to_row_addr_r_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_addr_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_addr[1]~1 .extended_lut = "off";
defparam \afi_addr[1]~1 .lut_mask = 64'h0010001000100010;
defparam \afi_addr[1]~1 .shared_arith = "off";

arriaii_lcell_comb \afi_addr[2]~2 (
	.dataa(!ctl_init_success),
	.datab(!do_activate_r),
	.datac(!always1),
	.datad(!to_col_addr_r_2),
	.datae(!to_row_addr_r_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_addr_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_addr[2]~2 .extended_lut = "off";
defparam \afi_addr[2]~2 .lut_mask = 64'h0005101500051015;
defparam \afi_addr[2]~2 .shared_arith = "off";

arriaii_lcell_comb \afi_addr[3]~3 (
	.dataa(!ctl_init_success),
	.datab(!do_activate_r),
	.datac(!always1),
	.datad(!to_col_addr_r_3),
	.datae(!to_row_addr_r_3),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_addr_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_addr[3]~3 .extended_lut = "off";
defparam \afi_addr[3]~3 .lut_mask = 64'h0005101500051015;
defparam \afi_addr[3]~3 .shared_arith = "off";

arriaii_lcell_comb \afi_addr[4]~4 (
	.dataa(!ctl_init_success),
	.datab(!do_activate_r),
	.datac(!always1),
	.datad(!to_col_addr_r_4),
	.datae(!to_row_addr_r_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_addr_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_addr[4]~4 .extended_lut = "off";
defparam \afi_addr[4]~4 .lut_mask = 64'h0005101500051015;
defparam \afi_addr[4]~4 .shared_arith = "off";

arriaii_lcell_comb \afi_addr[5]~5 (
	.dataa(!ctl_init_success),
	.datab(!do_activate_r),
	.datac(!always1),
	.datad(!to_col_addr_r_5),
	.datae(!to_row_addr_r_5),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_addr_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_addr[5]~5 .extended_lut = "off";
defparam \afi_addr[5]~5 .lut_mask = 64'h0005101500051015;
defparam \afi_addr[5]~5 .shared_arith = "off";

arriaii_lcell_comb \afi_addr[6]~6 (
	.dataa(!ctl_init_success),
	.datab(!do_activate_r),
	.datac(!always1),
	.datad(!to_col_addr_r_6),
	.datae(!to_row_addr_r_6),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_addr_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_addr[6]~6 .extended_lut = "off";
defparam \afi_addr[6]~6 .lut_mask = 64'h0005101500051015;
defparam \afi_addr[6]~6 .shared_arith = "off";

arriaii_lcell_comb \afi_addr[7]~7 (
	.dataa(!ctl_init_success),
	.datab(!do_activate_r),
	.datac(!always1),
	.datad(!to_col_addr_r_7),
	.datae(!to_row_addr_r_7),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_addr_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_addr[7]~7 .extended_lut = "off";
defparam \afi_addr[7]~7 .lut_mask = 64'h0005101500051015;
defparam \afi_addr[7]~7 .shared_arith = "off";

arriaii_lcell_comb \afi_addr[8]~8 (
	.dataa(!ctl_init_success),
	.datab(!do_activate_r),
	.datac(!always1),
	.datad(!to_col_addr_r_8),
	.datae(!to_row_addr_r_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_addr_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_addr[8]~8 .extended_lut = "off";
defparam \afi_addr[8]~8 .lut_mask = 64'h0005101500051015;
defparam \afi_addr[8]~8 .shared_arith = "off";

arriaii_lcell_comb \afi_addr[9]~9 (
	.dataa(!ctl_init_success),
	.datab(!do_activate_r),
	.datac(!always1),
	.datad(!to_col_addr_r_9),
	.datae(!to_row_addr_r_9),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_addr_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_addr[9]~9 .extended_lut = "off";
defparam \afi_addr[9]~9 .lut_mask = 64'h0005101500051015;
defparam \afi_addr[9]~9 .shared_arith = "off";

arriaii_lcell_comb \afi_addr[10]~10 (
	.dataa(!ctl_init_success),
	.datab(!do_precharge_all_r),
	.datac(!do_auto_precharge_r),
	.datad(!do_activate_r),
	.datae(!always1),
	.dataf(!to_row_addr_r_10),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_addr_10),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_addr[10]~10 .extended_lut = "off";
defparam \afi_addr[10]~10 .lut_mask = 64'h1100050511550505;
defparam \afi_addr[10]~10 .shared_arith = "off";

arriaii_lcell_comb \afi_addr[11]~11 (
	.dataa(!ctl_init_success),
	.datab(!do_activate_r),
	.datac(!always1),
	.datad(!to_row_addr_r_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_addr_11),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_addr[11]~11 .extended_lut = "off";
defparam \afi_addr[11]~11 .lut_mask = 64'h0010001000100010;
defparam \afi_addr[11]~11 .shared_arith = "off";

arriaii_lcell_comb \afi_addr[12]~12 (
	.dataa(!ctl_init_success),
	.datab(!do_activate_r),
	.datac(!do_burst_chop_r),
	.datad(!always1),
	.datae(!to_row_addr_r_12),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_addr_12),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_addr[12]~12 .extended_lut = "off";
defparam \afi_addr[12]~12 .lut_mask = 64'h0050115000501150;
defparam \afi_addr[12]~12 .shared_arith = "off";

arriaii_lcell_comb \afi_addr[13]~13 (
	.dataa(!ctl_init_success),
	.datab(!do_activate_r),
	.datac(!always1),
	.datad(!to_row_addr_r_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_addr_13),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_addr[13]~13 .extended_lut = "off";
defparam \afi_addr[13]~13 .lut_mask = 64'h0010001000100010;
defparam \afi_addr[13]~13 .shared_arith = "off";

arriaii_lcell_comb \afi_ba[0]~0 (
	.dataa(!ctl_init_success),
	.datab(!do_precharge_all_r),
	.datac(!to_bank_addr_r_0),
	.datad(!do_activate_r),
	.datae(!always1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_ba_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_ba[0]~0 .extended_lut = "off";
defparam \afi_ba[0]~0 .lut_mask = 64'h0105050501050505;
defparam \afi_ba[0]~0 .shared_arith = "off";

arriaii_lcell_comb \afi_ba[1]~1 (
	.dataa(!ctl_init_success),
	.datab(!do_precharge_all_r),
	.datac(!to_bank_addr_r_1),
	.datad(!do_activate_r),
	.datae(!always1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_ba_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_ba[1]~1 .extended_lut = "off";
defparam \afi_ba[1]~1 .lut_mask = 64'h0105050501050505;
defparam \afi_ba[1]~1 .shared_arith = "off";

arriaii_lcell_comb \afi_ba[2]~2 (
	.dataa(!ctl_init_success),
	.datab(!do_precharge_all_r),
	.datac(!to_bank_addr_r_2),
	.datad(!do_activate_r),
	.datae(!always1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_ba_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_ba[2]~2 .extended_lut = "off";
defparam \afi_ba[2]~2 .lut_mask = 64'h0105050501050505;
defparam \afi_ba[2]~2 .shared_arith = "off";

arriaii_lcell_comb \afi_ras_n[0]~0 (
	.dataa(!ctl_init_success),
	.datab(!do_precharge_all_r),
	.datac(!do_refresh_r),
	.datad(!do_activate_r),
	.datae(!always1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_ras_n_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_ras_n[0]~0 .extended_lut = "off";
defparam \afi_ras_n[0]~0 .lut_mask = 64'hEAAAFFFFEAAAFFFF;
defparam \afi_ras_n[0]~0 .shared_arith = "off";

arriaii_lcell_comb \afi_cas_n[0]~0 (
	.dataa(!ctl_init_success),
	.datab(!do_precharge_all_r),
	.datac(!do_refresh_r),
	.datad(!do_activate_r),
	.datae(!always1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_cas_n_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_cas_n[0]~0 .extended_lut = "off";
defparam \afi_cas_n[0]~0 .lut_mask = 64'hFBFFAAAAFBFFAAAA;
defparam \afi_cas_n[0]~0 .shared_arith = "off";

arriaii_lcell_comb \afi_we_n[0]~0 (
	.dataa(!ctl_init_success),
	.datab(!do_precharge_all_r),
	.datac(!do_read_r),
	.datad(!do_write_r),
	.datae(!do_activate_r),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_we_n_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_we_n[0]~0 .extended_lut = "off";
defparam \afi_we_n[0]~0 .lut_mask = 64'hEFAFFFAFEFAFFFAF;
defparam \afi_we_n[0]~0 .shared_arith = "off";

endmodule

module ddr3_int_alt_ddrx_afi_block (
	ctl_clk,
	do_read_r,
	do_write_r,
	do_burst_chop_r,
	q_b_132,
	q_b_140,
	q_b_128,
	q_b_136,
	q_b_133,
	q_b_141,
	q_b_129,
	q_b_137,
	q_b_134,
	q_b_142,
	q_b_130,
	q_b_138,
	q_b_135,
	q_b_143,
	q_b_131,
	q_b_139,
	ecc_wdata_fifo_read1,
	rdwr_data_valid,
	ctl_reset_n,
	doing_read1,
	wd_lat_2,
	afi_wlat,
	wd_lat_0,
	afi_dm_4,
	afi_dm_12,
	afi_dm_0,
	afi_dm_8,
	afi_dm_5,
	afi_dm_13,
	afi_dm_1,
	afi_dm_9,
	afi_dm_6,
	afi_dm_14,
	afi_dm_2,
	afi_dm_10,
	afi_dm_7,
	afi_dm_15,
	afi_dm_3,
	afi_dm_11,
	int_wdata_valid1,
	int_dqs_burst1,
	int_dqs_burst_hr1)/* synthesis synthesis_greybox=0 */;
input 	ctl_clk;
input 	do_read_r;
input 	do_write_r;
input 	do_burst_chop_r;
input 	q_b_132;
input 	q_b_140;
input 	q_b_128;
input 	q_b_136;
input 	q_b_133;
input 	q_b_141;
input 	q_b_129;
input 	q_b_137;
input 	q_b_134;
input 	q_b_142;
input 	q_b_130;
input 	q_b_138;
input 	q_b_135;
input 	q_b_143;
input 	q_b_131;
input 	q_b_139;
output 	ecc_wdata_fifo_read1;
input 	rdwr_data_valid;
input 	ctl_reset_n;
output 	doing_read1;
input 	wd_lat_2;
input 	[4:0] afi_wlat;
input 	wd_lat_0;
output 	afi_dm_4;
output 	afi_dm_12;
output 	afi_dm_0;
output 	afi_dm_8;
output 	afi_dm_5;
output 	afi_dm_13;
output 	afi_dm_1;
output 	afi_dm_9;
output 	afi_dm_6;
output 	afi_dm_14;
output 	afi_dm_2;
output 	afi_dm_10;
output 	afi_dm_7;
output 	afi_dm_15;
output 	afi_dm_3;
output 	afi_dm_11;
output 	int_wdata_valid1;
output 	int_dqs_burst1;
output 	int_dqs_burst_hr1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Mux0~0_combout ;
wire \Mux0~4_combout ;
wire \rdwr_data_valid_pipe[31]~q ;
wire \rdwr_data_valid_pipe[29]~q ;
wire \rdwr_data_valid_pipe[30]~q ;
wire \afi_wlat_r[2]~q ;
wire \rdwr_data_valid_pipe[27]~q ;
wire \rdwr_data_valid_pipe[25]~q ;
wire \rdwr_data_valid_pipe[26]~q ;
wire \rdwr_data_valid_pipe[24]~q ;
wire \rdwr_data_valid_pipe[28]~q ;
wire \rdwr_data_valid_pipe[23]~q ;
wire \doing_write_pipe[25]~q ;
wire \Mux1~0_combout ;
wire \doing_write_pipe[29]~q ;
wire \doing_write_pipe[28]~q ;
wire \Mux1~5_combout ;
wire \doing_write_pipe[27]~q ;
wire \doing_write_pipe[26]~q ;
wire \Mux1~10_combout ;
wire \doing_write_pipe[31]~q ;
wire \doing_write_pipe[30]~q ;
wire \Mux1~15_combout ;
wire \Mux1~21_combout ;
wire \Mux1~25_combout ;
wire \Mux1~29_combout ;
wire \Mux1~33_combout ;
wire \afi_wlat_r[2]~0_combout ;
wire \rdwr_data_valid_pipe[0]~q ;
wire \rdwr_data_valid_pipe[1]~q ;
wire \rdwr_data_valid_pipe[2]~q ;
wire \rdwr_data_valid_pipe[3]~q ;
wire \rdwr_data_valid_pipe[4]~q ;
wire \rdwr_data_valid_pipe[5]~q ;
wire \rdwr_data_valid_pipe[6]~q ;
wire \rdwr_data_valid_pipe[7]~q ;
wire \rdwr_data_valid_pipe[8]~q ;
wire \rdwr_data_valid_pipe[9]~q ;
wire \rdwr_data_valid_pipe[10]~q ;
wire \rdwr_data_valid_pipe[11]~q ;
wire \rdwr_data_valid_pipe[12]~q ;
wire \rdwr_data_valid_pipe[13]~q ;
wire \rdwr_data_valid_pipe[14]~q ;
wire \rdwr_data_valid_pipe[15]~q ;
wire \rdwr_data_valid_pipe[16]~q ;
wire \rdwr_data_valid_pipe[17]~q ;
wire \rdwr_data_valid_pipe[18]~q ;
wire \rdwr_data_valid_pipe[19]~q ;
wire \rdwr_data_valid_pipe[20]~q ;
wire \rdwr_data_valid_pipe[21]~q ;
wire \afi_wlat_r[1]~q ;
wire \Add0~0_combout ;
wire \afi_wlat_r[0]~1_combout ;
wire \afi_wlat_r[0]~q ;
wire \Mux0~8_combout ;
wire \rdwr_data_valid_pipe[22]~q ;
wire \Mux0~12_combout ;
wire \Mux0~16_combout ;
wire \Mux0~20_combout ;
wire \Mux0~24_combout ;
wire \Mux0~28_combout ;
wire \afi_wlat_r[3]~q ;
wire \Add0~1_combout ;
wire \afi_wlat_r[4]~q ;
wire \Add0~2_combout ;
wire \Mux0~32_combout ;
wire \doing_write~0_combout ;
wire \doing_write~q ;
wire \always8~0_combout ;
wire \doing_write_pipe[0]~q ;
wire \doing_write_pipe[1]~q ;
wire \doing_write_pipe[2]~q ;
wire \doing_write_pipe[3]~q ;
wire \doing_write_pipe[4]~q ;
wire \doing_write_pipe[5]~q ;
wire \doing_write_pipe[6]~q ;
wire \doing_write_pipe[7]~q ;
wire \doing_write_pipe[8]~q ;
wire \doing_write_pipe[9]~q ;
wire \doing_write_pipe[10]~q ;
wire \doing_write_pipe[11]~q ;
wire \doing_write_pipe[12]~q ;
wire \doing_write_pipe[13]~q ;
wire \doing_write_pipe[14]~q ;
wire \doing_write_pipe[15]~q ;
wire \doing_write_pipe[16]~q ;
wire \doing_write_pipe[17]~q ;
wire \Mux1~1_combout ;
wire \Mux1~2_combout ;
wire \Mux1~3_combout ;
wire \Mux1~4_combout ;
wire \doing_write_pipe[18]~q ;
wire \doing_write_pipe[19]~q ;
wire \doing_write_pipe[20]~q ;
wire \doing_write_pipe[21]~q ;
wire \Mux1~6_combout ;
wire \Mux1~7_combout ;
wire \Mux1~8_combout ;
wire \Mux1~9_combout ;
wire \Mux1~11_combout ;
wire \Mux1~12_combout ;
wire \Mux1~13_combout ;
wire \Mux1~14_combout ;
wire \doing_write_pipe[22]~q ;
wire \doing_write_pipe[23]~q ;
wire \Mux1~16_combout ;
wire \Mux1~17_combout ;
wire \Mux1~18_combout ;
wire \Mux1~19_combout ;
wire \Mux1~20_combout ;
wire \Equal0~0_combout ;
wire \ecc_wdata_fifo_read~0_combout ;
wire \doing_read~0_combout ;
wire \int_real_wdata_valid~q ;
wire \Mux1~22_combout ;
wire \Mux1~23_combout ;
wire \Mux1~24_combout ;
wire \Mux3~0_combout ;
wire \Mux1~26_combout ;
wire \Mux1~27_combout ;
wire \Mux1~28_combout ;
wire \Mux3~1_combout ;
wire \Mux1~30_combout ;
wire \Mux1~31_combout ;
wire \Mux1~32_combout ;
wire \Mux3~2_combout ;
wire \doing_write_pipe[24]~q ;
wire \Mux1~34_combout ;
wire \Mux1~35_combout ;
wire \Mux1~36_combout ;
wire \Mux3~3_combout ;
wire \Mux3~4_combout ;
wire \int_wdata_valid~0_combout ;
wire \int_dqs_burst~0_combout ;


arriaii_lcell_comb \Mux0~0 (
	.dataa(!\rdwr_data_valid_pipe[27]~q ),
	.datab(!\rdwr_data_valid_pipe[25]~q ),
	.datac(!\rdwr_data_valid_pipe[24]~q ),
	.datad(!\afi_wlat_r[0]~q ),
	.datae(!\afi_wlat_r[1]~q ),
	.dataf(!\Add0~0_combout ),
	.datag(!\rdwr_data_valid_pipe[26]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~0 .extended_lut = "on";
defparam \Mux0~0 .lut_mask = 64'h0F550F3300FF00FF;
defparam \Mux0~0 .shared_arith = "off";

arriaii_lcell_comb \Mux0~4 (
	.dataa(!\rdwr_data_valid_pipe[31]~q ),
	.datab(!\rdwr_data_valid_pipe[29]~q ),
	.datac(!\rdwr_data_valid_pipe[28]~q ),
	.datad(!\Add0~0_combout ),
	.datae(!\afi_wlat_r[1]~q ),
	.dataf(!\Mux0~0_combout ),
	.datag(!\rdwr_data_valid_pipe[30]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~4 .extended_lut = "on";
defparam \Mux0~4 .lut_mask = 64'h000F000FFF55FF33;
defparam \Mux0~4 .shared_arith = "off";

dffeas \rdwr_data_valid_pipe[31] (
	.clk(ctl_clk),
	.d(\rdwr_data_valid_pipe[30]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_data_valid_pipe[31]~q ),
	.prn(vcc));
defparam \rdwr_data_valid_pipe[31] .is_wysiwyg = "true";
defparam \rdwr_data_valid_pipe[31] .power_up = "low";

dffeas \rdwr_data_valid_pipe[29] (
	.clk(ctl_clk),
	.d(\rdwr_data_valid_pipe[28]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_data_valid_pipe[29]~q ),
	.prn(vcc));
defparam \rdwr_data_valid_pipe[29] .is_wysiwyg = "true";
defparam \rdwr_data_valid_pipe[29] .power_up = "low";

dffeas \rdwr_data_valid_pipe[30] (
	.clk(ctl_clk),
	.d(\rdwr_data_valid_pipe[29]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_data_valid_pipe[30]~q ),
	.prn(vcc));
defparam \rdwr_data_valid_pipe[30] .is_wysiwyg = "true";
defparam \rdwr_data_valid_pipe[30] .power_up = "low";

dffeas \afi_wlat_r[2] (
	.clk(ctl_clk),
	.d(\afi_wlat_r[2]~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\afi_wlat_r[2]~q ),
	.prn(vcc));
defparam \afi_wlat_r[2] .is_wysiwyg = "true";
defparam \afi_wlat_r[2] .power_up = "low";

dffeas \rdwr_data_valid_pipe[27] (
	.clk(ctl_clk),
	.d(\rdwr_data_valid_pipe[26]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_data_valid_pipe[27]~q ),
	.prn(vcc));
defparam \rdwr_data_valid_pipe[27] .is_wysiwyg = "true";
defparam \rdwr_data_valid_pipe[27] .power_up = "low";

dffeas \rdwr_data_valid_pipe[25] (
	.clk(ctl_clk),
	.d(\rdwr_data_valid_pipe[24]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_data_valid_pipe[25]~q ),
	.prn(vcc));
defparam \rdwr_data_valid_pipe[25] .is_wysiwyg = "true";
defparam \rdwr_data_valid_pipe[25] .power_up = "low";

dffeas \rdwr_data_valid_pipe[26] (
	.clk(ctl_clk),
	.d(\rdwr_data_valid_pipe[25]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_data_valid_pipe[26]~q ),
	.prn(vcc));
defparam \rdwr_data_valid_pipe[26] .is_wysiwyg = "true";
defparam \rdwr_data_valid_pipe[26] .power_up = "low";

dffeas \rdwr_data_valid_pipe[24] (
	.clk(ctl_clk),
	.d(\rdwr_data_valid_pipe[23]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_data_valid_pipe[24]~q ),
	.prn(vcc));
defparam \rdwr_data_valid_pipe[24] .is_wysiwyg = "true";
defparam \rdwr_data_valid_pipe[24] .power_up = "low";

dffeas \rdwr_data_valid_pipe[28] (
	.clk(ctl_clk),
	.d(\rdwr_data_valid_pipe[27]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_data_valid_pipe[28]~q ),
	.prn(vcc));
defparam \rdwr_data_valid_pipe[28] .is_wysiwyg = "true";
defparam \rdwr_data_valid_pipe[28] .power_up = "low";

dffeas \rdwr_data_valid_pipe[23] (
	.clk(ctl_clk),
	.d(\rdwr_data_valid_pipe[22]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_data_valid_pipe[23]~q ),
	.prn(vcc));
defparam \rdwr_data_valid_pipe[23] .is_wysiwyg = "true";
defparam \rdwr_data_valid_pipe[23] .power_up = "low";

dffeas \doing_write_pipe[25] (
	.clk(ctl_clk),
	.d(\doing_write_pipe[24]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write_pipe[25]~q ),
	.prn(vcc));
defparam \doing_write_pipe[25] .is_wysiwyg = "true";
defparam \doing_write_pipe[25] .power_up = "low";

arriaii_lcell_comb \Mux1~0 (
	.dataa(!\afi_wlat_r[0]~q ),
	.datab(!\doing_write_pipe[25]~q ),
	.datac(!\doing_write_pipe[24]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~0 .extended_lut = "off";
defparam \Mux1~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \Mux1~0 .shared_arith = "off";

dffeas \doing_write_pipe[29] (
	.clk(ctl_clk),
	.d(\doing_write_pipe[28]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write_pipe[29]~q ),
	.prn(vcc));
defparam \doing_write_pipe[29] .is_wysiwyg = "true";
defparam \doing_write_pipe[29] .power_up = "low";

dffeas \doing_write_pipe[28] (
	.clk(ctl_clk),
	.d(\doing_write_pipe[27]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write_pipe[28]~q ),
	.prn(vcc));
defparam \doing_write_pipe[28] .is_wysiwyg = "true";
defparam \doing_write_pipe[28] .power_up = "low";

arriaii_lcell_comb \Mux1~5 (
	.dataa(!\afi_wlat_r[0]~q ),
	.datab(!\doing_write_pipe[29]~q ),
	.datac(!\doing_write_pipe[28]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~5 .extended_lut = "off";
defparam \Mux1~5 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \Mux1~5 .shared_arith = "off";

dffeas \doing_write_pipe[27] (
	.clk(ctl_clk),
	.d(\doing_write_pipe[26]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write_pipe[27]~q ),
	.prn(vcc));
defparam \doing_write_pipe[27] .is_wysiwyg = "true";
defparam \doing_write_pipe[27] .power_up = "low";

dffeas \doing_write_pipe[26] (
	.clk(ctl_clk),
	.d(\doing_write_pipe[25]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write_pipe[26]~q ),
	.prn(vcc));
defparam \doing_write_pipe[26] .is_wysiwyg = "true";
defparam \doing_write_pipe[26] .power_up = "low";

arriaii_lcell_comb \Mux1~10 (
	.dataa(!\afi_wlat_r[0]~q ),
	.datab(!\doing_write_pipe[27]~q ),
	.datac(!\doing_write_pipe[26]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~10 .extended_lut = "off";
defparam \Mux1~10 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \Mux1~10 .shared_arith = "off";

dffeas \doing_write_pipe[31] (
	.clk(ctl_clk),
	.d(\doing_write_pipe[30]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write_pipe[31]~q ),
	.prn(vcc));
defparam \doing_write_pipe[31] .is_wysiwyg = "true";
defparam \doing_write_pipe[31] .power_up = "low";

dffeas \doing_write_pipe[30] (
	.clk(ctl_clk),
	.d(\doing_write_pipe[29]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write_pipe[30]~q ),
	.prn(vcc));
defparam \doing_write_pipe[30] .is_wysiwyg = "true";
defparam \doing_write_pipe[30] .power_up = "low";

arriaii_lcell_comb \Mux1~15 (
	.dataa(!\afi_wlat_r[0]~q ),
	.datab(!\doing_write_pipe[31]~q ),
	.datac(!\doing_write_pipe[30]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~15 .extended_lut = "off";
defparam \Mux1~15 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \Mux1~15 .shared_arith = "off";

arriaii_lcell_comb \Mux1~21 (
	.dataa(!\afi_wlat_r[0]~q ),
	.datab(!\doing_write_pipe[25]~q ),
	.datac(!\doing_write_pipe[26]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~21 .extended_lut = "off";
defparam \Mux1~21 .lut_mask = 64'h2727272727272727;
defparam \Mux1~21 .shared_arith = "off";

arriaii_lcell_comb \Mux1~25 (
	.dataa(!\afi_wlat_r[0]~q ),
	.datab(!\doing_write_pipe[29]~q ),
	.datac(!\doing_write_pipe[30]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~25 .extended_lut = "off";
defparam \Mux1~25 .lut_mask = 64'h2727272727272727;
defparam \Mux1~25 .shared_arith = "off";

arriaii_lcell_comb \Mux1~29 (
	.dataa(!\afi_wlat_r[0]~q ),
	.datab(!\doing_write_pipe[28]~q ),
	.datac(!\doing_write_pipe[27]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~29 .extended_lut = "off";
defparam \Mux1~29 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \Mux1~29 .shared_arith = "off";

arriaii_lcell_comb \Mux1~33 (
	.dataa(!\afi_wlat_r[0]~q ),
	.datab(!\doing_write_pipe[0]~q ),
	.datac(!\doing_write_pipe[31]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~33 .extended_lut = "off";
defparam \Mux1~33 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \Mux1~33 .shared_arith = "off";

arriaii_lcell_comb \afi_wlat_r[2]~0 (
	.dataa(!wd_lat_2),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\afi_wlat_r[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_wlat_r[2]~0 .extended_lut = "off";
defparam \afi_wlat_r[2]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \afi_wlat_r[2]~0 .shared_arith = "off";

dffeas ecc_wdata_fifo_read(
	.clk(ctl_clk),
	.d(\ecc_wdata_fifo_read~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ecc_wdata_fifo_read1),
	.prn(vcc));
defparam ecc_wdata_fifo_read.is_wysiwyg = "true";
defparam ecc_wdata_fifo_read.power_up = "low";

dffeas doing_read(
	.clk(ctl_clk),
	.d(\doing_read~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(doing_read1),
	.prn(vcc));
defparam doing_read.is_wysiwyg = "true";
defparam doing_read.power_up = "low";

arriaii_lcell_comb \afi_dm[4] (
	.dataa(!q_b_132),
	.datab(!\int_real_wdata_valid~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_dm_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_dm[4] .extended_lut = "off";
defparam \afi_dm[4] .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \afi_dm[4] .shared_arith = "off";

arriaii_lcell_comb \afi_dm[12] (
	.dataa(!\int_real_wdata_valid~q ),
	.datab(!q_b_140),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_dm_12),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_dm[12] .extended_lut = "off";
defparam \afi_dm[12] .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \afi_dm[12] .shared_arith = "off";

arriaii_lcell_comb \afi_dm[0] (
	.dataa(!\int_real_wdata_valid~q ),
	.datab(!q_b_128),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_dm_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_dm[0] .extended_lut = "off";
defparam \afi_dm[0] .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \afi_dm[0] .shared_arith = "off";

arriaii_lcell_comb \afi_dm[8] (
	.dataa(!\int_real_wdata_valid~q ),
	.datab(!q_b_136),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_dm_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_dm[8] .extended_lut = "off";
defparam \afi_dm[8] .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \afi_dm[8] .shared_arith = "off";

arriaii_lcell_comb \afi_dm[5] (
	.dataa(!\int_real_wdata_valid~q ),
	.datab(!q_b_133),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_dm_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_dm[5] .extended_lut = "off";
defparam \afi_dm[5] .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \afi_dm[5] .shared_arith = "off";

arriaii_lcell_comb \afi_dm[13] (
	.dataa(!\int_real_wdata_valid~q ),
	.datab(!q_b_141),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_dm_13),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_dm[13] .extended_lut = "off";
defparam \afi_dm[13] .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \afi_dm[13] .shared_arith = "off";

arriaii_lcell_comb \afi_dm[1] (
	.dataa(!\int_real_wdata_valid~q ),
	.datab(!q_b_129),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_dm_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_dm[1] .extended_lut = "off";
defparam \afi_dm[1] .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \afi_dm[1] .shared_arith = "off";

arriaii_lcell_comb \afi_dm[9] (
	.dataa(!\int_real_wdata_valid~q ),
	.datab(!q_b_137),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_dm_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_dm[9] .extended_lut = "off";
defparam \afi_dm[9] .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \afi_dm[9] .shared_arith = "off";

arriaii_lcell_comb \afi_dm[6] (
	.dataa(!\int_real_wdata_valid~q ),
	.datab(!q_b_134),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_dm_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_dm[6] .extended_lut = "off";
defparam \afi_dm[6] .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \afi_dm[6] .shared_arith = "off";

arriaii_lcell_comb \afi_dm[14] (
	.dataa(!\int_real_wdata_valid~q ),
	.datab(!q_b_142),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_dm_14),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_dm[14] .extended_lut = "off";
defparam \afi_dm[14] .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \afi_dm[14] .shared_arith = "off";

arriaii_lcell_comb \afi_dm[2] (
	.dataa(!\int_real_wdata_valid~q ),
	.datab(!q_b_130),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_dm_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_dm[2] .extended_lut = "off";
defparam \afi_dm[2] .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \afi_dm[2] .shared_arith = "off";

arriaii_lcell_comb \afi_dm[10] (
	.dataa(!\int_real_wdata_valid~q ),
	.datab(!q_b_138),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_dm_10),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_dm[10] .extended_lut = "off";
defparam \afi_dm[10] .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \afi_dm[10] .shared_arith = "off";

arriaii_lcell_comb \afi_dm[7] (
	.dataa(!\int_real_wdata_valid~q ),
	.datab(!q_b_135),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_dm_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_dm[7] .extended_lut = "off";
defparam \afi_dm[7] .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \afi_dm[7] .shared_arith = "off";

arriaii_lcell_comb \afi_dm[15] (
	.dataa(!\int_real_wdata_valid~q ),
	.datab(!q_b_143),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_dm_15),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_dm[15] .extended_lut = "off";
defparam \afi_dm[15] .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \afi_dm[15] .shared_arith = "off";

arriaii_lcell_comb \afi_dm[3] (
	.dataa(!\int_real_wdata_valid~q ),
	.datab(!q_b_131),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_dm_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_dm[3] .extended_lut = "off";
defparam \afi_dm[3] .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \afi_dm[3] .shared_arith = "off";

arriaii_lcell_comb \afi_dm[11] (
	.dataa(!\int_real_wdata_valid~q ),
	.datab(!q_b_139),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(afi_dm_11),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_dm[11] .extended_lut = "off";
defparam \afi_dm[11] .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \afi_dm[11] .shared_arith = "off";

dffeas int_wdata_valid(
	.clk(ctl_clk),
	.d(\int_wdata_valid~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(int_wdata_valid1),
	.prn(vcc));
defparam int_wdata_valid.is_wysiwyg = "true";
defparam int_wdata_valid.power_up = "low";

dffeas int_dqs_burst(
	.clk(ctl_clk),
	.d(\int_dqs_burst~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(int_dqs_burst1),
	.prn(vcc));
defparam int_dqs_burst.is_wysiwyg = "true";
defparam int_dqs_burst.power_up = "low";

dffeas int_dqs_burst_hr(
	.clk(ctl_clk),
	.d(\Mux3~4_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(int_dqs_burst_hr1),
	.prn(vcc));
defparam int_dqs_burst_hr.is_wysiwyg = "true";
defparam int_dqs_burst_hr.power_up = "low";

dffeas \rdwr_data_valid_pipe[0] (
	.clk(ctl_clk),
	.d(rdwr_data_valid),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_data_valid_pipe[0]~q ),
	.prn(vcc));
defparam \rdwr_data_valid_pipe[0] .is_wysiwyg = "true";
defparam \rdwr_data_valid_pipe[0] .power_up = "low";

dffeas \rdwr_data_valid_pipe[1] (
	.clk(ctl_clk),
	.d(\rdwr_data_valid_pipe[0]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_data_valid_pipe[1]~q ),
	.prn(vcc));
defparam \rdwr_data_valid_pipe[1] .is_wysiwyg = "true";
defparam \rdwr_data_valid_pipe[1] .power_up = "low";

dffeas \rdwr_data_valid_pipe[2] (
	.clk(ctl_clk),
	.d(\rdwr_data_valid_pipe[1]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_data_valid_pipe[2]~q ),
	.prn(vcc));
defparam \rdwr_data_valid_pipe[2] .is_wysiwyg = "true";
defparam \rdwr_data_valid_pipe[2] .power_up = "low";

dffeas \rdwr_data_valid_pipe[3] (
	.clk(ctl_clk),
	.d(\rdwr_data_valid_pipe[2]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_data_valid_pipe[3]~q ),
	.prn(vcc));
defparam \rdwr_data_valid_pipe[3] .is_wysiwyg = "true";
defparam \rdwr_data_valid_pipe[3] .power_up = "low";

dffeas \rdwr_data_valid_pipe[4] (
	.clk(ctl_clk),
	.d(\rdwr_data_valid_pipe[3]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_data_valid_pipe[4]~q ),
	.prn(vcc));
defparam \rdwr_data_valid_pipe[4] .is_wysiwyg = "true";
defparam \rdwr_data_valid_pipe[4] .power_up = "low";

dffeas \rdwr_data_valid_pipe[5] (
	.clk(ctl_clk),
	.d(\rdwr_data_valid_pipe[4]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_data_valid_pipe[5]~q ),
	.prn(vcc));
defparam \rdwr_data_valid_pipe[5] .is_wysiwyg = "true";
defparam \rdwr_data_valid_pipe[5] .power_up = "low";

dffeas \rdwr_data_valid_pipe[6] (
	.clk(ctl_clk),
	.d(\rdwr_data_valid_pipe[5]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_data_valid_pipe[6]~q ),
	.prn(vcc));
defparam \rdwr_data_valid_pipe[6] .is_wysiwyg = "true";
defparam \rdwr_data_valid_pipe[6] .power_up = "low";

dffeas \rdwr_data_valid_pipe[7] (
	.clk(ctl_clk),
	.d(\rdwr_data_valid_pipe[6]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_data_valid_pipe[7]~q ),
	.prn(vcc));
defparam \rdwr_data_valid_pipe[7] .is_wysiwyg = "true";
defparam \rdwr_data_valid_pipe[7] .power_up = "low";

dffeas \rdwr_data_valid_pipe[8] (
	.clk(ctl_clk),
	.d(\rdwr_data_valid_pipe[7]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_data_valid_pipe[8]~q ),
	.prn(vcc));
defparam \rdwr_data_valid_pipe[8] .is_wysiwyg = "true";
defparam \rdwr_data_valid_pipe[8] .power_up = "low";

dffeas \rdwr_data_valid_pipe[9] (
	.clk(ctl_clk),
	.d(\rdwr_data_valid_pipe[8]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_data_valid_pipe[9]~q ),
	.prn(vcc));
defparam \rdwr_data_valid_pipe[9] .is_wysiwyg = "true";
defparam \rdwr_data_valid_pipe[9] .power_up = "low";

dffeas \rdwr_data_valid_pipe[10] (
	.clk(ctl_clk),
	.d(\rdwr_data_valid_pipe[9]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_data_valid_pipe[10]~q ),
	.prn(vcc));
defparam \rdwr_data_valid_pipe[10] .is_wysiwyg = "true";
defparam \rdwr_data_valid_pipe[10] .power_up = "low";

dffeas \rdwr_data_valid_pipe[11] (
	.clk(ctl_clk),
	.d(\rdwr_data_valid_pipe[10]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_data_valid_pipe[11]~q ),
	.prn(vcc));
defparam \rdwr_data_valid_pipe[11] .is_wysiwyg = "true";
defparam \rdwr_data_valid_pipe[11] .power_up = "low";

dffeas \rdwr_data_valid_pipe[12] (
	.clk(ctl_clk),
	.d(\rdwr_data_valid_pipe[11]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_data_valid_pipe[12]~q ),
	.prn(vcc));
defparam \rdwr_data_valid_pipe[12] .is_wysiwyg = "true";
defparam \rdwr_data_valid_pipe[12] .power_up = "low";

dffeas \rdwr_data_valid_pipe[13] (
	.clk(ctl_clk),
	.d(\rdwr_data_valid_pipe[12]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_data_valid_pipe[13]~q ),
	.prn(vcc));
defparam \rdwr_data_valid_pipe[13] .is_wysiwyg = "true";
defparam \rdwr_data_valid_pipe[13] .power_up = "low";

dffeas \rdwr_data_valid_pipe[14] (
	.clk(ctl_clk),
	.d(\rdwr_data_valid_pipe[13]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_data_valid_pipe[14]~q ),
	.prn(vcc));
defparam \rdwr_data_valid_pipe[14] .is_wysiwyg = "true";
defparam \rdwr_data_valid_pipe[14] .power_up = "low";

dffeas \rdwr_data_valid_pipe[15] (
	.clk(ctl_clk),
	.d(\rdwr_data_valid_pipe[14]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_data_valid_pipe[15]~q ),
	.prn(vcc));
defparam \rdwr_data_valid_pipe[15] .is_wysiwyg = "true";
defparam \rdwr_data_valid_pipe[15] .power_up = "low";

dffeas \rdwr_data_valid_pipe[16] (
	.clk(ctl_clk),
	.d(\rdwr_data_valid_pipe[15]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_data_valid_pipe[16]~q ),
	.prn(vcc));
defparam \rdwr_data_valid_pipe[16] .is_wysiwyg = "true";
defparam \rdwr_data_valid_pipe[16] .power_up = "low";

dffeas \rdwr_data_valid_pipe[17] (
	.clk(ctl_clk),
	.d(\rdwr_data_valid_pipe[16]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_data_valid_pipe[17]~q ),
	.prn(vcc));
defparam \rdwr_data_valid_pipe[17] .is_wysiwyg = "true";
defparam \rdwr_data_valid_pipe[17] .power_up = "low";

dffeas \rdwr_data_valid_pipe[18] (
	.clk(ctl_clk),
	.d(\rdwr_data_valid_pipe[17]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_data_valid_pipe[18]~q ),
	.prn(vcc));
defparam \rdwr_data_valid_pipe[18] .is_wysiwyg = "true";
defparam \rdwr_data_valid_pipe[18] .power_up = "low";

dffeas \rdwr_data_valid_pipe[19] (
	.clk(ctl_clk),
	.d(\rdwr_data_valid_pipe[18]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_data_valid_pipe[19]~q ),
	.prn(vcc));
defparam \rdwr_data_valid_pipe[19] .is_wysiwyg = "true";
defparam \rdwr_data_valid_pipe[19] .power_up = "low";

dffeas \rdwr_data_valid_pipe[20] (
	.clk(ctl_clk),
	.d(\rdwr_data_valid_pipe[19]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_data_valid_pipe[20]~q ),
	.prn(vcc));
defparam \rdwr_data_valid_pipe[20] .is_wysiwyg = "true";
defparam \rdwr_data_valid_pipe[20] .power_up = "low";

dffeas \rdwr_data_valid_pipe[21] (
	.clk(ctl_clk),
	.d(\rdwr_data_valid_pipe[20]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_data_valid_pipe[21]~q ),
	.prn(vcc));
defparam \rdwr_data_valid_pipe[21] .is_wysiwyg = "true";
defparam \rdwr_data_valid_pipe[21] .power_up = "low";

dffeas \afi_wlat_r[1] (
	.clk(ctl_clk),
	.d(afi_wlat[1]),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\afi_wlat_r[1]~q ),
	.prn(vcc));
defparam \afi_wlat_r[1] .is_wysiwyg = "true";
defparam \afi_wlat_r[1] .power_up = "low";

arriaii_lcell_comb \Add0~0 (
	.dataa(!\afi_wlat_r[2]~q ),
	.datab(!\afi_wlat_r[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h9999999999999999;
defparam \Add0~0 .shared_arith = "off";

arriaii_lcell_comb \afi_wlat_r[0]~1 (
	.dataa(!wd_lat_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\afi_wlat_r[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \afi_wlat_r[0]~1 .extended_lut = "off";
defparam \afi_wlat_r[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \afi_wlat_r[0]~1 .shared_arith = "off";

dffeas \afi_wlat_r[0] (
	.clk(ctl_clk),
	.d(\afi_wlat_r[0]~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\afi_wlat_r[0]~q ),
	.prn(vcc));
defparam \afi_wlat_r[0] .is_wysiwyg = "true";
defparam \afi_wlat_r[0] .power_up = "low";

arriaii_lcell_comb \Mux0~8 (
	.dataa(!\rdwr_data_valid_pipe[19]~q ),
	.datab(!\rdwr_data_valid_pipe[17]~q ),
	.datac(!\rdwr_data_valid_pipe[16]~q ),
	.datad(!\afi_wlat_r[0]~q ),
	.datae(!\afi_wlat_r[1]~q ),
	.dataf(!\Add0~0_combout ),
	.datag(!\rdwr_data_valid_pipe[18]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~8 .extended_lut = "on";
defparam \Mux0~8 .lut_mask = 64'h0F550F3300FF00FF;
defparam \Mux0~8 .shared_arith = "off";

dffeas \rdwr_data_valid_pipe[22] (
	.clk(ctl_clk),
	.d(\rdwr_data_valid_pipe[21]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_data_valid_pipe[22]~q ),
	.prn(vcc));
defparam \rdwr_data_valid_pipe[22] .is_wysiwyg = "true";
defparam \rdwr_data_valid_pipe[22] .power_up = "low";

arriaii_lcell_comb \Mux0~12 (
	.dataa(!\rdwr_data_valid_pipe[23]~q ),
	.datab(!\rdwr_data_valid_pipe[21]~q ),
	.datac(!\rdwr_data_valid_pipe[20]~q ),
	.datad(!\Add0~0_combout ),
	.datae(!\afi_wlat_r[1]~q ),
	.dataf(!\Mux0~8_combout ),
	.datag(!\rdwr_data_valid_pipe[22]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~12 .extended_lut = "on";
defparam \Mux0~12 .lut_mask = 64'h000F000FFF55FF33;
defparam \Mux0~12 .shared_arith = "off";

arriaii_lcell_comb \Mux0~16 (
	.dataa(!\rdwr_data_valid_pipe[11]~q ),
	.datab(!\rdwr_data_valid_pipe[9]~q ),
	.datac(!\rdwr_data_valid_pipe[8]~q ),
	.datad(!\afi_wlat_r[0]~q ),
	.datae(!\afi_wlat_r[1]~q ),
	.dataf(!\Add0~0_combout ),
	.datag(!\rdwr_data_valid_pipe[10]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~16 .extended_lut = "on";
defparam \Mux0~16 .lut_mask = 64'h0F550F3300FF00FF;
defparam \Mux0~16 .shared_arith = "off";

arriaii_lcell_comb \Mux0~20 (
	.dataa(!\rdwr_data_valid_pipe[15]~q ),
	.datab(!\rdwr_data_valid_pipe[13]~q ),
	.datac(!\rdwr_data_valid_pipe[12]~q ),
	.datad(!\Add0~0_combout ),
	.datae(!\afi_wlat_r[1]~q ),
	.dataf(!\Mux0~16_combout ),
	.datag(!\rdwr_data_valid_pipe[14]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~20 .extended_lut = "on";
defparam \Mux0~20 .lut_mask = 64'h000F000FFF55FF33;
defparam \Mux0~20 .shared_arith = "off";

arriaii_lcell_comb \Mux0~24 (
	.dataa(!\rdwr_data_valid_pipe[3]~q ),
	.datab(!\rdwr_data_valid_pipe[1]~q ),
	.datac(!\rdwr_data_valid_pipe[0]~q ),
	.datad(!\afi_wlat_r[0]~q ),
	.datae(!\afi_wlat_r[1]~q ),
	.dataf(!\Add0~0_combout ),
	.datag(!\rdwr_data_valid_pipe[2]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~24 .extended_lut = "on";
defparam \Mux0~24 .lut_mask = 64'h0F550F3300FF00FF;
defparam \Mux0~24 .shared_arith = "off";

arriaii_lcell_comb \Mux0~28 (
	.dataa(!\rdwr_data_valid_pipe[7]~q ),
	.datab(!\rdwr_data_valid_pipe[5]~q ),
	.datac(!\rdwr_data_valid_pipe[4]~q ),
	.datad(!\Add0~0_combout ),
	.datae(!\afi_wlat_r[1]~q ),
	.dataf(!\Mux0~24_combout ),
	.datag(!\rdwr_data_valid_pipe[6]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~28 .extended_lut = "on";
defparam \Mux0~28 .lut_mask = 64'h000F000FFF55FF33;
defparam \Mux0~28 .shared_arith = "off";

dffeas \afi_wlat_r[3] (
	.clk(ctl_clk),
	.d(afi_wlat[3]),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\afi_wlat_r[3]~q ),
	.prn(vcc));
defparam \afi_wlat_r[3] .is_wysiwyg = "true";
defparam \afi_wlat_r[3] .power_up = "low";

arriaii_lcell_comb \Add0~1 (
	.dataa(!\afi_wlat_r[2]~q ),
	.datab(!\afi_wlat_r[1]~q ),
	.datac(!\afi_wlat_r[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h7878787878787878;
defparam \Add0~1 .shared_arith = "off";

dffeas \afi_wlat_r[4] (
	.clk(ctl_clk),
	.d(afi_wlat[4]),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\afi_wlat_r[4]~q ),
	.prn(vcc));
defparam \afi_wlat_r[4] .is_wysiwyg = "true";
defparam \afi_wlat_r[4] .power_up = "low";

arriaii_lcell_comb \Add0~2 (
	.dataa(!\afi_wlat_r[2]~q ),
	.datab(!\afi_wlat_r[1]~q ),
	.datac(!\afi_wlat_r[3]~q ),
	.datad(!\afi_wlat_r[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h7F807F807F807F80;
defparam \Add0~2 .shared_arith = "off";

arriaii_lcell_comb \Mux0~32 (
	.dataa(!\Mux0~4_combout ),
	.datab(!\Mux0~12_combout ),
	.datac(!\Mux0~20_combout ),
	.datad(!\Mux0~28_combout ),
	.datae(!\Add0~1_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~32 .extended_lut = "off";
defparam \Mux0~32 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux0~32 .shared_arith = "off";

arriaii_lcell_comb \doing_write~0 (
	.dataa(!do_write_r),
	.datab(!do_burst_chop_r),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_write~0 .extended_lut = "off";
defparam \doing_write~0 .lut_mask = 64'h4444444444444444;
defparam \doing_write~0 .shared_arith = "off";

dffeas doing_write(
	.clk(ctl_clk),
	.d(\doing_write~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write~q ),
	.prn(vcc));
defparam doing_write.is_wysiwyg = "true";
defparam doing_write.power_up = "low";

arriaii_lcell_comb \always8~0 (
	.dataa(!do_write_r),
	.datab(!\doing_write~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always8~0 .extended_lut = "off";
defparam \always8~0 .lut_mask = 64'h7777777777777777;
defparam \always8~0 .shared_arith = "off";

dffeas \doing_write_pipe[0] (
	.clk(ctl_clk),
	.d(\always8~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write_pipe[0]~q ),
	.prn(vcc));
defparam \doing_write_pipe[0] .is_wysiwyg = "true";
defparam \doing_write_pipe[0] .power_up = "low";

dffeas \doing_write_pipe[1] (
	.clk(ctl_clk),
	.d(\doing_write_pipe[0]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write_pipe[1]~q ),
	.prn(vcc));
defparam \doing_write_pipe[1] .is_wysiwyg = "true";
defparam \doing_write_pipe[1] .power_up = "low";

dffeas \doing_write_pipe[2] (
	.clk(ctl_clk),
	.d(\doing_write_pipe[1]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write_pipe[2]~q ),
	.prn(vcc));
defparam \doing_write_pipe[2] .is_wysiwyg = "true";
defparam \doing_write_pipe[2] .power_up = "low";

dffeas \doing_write_pipe[3] (
	.clk(ctl_clk),
	.d(\doing_write_pipe[2]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write_pipe[3]~q ),
	.prn(vcc));
defparam \doing_write_pipe[3] .is_wysiwyg = "true";
defparam \doing_write_pipe[3] .power_up = "low";

dffeas \doing_write_pipe[4] (
	.clk(ctl_clk),
	.d(\doing_write_pipe[3]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write_pipe[4]~q ),
	.prn(vcc));
defparam \doing_write_pipe[4] .is_wysiwyg = "true";
defparam \doing_write_pipe[4] .power_up = "low";

dffeas \doing_write_pipe[5] (
	.clk(ctl_clk),
	.d(\doing_write_pipe[4]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write_pipe[5]~q ),
	.prn(vcc));
defparam \doing_write_pipe[5] .is_wysiwyg = "true";
defparam \doing_write_pipe[5] .power_up = "low";

dffeas \doing_write_pipe[6] (
	.clk(ctl_clk),
	.d(\doing_write_pipe[5]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write_pipe[6]~q ),
	.prn(vcc));
defparam \doing_write_pipe[6] .is_wysiwyg = "true";
defparam \doing_write_pipe[6] .power_up = "low";

dffeas \doing_write_pipe[7] (
	.clk(ctl_clk),
	.d(\doing_write_pipe[6]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write_pipe[7]~q ),
	.prn(vcc));
defparam \doing_write_pipe[7] .is_wysiwyg = "true";
defparam \doing_write_pipe[7] .power_up = "low";

dffeas \doing_write_pipe[8] (
	.clk(ctl_clk),
	.d(\doing_write_pipe[7]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write_pipe[8]~q ),
	.prn(vcc));
defparam \doing_write_pipe[8] .is_wysiwyg = "true";
defparam \doing_write_pipe[8] .power_up = "low";

dffeas \doing_write_pipe[9] (
	.clk(ctl_clk),
	.d(\doing_write_pipe[8]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write_pipe[9]~q ),
	.prn(vcc));
defparam \doing_write_pipe[9] .is_wysiwyg = "true";
defparam \doing_write_pipe[9] .power_up = "low";

dffeas \doing_write_pipe[10] (
	.clk(ctl_clk),
	.d(\doing_write_pipe[9]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write_pipe[10]~q ),
	.prn(vcc));
defparam \doing_write_pipe[10] .is_wysiwyg = "true";
defparam \doing_write_pipe[10] .power_up = "low";

dffeas \doing_write_pipe[11] (
	.clk(ctl_clk),
	.d(\doing_write_pipe[10]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write_pipe[11]~q ),
	.prn(vcc));
defparam \doing_write_pipe[11] .is_wysiwyg = "true";
defparam \doing_write_pipe[11] .power_up = "low";

dffeas \doing_write_pipe[12] (
	.clk(ctl_clk),
	.d(\doing_write_pipe[11]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write_pipe[12]~q ),
	.prn(vcc));
defparam \doing_write_pipe[12] .is_wysiwyg = "true";
defparam \doing_write_pipe[12] .power_up = "low";

dffeas \doing_write_pipe[13] (
	.clk(ctl_clk),
	.d(\doing_write_pipe[12]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write_pipe[13]~q ),
	.prn(vcc));
defparam \doing_write_pipe[13] .is_wysiwyg = "true";
defparam \doing_write_pipe[13] .power_up = "low";

dffeas \doing_write_pipe[14] (
	.clk(ctl_clk),
	.d(\doing_write_pipe[13]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write_pipe[14]~q ),
	.prn(vcc));
defparam \doing_write_pipe[14] .is_wysiwyg = "true";
defparam \doing_write_pipe[14] .power_up = "low";

dffeas \doing_write_pipe[15] (
	.clk(ctl_clk),
	.d(\doing_write_pipe[14]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write_pipe[15]~q ),
	.prn(vcc));
defparam \doing_write_pipe[15] .is_wysiwyg = "true";
defparam \doing_write_pipe[15] .power_up = "low";

dffeas \doing_write_pipe[16] (
	.clk(ctl_clk),
	.d(\doing_write_pipe[15]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write_pipe[16]~q ),
	.prn(vcc));
defparam \doing_write_pipe[16] .is_wysiwyg = "true";
defparam \doing_write_pipe[16] .power_up = "low";

dffeas \doing_write_pipe[17] (
	.clk(ctl_clk),
	.d(\doing_write_pipe[16]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write_pipe[17]~q ),
	.prn(vcc));
defparam \doing_write_pipe[17] .is_wysiwyg = "true";
defparam \doing_write_pipe[17] .power_up = "low";

arriaii_lcell_comb \Mux1~1 (
	.dataa(!\afi_wlat_r[0]~q ),
	.datab(!\doing_write_pipe[17]~q ),
	.datac(!\doing_write_pipe[16]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~1 .extended_lut = "off";
defparam \Mux1~1 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \Mux1~1 .shared_arith = "off";

arriaii_lcell_comb \Mux1~2 (
	.dataa(!\afi_wlat_r[0]~q ),
	.datab(!\doing_write_pipe[9]~q ),
	.datac(!\doing_write_pipe[8]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~2 .extended_lut = "off";
defparam \Mux1~2 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \Mux1~2 .shared_arith = "off";

arriaii_lcell_comb \Mux1~3 (
	.dataa(!\afi_wlat_r[0]~q ),
	.datab(!\doing_write_pipe[1]~q ),
	.datac(!\doing_write_pipe[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~3 .extended_lut = "off";
defparam \Mux1~3 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \Mux1~3 .shared_arith = "off";

arriaii_lcell_comb \Mux1~4 (
	.dataa(!\Mux1~0_combout ),
	.datab(!\Mux1~1_combout ),
	.datac(!\Mux1~2_combout ),
	.datad(!\Mux1~3_combout ),
	.datae(!\Add0~1_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~4 .extended_lut = "off";
defparam \Mux1~4 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux1~4 .shared_arith = "off";

dffeas \doing_write_pipe[18] (
	.clk(ctl_clk),
	.d(\doing_write_pipe[17]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write_pipe[18]~q ),
	.prn(vcc));
defparam \doing_write_pipe[18] .is_wysiwyg = "true";
defparam \doing_write_pipe[18] .power_up = "low";

dffeas \doing_write_pipe[19] (
	.clk(ctl_clk),
	.d(\doing_write_pipe[18]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write_pipe[19]~q ),
	.prn(vcc));
defparam \doing_write_pipe[19] .is_wysiwyg = "true";
defparam \doing_write_pipe[19] .power_up = "low";

dffeas \doing_write_pipe[20] (
	.clk(ctl_clk),
	.d(\doing_write_pipe[19]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write_pipe[20]~q ),
	.prn(vcc));
defparam \doing_write_pipe[20] .is_wysiwyg = "true";
defparam \doing_write_pipe[20] .power_up = "low";

dffeas \doing_write_pipe[21] (
	.clk(ctl_clk),
	.d(\doing_write_pipe[20]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write_pipe[21]~q ),
	.prn(vcc));
defparam \doing_write_pipe[21] .is_wysiwyg = "true";
defparam \doing_write_pipe[21] .power_up = "low";

arriaii_lcell_comb \Mux1~6 (
	.dataa(!\afi_wlat_r[0]~q ),
	.datab(!\doing_write_pipe[21]~q ),
	.datac(!\doing_write_pipe[20]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~6 .extended_lut = "off";
defparam \Mux1~6 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \Mux1~6 .shared_arith = "off";

arriaii_lcell_comb \Mux1~7 (
	.dataa(!\afi_wlat_r[0]~q ),
	.datab(!\doing_write_pipe[13]~q ),
	.datac(!\doing_write_pipe[12]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~7 .extended_lut = "off";
defparam \Mux1~7 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \Mux1~7 .shared_arith = "off";

arriaii_lcell_comb \Mux1~8 (
	.dataa(!\afi_wlat_r[0]~q ),
	.datab(!\doing_write_pipe[5]~q ),
	.datac(!\doing_write_pipe[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~8 .extended_lut = "off";
defparam \Mux1~8 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \Mux1~8 .shared_arith = "off";

arriaii_lcell_comb \Mux1~9 (
	.dataa(!\Mux1~5_combout ),
	.datab(!\Mux1~6_combout ),
	.datac(!\Mux1~7_combout ),
	.datad(!\Mux1~8_combout ),
	.datae(!\Add0~1_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~9 .extended_lut = "off";
defparam \Mux1~9 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux1~9 .shared_arith = "off";

arriaii_lcell_comb \Mux1~11 (
	.dataa(!\afi_wlat_r[0]~q ),
	.datab(!\doing_write_pipe[19]~q ),
	.datac(!\doing_write_pipe[18]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~11 .extended_lut = "off";
defparam \Mux1~11 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \Mux1~11 .shared_arith = "off";

arriaii_lcell_comb \Mux1~12 (
	.dataa(!\afi_wlat_r[0]~q ),
	.datab(!\doing_write_pipe[11]~q ),
	.datac(!\doing_write_pipe[10]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~12 .extended_lut = "off";
defparam \Mux1~12 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \Mux1~12 .shared_arith = "off";

arriaii_lcell_comb \Mux1~13 (
	.dataa(!\afi_wlat_r[0]~q ),
	.datab(!\doing_write_pipe[3]~q ),
	.datac(!\doing_write_pipe[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~13 .extended_lut = "off";
defparam \Mux1~13 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \Mux1~13 .shared_arith = "off";

arriaii_lcell_comb \Mux1~14 (
	.dataa(!\Mux1~10_combout ),
	.datab(!\Mux1~11_combout ),
	.datac(!\Mux1~12_combout ),
	.datad(!\Mux1~13_combout ),
	.datae(!\Add0~1_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~14 .extended_lut = "off";
defparam \Mux1~14 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux1~14 .shared_arith = "off";

dffeas \doing_write_pipe[22] (
	.clk(ctl_clk),
	.d(\doing_write_pipe[21]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write_pipe[22]~q ),
	.prn(vcc));
defparam \doing_write_pipe[22] .is_wysiwyg = "true";
defparam \doing_write_pipe[22] .power_up = "low";

dffeas \doing_write_pipe[23] (
	.clk(ctl_clk),
	.d(\doing_write_pipe[22]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write_pipe[23]~q ),
	.prn(vcc));
defparam \doing_write_pipe[23] .is_wysiwyg = "true";
defparam \doing_write_pipe[23] .power_up = "low";

arriaii_lcell_comb \Mux1~16 (
	.dataa(!\afi_wlat_r[0]~q ),
	.datab(!\doing_write_pipe[23]~q ),
	.datac(!\doing_write_pipe[22]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~16 .extended_lut = "off";
defparam \Mux1~16 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \Mux1~16 .shared_arith = "off";

arriaii_lcell_comb \Mux1~17 (
	.dataa(!\afi_wlat_r[0]~q ),
	.datab(!\doing_write_pipe[15]~q ),
	.datac(!\doing_write_pipe[14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~17 .extended_lut = "off";
defparam \Mux1~17 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \Mux1~17 .shared_arith = "off";

arriaii_lcell_comb \Mux1~18 (
	.dataa(!\afi_wlat_r[0]~q ),
	.datab(!\doing_write_pipe[7]~q ),
	.datac(!\doing_write_pipe[6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~18 .extended_lut = "off";
defparam \Mux1~18 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \Mux1~18 .shared_arith = "off";

arriaii_lcell_comb \Mux1~19 (
	.dataa(!\Mux1~15_combout ),
	.datab(!\Mux1~16_combout ),
	.datac(!\Mux1~17_combout ),
	.datad(!\Mux1~18_combout ),
	.datae(!\Add0~1_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~19 .extended_lut = "off";
defparam \Mux1~19 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux1~19 .shared_arith = "off";

arriaii_lcell_comb \Mux1~20 (
	.dataa(!\afi_wlat_r[2]~q ),
	.datab(!\afi_wlat_r[1]~q ),
	.datac(!\Mux1~4_combout ),
	.datad(!\Mux1~9_combout ),
	.datae(!\Mux1~14_combout ),
	.dataf(!\Mux1~19_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~20 .extended_lut = "off";
defparam \Mux1~20 .lut_mask = 64'h021346578A9BCEDF;
defparam \Mux1~20 .shared_arith = "off";

arriaii_lcell_comb \Equal0~0 (
	.dataa(!\afi_wlat_r[2]~q ),
	.datab(!\afi_wlat_r[1]~q ),
	.datac(!\afi_wlat_r[3]~q ),
	.datad(!\afi_wlat_r[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h8000800080008000;
defparam \Equal0~0 .shared_arith = "off";

arriaii_lcell_comb \ecc_wdata_fifo_read~0 (
	.dataa(!\Mux0~32_combout ),
	.datab(!\Mux1~20_combout ),
	.datac(!\Equal0~0_combout ),
	.datad(!rdwr_data_valid),
	.datae(!\always8~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ecc_wdata_fifo_read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ecc_wdata_fifo_read~0 .extended_lut = "off";
defparam \ecc_wdata_fifo_read~0 .lut_mask = 64'h1010101F1010101F;
defparam \ecc_wdata_fifo_read~0 .shared_arith = "off";

arriaii_lcell_comb \doing_read~0 (
	.dataa(!do_read_r),
	.datab(!do_burst_chop_r),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_read~0 .extended_lut = "off";
defparam \doing_read~0 .lut_mask = 64'h4444444444444444;
defparam \doing_read~0 .shared_arith = "off";

dffeas int_real_wdata_valid(
	.clk(ctl_clk),
	.d(ecc_wdata_fifo_read1),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\int_real_wdata_valid~q ),
	.prn(vcc));
defparam int_real_wdata_valid.is_wysiwyg = "true";
defparam int_real_wdata_valid.power_up = "low";

arriaii_lcell_comb \Mux1~22 (
	.dataa(!\afi_wlat_r[0]~q ),
	.datab(!\doing_write_pipe[17]~q ),
	.datac(!\doing_write_pipe[18]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~22 .extended_lut = "off";
defparam \Mux1~22 .lut_mask = 64'h2727272727272727;
defparam \Mux1~22 .shared_arith = "off";

arriaii_lcell_comb \Mux1~23 (
	.dataa(!\afi_wlat_r[0]~q ),
	.datab(!\doing_write_pipe[9]~q ),
	.datac(!\doing_write_pipe[10]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~23 .extended_lut = "off";
defparam \Mux1~23 .lut_mask = 64'h2727272727272727;
defparam \Mux1~23 .shared_arith = "off";

arriaii_lcell_comb \Mux1~24 (
	.dataa(!\afi_wlat_r[0]~q ),
	.datab(!\doing_write_pipe[1]~q ),
	.datac(!\doing_write_pipe[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~24 .extended_lut = "off";
defparam \Mux1~24 .lut_mask = 64'h2727272727272727;
defparam \Mux1~24 .shared_arith = "off";

arriaii_lcell_comb \Mux3~0 (
	.dataa(!\Mux1~21_combout ),
	.datab(!\Mux1~22_combout ),
	.datac(!\Mux1~23_combout ),
	.datad(!\Mux1~24_combout ),
	.datae(!\Add0~1_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux3~0 .extended_lut = "off";
defparam \Mux3~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux3~0 .shared_arith = "off";

arriaii_lcell_comb \Mux1~26 (
	.dataa(!\afi_wlat_r[0]~q ),
	.datab(!\doing_write_pipe[21]~q ),
	.datac(!\doing_write_pipe[22]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~26 .extended_lut = "off";
defparam \Mux1~26 .lut_mask = 64'h2727272727272727;
defparam \Mux1~26 .shared_arith = "off";

arriaii_lcell_comb \Mux1~27 (
	.dataa(!\afi_wlat_r[0]~q ),
	.datab(!\doing_write_pipe[13]~q ),
	.datac(!\doing_write_pipe[14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~27 .extended_lut = "off";
defparam \Mux1~27 .lut_mask = 64'h2727272727272727;
defparam \Mux1~27 .shared_arith = "off";

arriaii_lcell_comb \Mux1~28 (
	.dataa(!\afi_wlat_r[0]~q ),
	.datab(!\doing_write_pipe[5]~q ),
	.datac(!\doing_write_pipe[6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~28 .extended_lut = "off";
defparam \Mux1~28 .lut_mask = 64'h2727272727272727;
defparam \Mux1~28 .shared_arith = "off";

arriaii_lcell_comb \Mux3~1 (
	.dataa(!\Mux1~25_combout ),
	.datab(!\Mux1~26_combout ),
	.datac(!\Mux1~27_combout ),
	.datad(!\Mux1~28_combout ),
	.datae(!\Add0~1_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux3~1 .extended_lut = "off";
defparam \Mux3~1 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux3~1 .shared_arith = "off";

arriaii_lcell_comb \Mux1~30 (
	.dataa(!\afi_wlat_r[0]~q ),
	.datab(!\doing_write_pipe[20]~q ),
	.datac(!\doing_write_pipe[19]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~30 .extended_lut = "off";
defparam \Mux1~30 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \Mux1~30 .shared_arith = "off";

arriaii_lcell_comb \Mux1~31 (
	.dataa(!\afi_wlat_r[0]~q ),
	.datab(!\doing_write_pipe[12]~q ),
	.datac(!\doing_write_pipe[11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~31 .extended_lut = "off";
defparam \Mux1~31 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \Mux1~31 .shared_arith = "off";

arriaii_lcell_comb \Mux1~32 (
	.dataa(!\afi_wlat_r[0]~q ),
	.datab(!\doing_write_pipe[4]~q ),
	.datac(!\doing_write_pipe[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~32 .extended_lut = "off";
defparam \Mux1~32 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \Mux1~32 .shared_arith = "off";

arriaii_lcell_comb \Mux3~2 (
	.dataa(!\Mux1~29_combout ),
	.datab(!\Mux1~30_combout ),
	.datac(!\Mux1~31_combout ),
	.datad(!\Mux1~32_combout ),
	.datae(!\Add0~1_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux3~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux3~2 .extended_lut = "off";
defparam \Mux3~2 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux3~2 .shared_arith = "off";

dffeas \doing_write_pipe[24] (
	.clk(ctl_clk),
	.d(\doing_write_pipe[23]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_write_pipe[24]~q ),
	.prn(vcc));
defparam \doing_write_pipe[24] .is_wysiwyg = "true";
defparam \doing_write_pipe[24] .power_up = "low";

arriaii_lcell_comb \Mux1~34 (
	.dataa(!\afi_wlat_r[0]~q ),
	.datab(!\doing_write_pipe[24]~q ),
	.datac(!\doing_write_pipe[23]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~34 .extended_lut = "off";
defparam \Mux1~34 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \Mux1~34 .shared_arith = "off";

arriaii_lcell_comb \Mux1~35 (
	.dataa(!\afi_wlat_r[0]~q ),
	.datab(!\doing_write_pipe[16]~q ),
	.datac(!\doing_write_pipe[15]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~35 .extended_lut = "off";
defparam \Mux1~35 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \Mux1~35 .shared_arith = "off";

arriaii_lcell_comb \Mux1~36 (
	.dataa(!\afi_wlat_r[0]~q ),
	.datab(!\doing_write_pipe[8]~q ),
	.datac(!\doing_write_pipe[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~36 .extended_lut = "off";
defparam \Mux1~36 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \Mux1~36 .shared_arith = "off";

arriaii_lcell_comb \Mux3~3 (
	.dataa(!\Mux1~33_combout ),
	.datab(!\Mux1~34_combout ),
	.datac(!\Mux1~35_combout ),
	.datad(!\Mux1~36_combout ),
	.datae(!\Add0~1_combout ),
	.dataf(!\Add0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux3~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux3~3 .extended_lut = "off";
defparam \Mux3~3 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux3~3 .shared_arith = "off";

arriaii_lcell_comb \Mux3~4 (
	.dataa(!\afi_wlat_r[2]~q ),
	.datab(!\afi_wlat_r[1]~q ),
	.datac(!\Mux3~0_combout ),
	.datad(!\Mux3~1_combout ),
	.datae(!\Mux3~2_combout ),
	.dataf(!\Mux3~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux3~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux3~4 .extended_lut = "off";
defparam \Mux3~4 .lut_mask = 64'h021346578A9BCEDF;
defparam \Mux3~4 .shared_arith = "off";

arriaii_lcell_comb \int_wdata_valid~0 (
	.dataa(!do_write_r),
	.datab(!\afi_wlat_r[0]~q ),
	.datac(!\Mux1~3_combout ),
	.datad(!\Equal0~0_combout ),
	.datae(!\Mux3~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_wdata_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_wdata_valid~0 .extended_lut = "off";
defparam \int_wdata_valid~0 .lut_mask = 64'h004CFF7F004CFF7F;
defparam \int_wdata_valid~0 .shared_arith = "off";

arriaii_lcell_comb \int_dqs_burst~0 (
	.dataa(!do_write_r),
	.datab(!\doing_write_pipe[0]~q ),
	.datac(!\Mux1~20_combout ),
	.datad(!\Equal0~0_combout ),
	.datae(!\Mux3~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_dqs_burst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_dqs_burst~0 .extended_lut = "off";
defparam \int_dqs_burst~0 .lut_mask = 64'h0F77FF770F77FF77;
defparam \int_dqs_burst~0 .shared_arith = "off";

endmodule

module ddr3_int_alt_ddrx_bank_timer_wrapper (
	clk_0,
	auto_refresh_logic_per_chip0int_refresh_req,
	out_cmd_info_valid_0,
	do_read_r,
	do_auto_precharge_r,
	do_write_r,
	out_cmd_info_valid_2,
	out_cmd_info_valid_3,
	out_cmd_info_valid_4,
	out_cmd_info_valid_1,
	pipe_10_0,
	pipe_12_0,
	pipe_11_0,
	pipe_12_2,
	pipe_12_3,
	pipe_12_1,
	pipe_10_2,
	pipe_10_3,
	pipe_10_1,
	pipe_11_2,
	pipe_11_3,
	pipe_11_1,
	do_burst_chop_r,
	pipe_12_4,
	pipe_11_4,
	pipe_10_4,
	fetch,
	do_precharge_all_r,
	out_cs_can_refresh_0,
	pipefull_0,
	do_refresh_r,
	add_lat_on,
	out_cmd_can_activate_0,
	out_cmd_bank_is_open_0,
	can_al_activate_write,
	to_chip_r_0,
	always38,
	to_bank_addr_r_2,
	current_bank_2,
	to_bank_addr_r_0,
	current_bank_0,
	to_bank_addr_r_1,
	current_bank_1,
	always381,
	out_cmd_can_write_0,
	can_al_activate_read,
	out_cmd_can_read_0,
	out_cs_all_banks_closed_0,
	out_cs_can_precharge_all_0,
	do_activate_r,
	reset_reg_11,
	pipefull_1,
	reset_reg_9,
	reset_reg_12,
	out_cmd_can_activate_2,
	out_cmd_bank_is_open_2,
	out_cmd_can_activate_3,
	out_cmd_bank_is_open_3,
	out_cmd_can_activate_4,
	out_cmd_bank_is_open_4,
	out_cmd_can_activate_1,
	out_cmd_bank_is_open_1,
	reset_reg_8,
	pipefull_4,
	pipefull_2,
	reset_reg_10,
	pipefull_3,
	always1,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	clk_0;
output 	auto_refresh_logic_per_chip0int_refresh_req;
output 	out_cmd_info_valid_0;
input 	do_read_r;
input 	do_auto_precharge_r;
input 	do_write_r;
output 	out_cmd_info_valid_2;
output 	out_cmd_info_valid_3;
output 	out_cmd_info_valid_4;
output 	out_cmd_info_valid_1;
input 	pipe_10_0;
input 	pipe_12_0;
input 	pipe_11_0;
input 	pipe_12_2;
input 	pipe_12_3;
input 	pipe_12_1;
input 	pipe_10_2;
input 	pipe_10_3;
input 	pipe_10_1;
input 	pipe_11_2;
input 	pipe_11_3;
input 	pipe_11_1;
input 	do_burst_chop_r;
input 	pipe_12_4;
input 	pipe_11_4;
input 	pipe_10_4;
input 	fetch;
input 	do_precharge_all_r;
output 	out_cs_can_refresh_0;
input 	pipefull_0;
input 	do_refresh_r;
output 	add_lat_on;
output 	out_cmd_can_activate_0;
output 	out_cmd_bank_is_open_0;
output 	can_al_activate_write;
input 	to_chip_r_0;
input 	always38;
input 	to_bank_addr_r_2;
input 	current_bank_2;
input 	to_bank_addr_r_0;
input 	current_bank_0;
input 	to_bank_addr_r_1;
input 	current_bank_1;
input 	always381;
output 	out_cmd_can_write_0;
output 	can_al_activate_read;
output 	out_cmd_can_read_0;
output 	out_cs_all_banks_closed_0;
output 	out_cs_can_precharge_all_0;
input 	do_activate_r;
input 	reset_reg_11;
input 	pipefull_1;
input 	reset_reg_9;
input 	reset_reg_12;
output 	out_cmd_can_activate_2;
output 	out_cmd_bank_is_open_2;
output 	out_cmd_can_activate_3;
output 	out_cmd_bank_is_open_3;
output 	out_cmd_can_activate_4;
output 	out_cmd_bank_is_open_4;
output 	out_cmd_can_activate_1;
output 	out_cmd_bank_is_open_1;
input 	reset_reg_8;
input 	pipefull_4;
input 	pipefull_2;
input 	reset_reg_10;
input 	pipefull_3;
output 	always1;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \rank_monitor_inst|act_cmd_monitor_per_chip[0].act_cmd_cnt[0]~q ;
wire \rank_monitor_inst|act_trrd_ready[0]~q ;
wire \bank_timer_inst|Mux0~4_combout ;
wire \rank_monitor_inst|write_dqs_ready~q ;
wire \rank_monitor_inst|read_dqs_ready~q ;
wire \bank_timer_inst|Mux25~4_combout ;
wire \bank_timer_inst|Mux5~4_combout ;
wire \bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[7].bank_timer_info_inst|act_ready~combout ;
wire \bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[5].bank_timer_info_inst|act_ready~combout ;
wire \bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[6].bank_timer_info_inst|act_ready~combout ;
wire \bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[1].bank_timer_info_inst|act_ready~combout ;
wire \bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[0].bank_timer_info_inst|act_ready~combout ;
wire \rank_monitor_inst|power_saving_logic_per_chip[0].int_enter_power_saving_ready~q ;
wire \bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[4].bank_timer_info_inst|act_ready~combout ;
wire \bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[2].bank_timer_info_inst|act_ready~combout ;
wire \bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[3].bank_timer_info_inst|act_ready~combout ;
wire \rank_monitor_inst|Selector20~0_combout ;
wire \timing_param_inst|act_to_rdwr[1]~q ;
wire \cache_inst|int_cmd_info_valid~0_combout ;
wire \bank_timer_inst|Mux10~2_combout ;
wire \bank_timer_inst|Mux13~2_combout ;
wire \bank_timer_inst|always106~0_combout ;
wire \bypass_inst|always145~0_combout ;
wire \rank_monitor_inst|act_cmd_monitor_per_chip[0].act_cmd_cnt[1]~q ;
wire \rank_monitor_inst|act_cmd_monitor_per_chip[0].act_cmd_cnt[2]~q ;
wire \bank_timer_inst|Mux1~2_combout ;
wire \timing_param_inst|more_than_3_wr_to_pch~q ;
wire \bank_timer_inst|can_al_activate_write~0_combout ;
wire \bank_timer_inst|Mux12~0_combout ;
wire \bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[0].bank_timer_info_inst|rdwr_ready~q ;
wire \bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[4].bank_timer_info_inst|rdwr_ready~q ;
wire \bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[2].bank_timer_info_inst|rdwr_ready~q ;
wire \bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[6].bank_timer_info_inst|rdwr_ready~q ;
wire \bank_timer_inst|Mux9~0_combout ;
wire \rank_monitor_inst|write_to_read_finish_twtr[0]~q ;
wire \bank_timer_inst|can_al_activate_read~0_combout ;
wire \bank_timer_inst|cs_all_banks_closed[0]~q ;
wire \bypass_inst|always140~0_combout ;
wire \bank_timer_inst|Mux16~2_combout ;
wire \bank_timer_inst|Mux19~2_combout ;
wire \bank_timer_inst|Mux3~2_combout ;
wire \bank_timer_inst|Mux2~2_combout ;
wire \bank_timer_inst|Mux22~2_combout ;
wire \bank_timer_inst|Mux4~2_combout ;
wire \bypass_inst|always71~0_combout ;


ddr3_int_alt_ddrx_rank_monitor rank_monitor_inst(
	.ctl_clk(clk_0),
	.auto_refresh_logic_per_chip0int_refresh_req(auto_refresh_logic_per_chip0int_refresh_req),
	.do_read_r(do_read_r),
	.do_write_r(do_write_r),
	.act_cmd_monitor_per_chip0act_cmd_cnt0(\rank_monitor_inst|act_cmd_monitor_per_chip[0].act_cmd_cnt[0]~q ),
	.act_trrd_ready_0(\rank_monitor_inst|act_trrd_ready[0]~q ),
	.write_dqs_ready1(\rank_monitor_inst|write_dqs_ready~q ),
	.read_dqs_ready1(\rank_monitor_inst|read_dqs_ready~q ),
	.do_burst_chop_r(do_burst_chop_r),
	.do_precharge_all_r(do_precharge_all_r),
	.do_refresh_r(do_refresh_r),
	.add_lat_on(add_lat_on),
	.to_chip_r_0(to_chip_r_0),
	.power_saving_logic_per_chip0int_enter_power_saving_ready(\rank_monitor_inst|power_saving_logic_per_chip[0].int_enter_power_saving_ready~q ),
	.Selector20(\rank_monitor_inst|Selector20~0_combout ),
	.act_to_rdwr_1(\timing_param_inst|act_to_rdwr[1]~q ),
	.ctl_reset_n(reset_reg_9),
	.always145(\bypass_inst|always145~0_combout ),
	.act_cmd_monitor_per_chip0act_cmd_cnt1(\rank_monitor_inst|act_cmd_monitor_per_chip[0].act_cmd_cnt[1]~q ),
	.act_cmd_monitor_per_chip0act_cmd_cnt2(\rank_monitor_inst|act_cmd_monitor_per_chip[0].act_cmd_cnt[2]~q ),
	.write_to_read_finish_twtr_0(\rank_monitor_inst|write_to_read_finish_twtr[0]~q ),
	.always1(always1),
	.always71(\bypass_inst|always71~0_combout ),
	.GND_port(GND_port));

ddr3_int_alt_ddrx_cache cache_inst(
	.ctl_clk(clk_0),
	.fetch(fetch),
	.int_cmd_info_valid(\cache_inst|int_cmd_info_valid~0_combout ),
	.ctl_reset_n(reset_reg_10));

ddr3_int_alt_ddrx_bypass bypass_inst(
	.ctl_clk(clk_0),
	.out_cmd_info_valid_0(out_cmd_info_valid_0),
	.do_read(do_read_r),
	.do_auto_precharge(do_auto_precharge_r),
	.do_write(do_write_r),
	.out_cmd_info_valid_2(out_cmd_info_valid_2),
	.out_cmd_info_valid_3(out_cmd_info_valid_3),
	.out_cmd_info_valid_4(out_cmd_info_valid_4),
	.out_cmd_info_valid_1(out_cmd_info_valid_1),
	.pipe_10_0(pipe_10_0),
	.pipe_12_0(pipe_12_0),
	.pipe_11_0(pipe_11_0),
	.act_cmd_monitor_per_chip0act_cmd_cnt0(\rank_monitor_inst|act_cmd_monitor_per_chip[0].act_cmd_cnt[0]~q ),
	.act_trrd_ready_0(\rank_monitor_inst|act_trrd_ready[0]~q ),
	.Mux0(\bank_timer_inst|Mux0~4_combout ),
	.pipe_12_2(pipe_12_2),
	.pipe_12_3(pipe_12_3),
	.pipe_12_1(pipe_12_1),
	.pipe_10_2(pipe_10_2),
	.pipe_10_3(pipe_10_3),
	.pipe_10_1(pipe_10_1),
	.pipe_11_2(pipe_11_2),
	.pipe_11_3(pipe_11_3),
	.pipe_11_1(pipe_11_1),
	.pipe_12_4(pipe_12_4),
	.pipe_11_4(pipe_11_4),
	.pipe_10_4(pipe_10_4),
	.Mux25(\bank_timer_inst|Mux25~4_combout ),
	.Mux5(\bank_timer_inst|Mux5~4_combout ),
	.fetch(fetch),
	.do_precharge_all(do_precharge_all_r),
	.out_cs_can_refresh_0(out_cs_can_refresh_0),
	.pipefull_0(pipefull_0),
	.out_cmd_can_activate_0(out_cmd_can_activate_0),
	.out_cmd_bank_is_open_0(out_cmd_bank_is_open_0),
	.to_chip({to_chip_r_0}),
	.always38(always38),
	.to_bank_addr_r_2(to_bank_addr_r_2),
	.current_bank_2(current_bank_2),
	.to_bank_addr_r_0(to_bank_addr_r_0),
	.current_bank_0(current_bank_0),
	.to_bank_addr_r_1(to_bank_addr_r_1),
	.current_bank_1(current_bank_1),
	.always381(always381),
	.out_cmd_can_write_0(out_cmd_can_write_0),
	.out_cmd_can_read_0(out_cmd_can_read_0),
	.out_cs_all_banks_closed_0(out_cs_all_banks_closed_0),
	.out_cs_can_precharge_all_0(out_cs_can_precharge_all_0),
	.do_activate(do_activate_r),
	.act_ready(\bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[7].bank_timer_info_inst|act_ready~combout ),
	.act_ready1(\bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[5].bank_timer_info_inst|act_ready~combout ),
	.act_ready2(\bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[6].bank_timer_info_inst|act_ready~combout ),
	.act_ready3(\bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[1].bank_timer_info_inst|act_ready~combout ),
	.act_ready4(\bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[0].bank_timer_info_inst|act_ready~combout ),
	.power_saving_logic_per_chip0int_enter_power_saving_ready(\rank_monitor_inst|power_saving_logic_per_chip[0].int_enter_power_saving_ready~q ),
	.act_ready5(\bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[4].bank_timer_info_inst|act_ready~combout ),
	.act_ready6(\bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[2].bank_timer_info_inst|act_ready~combout ),
	.act_ready7(\bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[3].bank_timer_info_inst|act_ready~combout ),
	.Selector20(\rank_monitor_inst|Selector20~0_combout ),
	.ctl_reset_n(reset_reg_11),
	.pipefull_1(pipefull_1),
	.act_to_rdwr_1(\timing_param_inst|act_to_rdwr[1]~q ),
	.int_cmd_info_valid(\cache_inst|int_cmd_info_valid~0_combout ),
	.out_cmd_can_activate_2(out_cmd_can_activate_2),
	.out_cmd_bank_is_open_2(out_cmd_bank_is_open_2),
	.out_cmd_can_activate_3(out_cmd_can_activate_3),
	.out_cmd_bank_is_open_3(out_cmd_bank_is_open_3),
	.out_cmd_can_activate_4(out_cmd_can_activate_4),
	.out_cmd_bank_is_open_4(out_cmd_bank_is_open_4),
	.out_cmd_can_activate_1(out_cmd_can_activate_1),
	.out_cmd_bank_is_open_1(out_cmd_bank_is_open_1),
	.Mux10(\bank_timer_inst|Mux10~2_combout ),
	.Mux13(\bank_timer_inst|Mux13~2_combout ),
	.always106(\bank_timer_inst|always106~0_combout ),
	.always145(\bypass_inst|always145~0_combout ),
	.act_cmd_monitor_per_chip0act_cmd_cnt1(\rank_monitor_inst|act_cmd_monitor_per_chip[0].act_cmd_cnt[1]~q ),
	.act_cmd_monitor_per_chip0act_cmd_cnt2(\rank_monitor_inst|act_cmd_monitor_per_chip[0].act_cmd_cnt[2]~q ),
	.Mux1(\bank_timer_inst|Mux1~2_combout ),
	.can_al_activate_write(\bank_timer_inst|can_al_activate_write~0_combout ),
	.Mux12(\bank_timer_inst|Mux12~0_combout ),
	.rdwr_ready(\bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[0].bank_timer_info_inst|rdwr_ready~q ),
	.rdwr_ready1(\bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[4].bank_timer_info_inst|rdwr_ready~q ),
	.rdwr_ready2(\bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[2].bank_timer_info_inst|rdwr_ready~q ),
	.rdwr_ready3(\bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[6].bank_timer_info_inst|rdwr_ready~q ),
	.Mux9(\bank_timer_inst|Mux9~0_combout ),
	.can_al_activate_read(\bank_timer_inst|can_al_activate_read~0_combout ),
	.pipefull_4(pipefull_4),
	.cs_all_banks_closed_0(\bank_timer_inst|cs_all_banks_closed[0]~q ),
	.always140(\bypass_inst|always140~0_combout ),
	.pipefull_2(pipefull_2),
	.Mux16(\bank_timer_inst|Mux16~2_combout ),
	.Mux19(\bank_timer_inst|Mux19~2_combout ),
	.Mux3(\bank_timer_inst|Mux3~2_combout ),
	.Mux2(\bank_timer_inst|Mux2~2_combout ),
	.pipefull_3(pipefull_3),
	.Mux22(\bank_timer_inst|Mux22~2_combout ),
	.Mux4(\bank_timer_inst|Mux4~2_combout ),
	.always71(\bypass_inst|always71~0_combout ),
	.GND_port(GND_port));

ddr3_int_alt_ddrx_timing_param timing_param_inst(
	.clk_0(clk_0),
	.add_lat_on1(add_lat_on),
	.act_to_rdwr_1(\timing_param_inst|act_to_rdwr[1]~q ),
	.reset_reg_12(reset_reg_12),
	.more_than_3_wr_to_pch1(\timing_param_inst|more_than_3_wr_to_pch~q ));

ddr3_int_alt_ddrx_bank_timer bank_timer_inst(
	.clk_0(clk_0),
	.do_read_r(do_read_r),
	.do_auto_precharge_r(do_auto_precharge_r),
	.do_write_r(do_write_r),
	.pipe_10_0(pipe_10_0),
	.pipe_12_0(pipe_12_0),
	.pipe_11_0(pipe_11_0),
	.Mux0(\bank_timer_inst|Mux0~4_combout ),
	.write_dqs_ready(\rank_monitor_inst|write_dqs_ready~q ),
	.pipe_12_2(pipe_12_2),
	.pipe_12_3(pipe_12_3),
	.pipe_12_1(pipe_12_1),
	.pipe_10_2(pipe_10_2),
	.pipe_10_3(pipe_10_3),
	.pipe_10_1(pipe_10_1),
	.pipe_11_2(pipe_11_2),
	.pipe_11_3(pipe_11_3),
	.pipe_11_1(pipe_11_1),
	.read_dqs_ready(\rank_monitor_inst|read_dqs_ready~q ),
	.pipe_12_4(pipe_12_4),
	.pipe_11_4(pipe_11_4),
	.pipe_10_4(pipe_10_4),
	.Mux25(\bank_timer_inst|Mux25~4_combout ),
	.Mux5(\bank_timer_inst|Mux5~4_combout ),
	.do_precharge_all_r(do_precharge_all_r),
	.can_al_activate_write1(can_al_activate_write),
	.to_chip_r_0(to_chip_r_0),
	.always38(always38),
	.to_bank_addr_r_2(to_bank_addr_r_2),
	.current_bank_2(current_bank_2),
	.to_bank_addr_r_0(to_bank_addr_r_0),
	.current_bank_0(current_bank_0),
	.to_bank_addr_r_1(to_bank_addr_r_1),
	.current_bank_1(current_bank_1),
	.can_al_activate_read1(can_al_activate_read),
	.do_activate_r(do_activate_r),
	.act_ready(\bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[7].bank_timer_info_inst|act_ready~combout ),
	.act_ready1(\bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[5].bank_timer_info_inst|act_ready~combout ),
	.act_ready2(\bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[6].bank_timer_info_inst|act_ready~combout ),
	.act_ready3(\bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[1].bank_timer_info_inst|act_ready~combout ),
	.act_ready4(\bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[0].bank_timer_info_inst|act_ready~combout ),
	.act_ready5(\bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[4].bank_timer_info_inst|act_ready~combout ),
	.act_ready6(\bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[2].bank_timer_info_inst|act_ready~combout ),
	.act_ready7(\bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[3].bank_timer_info_inst|act_ready~combout ),
	.act_to_rdwr_1(\timing_param_inst|act_to_rdwr[1]~q ),
	.Mux10(\bank_timer_inst|Mux10~2_combout ),
	.Mux13(\bank_timer_inst|Mux13~2_combout ),
	.always106(\bank_timer_inst|always106~0_combout ),
	.always145(\bypass_inst|always145~0_combout ),
	.Mux1(\bank_timer_inst|Mux1~2_combout ),
	.more_than_3_wr_to_pch(\timing_param_inst|more_than_3_wr_to_pch~q ),
	.can_al_activate_write2(\bank_timer_inst|can_al_activate_write~0_combout ),
	.reset_reg_8(reset_reg_8),
	.Mux12(\bank_timer_inst|Mux12~0_combout ),
	.rdwr_ready(\bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[0].bank_timer_info_inst|rdwr_ready~q ),
	.rdwr_ready1(\bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[4].bank_timer_info_inst|rdwr_ready~q ),
	.rdwr_ready2(\bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[2].bank_timer_info_inst|rdwr_ready~q ),
	.rdwr_ready3(\bank_timer_inst|bank_timer_info_per_chip[0].bank_timer_info_per_bank[6].bank_timer_info_inst|rdwr_ready~q ),
	.Mux9(\bank_timer_inst|Mux9~0_combout ),
	.write_to_read_finish_twtr_0(\rank_monitor_inst|write_to_read_finish_twtr[0]~q ),
	.can_al_activate_read2(\bank_timer_inst|can_al_activate_read~0_combout ),
	.cs_all_banks_closed_0(\bank_timer_inst|cs_all_banks_closed[0]~q ),
	.always140(\bypass_inst|always140~0_combout ),
	.Mux16(\bank_timer_inst|Mux16~2_combout ),
	.Mux19(\bank_timer_inst|Mux19~2_combout ),
	.Mux3(\bank_timer_inst|Mux3~2_combout ),
	.Mux2(\bank_timer_inst|Mux2~2_combout ),
	.Mux22(\bank_timer_inst|Mux22~2_combout ),
	.Mux4(\bank_timer_inst|Mux4~2_combout ),
	.always1(always1),
	.GND_port(GND_port));

endmodule

module ddr3_int_alt_ddrx_bank_timer (
	clk_0,
	do_read_r,
	do_auto_precharge_r,
	do_write_r,
	pipe_10_0,
	pipe_12_0,
	pipe_11_0,
	Mux0,
	write_dqs_ready,
	pipe_12_2,
	pipe_12_3,
	pipe_12_1,
	pipe_10_2,
	pipe_10_3,
	pipe_10_1,
	pipe_11_2,
	pipe_11_3,
	pipe_11_1,
	read_dqs_ready,
	pipe_12_4,
	pipe_11_4,
	pipe_10_4,
	Mux25,
	Mux5,
	do_precharge_all_r,
	can_al_activate_write1,
	to_chip_r_0,
	always38,
	to_bank_addr_r_2,
	current_bank_2,
	to_bank_addr_r_0,
	current_bank_0,
	to_bank_addr_r_1,
	current_bank_1,
	can_al_activate_read1,
	do_activate_r,
	act_ready,
	act_ready1,
	act_ready2,
	act_ready3,
	act_ready4,
	act_ready5,
	act_ready6,
	act_ready7,
	act_to_rdwr_1,
	Mux10,
	Mux13,
	always106,
	always145,
	Mux1,
	more_than_3_wr_to_pch,
	can_al_activate_write2,
	reset_reg_8,
	Mux12,
	rdwr_ready,
	rdwr_ready1,
	rdwr_ready2,
	rdwr_ready3,
	Mux9,
	write_to_read_finish_twtr_0,
	can_al_activate_read2,
	cs_all_banks_closed_0,
	always140,
	Mux16,
	Mux19,
	Mux3,
	Mux2,
	Mux22,
	Mux4,
	always1,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	clk_0;
input 	do_read_r;
input 	do_auto_precharge_r;
input 	do_write_r;
input 	pipe_10_0;
input 	pipe_12_0;
input 	pipe_11_0;
output 	Mux0;
input 	write_dqs_ready;
input 	pipe_12_2;
input 	pipe_12_3;
input 	pipe_12_1;
input 	pipe_10_2;
input 	pipe_10_3;
input 	pipe_10_1;
input 	pipe_11_2;
input 	pipe_11_3;
input 	pipe_11_1;
input 	read_dqs_ready;
input 	pipe_12_4;
input 	pipe_11_4;
input 	pipe_10_4;
output 	Mux25;
output 	Mux5;
input 	do_precharge_all_r;
output 	can_al_activate_write1;
input 	to_chip_r_0;
input 	always38;
input 	to_bank_addr_r_2;
input 	current_bank_2;
input 	to_bank_addr_r_0;
input 	current_bank_0;
input 	to_bank_addr_r_1;
input 	current_bank_1;
output 	can_al_activate_read1;
input 	do_activate_r;
output 	act_ready;
output 	act_ready1;
output 	act_ready2;
output 	act_ready3;
output 	act_ready4;
output 	act_ready5;
output 	act_ready6;
output 	act_ready7;
input 	act_to_rdwr_1;
output 	Mux10;
output 	Mux13;
output 	always106;
input 	always145;
output 	Mux1;
input 	more_than_3_wr_to_pch;
output 	can_al_activate_write2;
input 	reset_reg_8;
output 	Mux12;
output 	rdwr_ready;
output 	rdwr_ready1;
output 	rdwr_ready2;
output 	rdwr_ready3;
output 	Mux9;
input 	write_to_read_finish_twtr_0;
output 	can_al_activate_read2;
output 	cs_all_banks_closed_0;
input 	always140;
output 	Mux16;
output 	Mux19;
output 	Mux3;
output 	Mux2;
output 	Mux22;
output 	Mux4;
output 	always1;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \bank_timer_info_per_chip[0].bank_timer_info_per_bank[5].bank_timer_info_inst|current_state~q ;
wire \bank_timer_info_per_chip[0].bank_timer_info_per_bank[7].bank_timer_info_inst|current_state~q ;
wire \bank_timer_info_per_chip[0].bank_timer_info_per_bank[4].bank_timer_info_inst|current_state~q ;
wire \bank_timer_info_per_chip[0].bank_timer_info_per_bank[1].bank_timer_info_inst|current_state~q ;
wire \bank_timer_info_per_chip[0].bank_timer_info_per_bank[3].bank_timer_info_inst|current_state~q ;
wire \bank_timer_info_per_chip[0].bank_timer_info_per_bank[0].bank_timer_info_inst|current_state~q ;
wire \bank_timer_info_per_chip[0].bank_timer_info_per_bank[2].bank_timer_info_inst|current_state~q ;
wire \bank_timer_info_per_chip[0].bank_timer_info_per_bank[6].bank_timer_info_inst|current_state~q ;
wire \bank_timer_info_per_chip[0].bank_timer_info_per_bank[1].bank_timer_info_inst|rdwr_ready~q ;
wire \bank_timer_info_per_chip[0].bank_timer_info_per_bank[5].bank_timer_info_inst|rdwr_ready~q ;
wire \bank_timer_info_per_chip[0].bank_timer_info_per_bank[3].bank_timer_info_inst|rdwr_ready~q ;
wire \bank_timer_info_per_chip[0].bank_timer_info_per_bank[7].bank_timer_info_inst|rdwr_ready~q ;
wire \Equal0~0_combout ;
wire \close[0][7]~combout ;
wire \open[0][7]~combout ;
wire \Equal0~1_combout ;
wire \close[0][5]~combout ;
wire \open[0][5]~combout ;
wire \Equal0~2_combout ;
wire \close[0][6]~combout ;
wire \open[0][6]~combout ;
wire \Equal0~3_combout ;
wire \close[0][1]~combout ;
wire \open[0][1]~combout ;
wire \Equal0~4_combout ;
wire \close[0][0]~combout ;
wire \open[0][0]~combout ;
wire \Equal0~5_combout ;
wire \close[0][4]~combout ;
wire \open[0][4]~combout ;
wire \Equal0~6_combout ;
wire \close[0][2]~combout ;
wire \open[0][2]~combout ;
wire \Equal0~7_combout ;
wire \close[0][3]~combout ;
wire \open[0][3]~combout ;
wire \bank_timer_info_per_chip[0].bank_timer_info_per_bank[0].bank_timer_info_inst|general_counter~0_combout ;
wire \Mux0~0_combout ;
wire \Mux25~0_combout ;
wire \Mux5~0_combout ;
wire \Mux10~0_combout ;
wire \Mux10~1_combout ;
wire \Mux13~0_combout ;
wire \Mux13~1_combout ;
wire \Mux1~0_combout ;
wire \Mux1~1_combout ;
wire \WideOr0~0_combout ;
wire \WideOr0~combout ;
wire \Mux16~0_combout ;
wire \Mux16~1_combout ;
wire \Mux19~0_combout ;
wire \Mux19~1_combout ;
wire \Mux3~0_combout ;
wire \Mux3~1_combout ;
wire \Mux2~0_combout ;
wire \Mux2~1_combout ;
wire \Mux22~0_combout ;
wire \Mux22~1_combout ;
wire \Mux4~0_combout ;
wire \Mux4~1_combout ;


ddr3_int_alt_ddrx_bank_timer_info_1 \bank_timer_info_per_chip[0].bank_timer_info_per_bank[1].bank_timer_info_inst (
	.ctl_clk(clk_0),
	.do_read_r(do_read_r),
	.do_write_r(do_write_r),
	.current_state1(\bank_timer_info_per_chip[0].bank_timer_info_per_bank[1].bank_timer_info_inst|current_state~q ),
	.do_precharge_all_r(do_precharge_all_r),
	.to_chip_r_0(to_chip_r_0),
	.always38(always38),
	.act_ready1(act_ready3),
	.act_to_rdwr_1(act_to_rdwr_1),
	.always106(always106),
	.always145(always145),
	.ctl_reset_n(reset_reg_8),
	.rdwr_ready1(\bank_timer_info_per_chip[0].bank_timer_info_per_bank[1].bank_timer_info_inst|rdwr_ready~q ),
	.always140(always140),
	.Equal0(\Equal0~3_combout ),
	.close_1_0(\close[0][1]~combout ),
	.open_1_0(\open[0][1]~combout ),
	.general_counter(\bank_timer_info_per_chip[0].bank_timer_info_per_bank[0].bank_timer_info_inst|general_counter~0_combout ),
	.GND_port(GND_port));

ddr3_int_alt_ddrx_bank_timer_info_2 \bank_timer_info_per_chip[0].bank_timer_info_per_bank[2].bank_timer_info_inst (
	.ctl_clk(clk_0),
	.do_read_r(do_read_r),
	.do_write_r(do_write_r),
	.current_state1(\bank_timer_info_per_chip[0].bank_timer_info_per_bank[2].bank_timer_info_inst|current_state~q ),
	.do_precharge_all_r(do_precharge_all_r),
	.to_chip_r_0(to_chip_r_0),
	.always38(always38),
	.act_ready1(act_ready6),
	.act_to_rdwr_1(act_to_rdwr_1),
	.always106(always106),
	.always145(always145),
	.ctl_reset_n(reset_reg_8),
	.rdwr_ready1(rdwr_ready2),
	.always140(always140),
	.Equal0(\Equal0~6_combout ),
	.close_2_0(\close[0][2]~combout ),
	.open_2_0(\open[0][2]~combout ),
	.general_counter(\bank_timer_info_per_chip[0].bank_timer_info_per_bank[0].bank_timer_info_inst|general_counter~0_combout ),
	.always1(always1),
	.GND_port(GND_port));

ddr3_int_alt_ddrx_bank_timer_info_3 \bank_timer_info_per_chip[0].bank_timer_info_per_bank[3].bank_timer_info_inst (
	.ctl_clk(clk_0),
	.do_read_r(do_read_r),
	.do_write_r(do_write_r),
	.current_state1(\bank_timer_info_per_chip[0].bank_timer_info_per_bank[3].bank_timer_info_inst|current_state~q ),
	.do_precharge_all_r(do_precharge_all_r),
	.to_chip_r_0(to_chip_r_0),
	.always38(always38),
	.act_ready1(act_ready7),
	.act_to_rdwr_1(act_to_rdwr_1),
	.always106(always106),
	.always145(always145),
	.ctl_reset_n(reset_reg_8),
	.rdwr_ready1(\bank_timer_info_per_chip[0].bank_timer_info_per_bank[3].bank_timer_info_inst|rdwr_ready~q ),
	.always140(always140),
	.Equal0(\Equal0~7_combout ),
	.close_3_0(\close[0][3]~combout ),
	.open_3_0(\open[0][3]~combout ),
	.general_counter(\bank_timer_info_per_chip[0].bank_timer_info_per_bank[0].bank_timer_info_inst|general_counter~0_combout ),
	.GND_port(GND_port));

ddr3_int_alt_ddrx_bank_timer_info_4 \bank_timer_info_per_chip[0].bank_timer_info_per_bank[4].bank_timer_info_inst (
	.ctl_clk(clk_0),
	.do_read_r(do_read_r),
	.do_write_r(do_write_r),
	.current_state1(\bank_timer_info_per_chip[0].bank_timer_info_per_bank[4].bank_timer_info_inst|current_state~q ),
	.do_precharge_all_r(do_precharge_all_r),
	.to_chip_r_0(to_chip_r_0),
	.always38(always38),
	.act_ready1(act_ready5),
	.act_to_rdwr_1(act_to_rdwr_1),
	.always106(always106),
	.always145(always145),
	.ctl_reset_n(reset_reg_8),
	.rdwr_ready1(rdwr_ready1),
	.always140(always140),
	.Equal0(\Equal0~5_combout ),
	.close_4_0(\close[0][4]~combout ),
	.open_4_0(\open[0][4]~combout ),
	.general_counter(\bank_timer_info_per_chip[0].bank_timer_info_per_bank[0].bank_timer_info_inst|general_counter~0_combout ),
	.GND_port(GND_port));

ddr3_int_alt_ddrx_bank_timer_info_5 \bank_timer_info_per_chip[0].bank_timer_info_per_bank[5].bank_timer_info_inst (
	.ctl_clk(clk_0),
	.do_read_r(do_read_r),
	.do_write_r(do_write_r),
	.current_state1(\bank_timer_info_per_chip[0].bank_timer_info_per_bank[5].bank_timer_info_inst|current_state~q ),
	.do_precharge_all_r(do_precharge_all_r),
	.to_chip_r_0(to_chip_r_0),
	.always38(always38),
	.act_ready1(act_ready1),
	.act_to_rdwr_1(act_to_rdwr_1),
	.always106(always106),
	.always145(always145),
	.ctl_reset_n(reset_reg_8),
	.rdwr_ready1(\bank_timer_info_per_chip[0].bank_timer_info_per_bank[5].bank_timer_info_inst|rdwr_ready~q ),
	.always140(always140),
	.Equal0(\Equal0~1_combout ),
	.close_5_0(\close[0][5]~combout ),
	.open_5_0(\open[0][5]~combout ),
	.general_counter(\bank_timer_info_per_chip[0].bank_timer_info_per_bank[0].bank_timer_info_inst|general_counter~0_combout ),
	.GND_port(GND_port));

ddr3_int_alt_ddrx_bank_timer_info_6 \bank_timer_info_per_chip[0].bank_timer_info_per_bank[6].bank_timer_info_inst (
	.ctl_clk(clk_0),
	.do_read_r(do_read_r),
	.do_write_r(do_write_r),
	.current_state1(\bank_timer_info_per_chip[0].bank_timer_info_per_bank[6].bank_timer_info_inst|current_state~q ),
	.do_precharge_all_r(do_precharge_all_r),
	.to_chip_r_0(to_chip_r_0),
	.always38(always38),
	.act_ready1(act_ready2),
	.act_to_rdwr_1(act_to_rdwr_1),
	.always106(always106),
	.always145(always145),
	.ctl_reset_n(reset_reg_8),
	.rdwr_ready1(rdwr_ready3),
	.always140(always140),
	.Equal0(\Equal0~2_combout ),
	.close_6_0(\close[0][6]~combout ),
	.open_6_0(\open[0][6]~combout ),
	.general_counter(\bank_timer_info_per_chip[0].bank_timer_info_per_bank[0].bank_timer_info_inst|general_counter~0_combout ),
	.GND_port(GND_port));

ddr3_int_alt_ddrx_bank_timer_info_7 \bank_timer_info_per_chip[0].bank_timer_info_per_bank[7].bank_timer_info_inst (
	.ctl_clk(clk_0),
	.do_read_r(do_read_r),
	.do_write_r(do_write_r),
	.current_state1(\bank_timer_info_per_chip[0].bank_timer_info_per_bank[7].bank_timer_info_inst|current_state~q ),
	.do_precharge_all_r(do_precharge_all_r),
	.to_chip_r_0(to_chip_r_0),
	.always38(always38),
	.act_ready1(act_ready),
	.act_to_rdwr_1(act_to_rdwr_1),
	.always106(always106),
	.always145(always145),
	.ctl_reset_n(reset_reg_8),
	.rdwr_ready1(\bank_timer_info_per_chip[0].bank_timer_info_per_bank[7].bank_timer_info_inst|rdwr_ready~q ),
	.always140(always140),
	.Equal0(\Equal0~0_combout ),
	.close_7_0(\close[0][7]~combout ),
	.open_7_0(\open[0][7]~combout ),
	.general_counter(\bank_timer_info_per_chip[0].bank_timer_info_per_bank[0].bank_timer_info_inst|general_counter~0_combout ),
	.GND_port(GND_port));

ddr3_int_alt_ddrx_bank_timer_info \bank_timer_info_per_chip[0].bank_timer_info_per_bank[0].bank_timer_info_inst (
	.ctl_clk(clk_0),
	.do_read_r(do_read_r),
	.do_auto_precharge_r(do_auto_precharge_r),
	.do_write_r(do_write_r),
	.current_state1(\bank_timer_info_per_chip[0].bank_timer_info_per_bank[0].bank_timer_info_inst|current_state~q ),
	.do_precharge_all_r(do_precharge_all_r),
	.to_chip_r_0(to_chip_r_0),
	.always38(always38),
	.act_ready1(act_ready4),
	.act_to_rdwr_1(act_to_rdwr_1),
	.always106(always106),
	.always145(always145),
	.ctl_reset_n(reset_reg_8),
	.rdwr_ready1(rdwr_ready),
	.always140(always140),
	.Equal0(\Equal0~4_combout ),
	.close_0_0(\close[0][0]~combout ),
	.open_0_0(\open[0][0]~combout ),
	.general_counter(\bank_timer_info_per_chip[0].bank_timer_info_per_bank[0].bank_timer_info_inst|general_counter~0_combout ),
	.GND_port(GND_port));

arriaii_lcell_comb \Equal0~0 (
	.dataa(!to_bank_addr_r_2),
	.datab(!to_bank_addr_r_0),
	.datac(!to_bank_addr_r_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h0101010101010101;
defparam \Equal0~0 .shared_arith = "off";

arriaii_lcell_comb \close[0][7] (
	.dataa(!always38),
	.datab(!always106),
	.datac(!\Equal0~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\close[0][7]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \close[0][7] .extended_lut = "off";
defparam \close[0][7] .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \close[0][7] .shared_arith = "off";

arriaii_lcell_comb \open[0][7] (
	.dataa(!to_chip_r_0),
	.datab(!do_activate_r),
	.datac(!to_bank_addr_r_2),
	.datad(!to_bank_addr_r_0),
	.datae(!to_bank_addr_r_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\open[0][7]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \open[0][7] .extended_lut = "off";
defparam \open[0][7] .lut_mask = 64'h0000000100000001;
defparam \open[0][7] .shared_arith = "off";

arriaii_lcell_comb \Equal0~1 (
	.dataa(!to_bank_addr_r_2),
	.datab(!to_bank_addr_r_0),
	.datac(!to_bank_addr_r_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~1 .extended_lut = "off";
defparam \Equal0~1 .lut_mask = 64'h1010101010101010;
defparam \Equal0~1 .shared_arith = "off";

arriaii_lcell_comb \close[0][5] (
	.dataa(!always38),
	.datab(!always106),
	.datac(!\Equal0~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\close[0][5]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \close[0][5] .extended_lut = "off";
defparam \close[0][5] .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \close[0][5] .shared_arith = "off";

arriaii_lcell_comb \open[0][5] (
	.dataa(!to_chip_r_0),
	.datab(!do_activate_r),
	.datac(!to_bank_addr_r_2),
	.datad(!to_bank_addr_r_0),
	.datae(!to_bank_addr_r_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\open[0][5]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \open[0][5] .extended_lut = "off";
defparam \open[0][5] .lut_mask = 64'h0001000000010000;
defparam \open[0][5] .shared_arith = "off";

arriaii_lcell_comb \Equal0~2 (
	.dataa(!to_bank_addr_r_2),
	.datab(!to_bank_addr_r_0),
	.datac(!to_bank_addr_r_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~2 .extended_lut = "off";
defparam \Equal0~2 .lut_mask = 64'h0404040404040404;
defparam \Equal0~2 .shared_arith = "off";

arriaii_lcell_comb \close[0][6] (
	.dataa(!always38),
	.datab(!always106),
	.datac(!\Equal0~2_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\close[0][6]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \close[0][6] .extended_lut = "off";
defparam \close[0][6] .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \close[0][6] .shared_arith = "off";

arriaii_lcell_comb \open[0][6] (
	.dataa(!to_chip_r_0),
	.datab(!do_activate_r),
	.datac(!to_bank_addr_r_2),
	.datad(!to_bank_addr_r_0),
	.datae(!to_bank_addr_r_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\open[0][6]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \open[0][6] .extended_lut = "off";
defparam \open[0][6] .lut_mask = 64'h0000010000000100;
defparam \open[0][6] .shared_arith = "off";

arriaii_lcell_comb \Equal0~3 (
	.dataa(!to_bank_addr_r_2),
	.datab(!to_bank_addr_r_0),
	.datac(!to_bank_addr_r_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~3 .extended_lut = "off";
defparam \Equal0~3 .lut_mask = 64'h2020202020202020;
defparam \Equal0~3 .shared_arith = "off";

arriaii_lcell_comb \close[0][1] (
	.dataa(!always38),
	.datab(!always106),
	.datac(!\Equal0~3_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\close[0][1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \close[0][1] .extended_lut = "off";
defparam \close[0][1] .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \close[0][1] .shared_arith = "off";

arriaii_lcell_comb \open[0][1] (
	.dataa(!to_chip_r_0),
	.datab(!do_activate_r),
	.datac(!to_bank_addr_r_2),
	.datad(!to_bank_addr_r_0),
	.datae(!to_bank_addr_r_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\open[0][1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \open[0][1] .extended_lut = "off";
defparam \open[0][1] .lut_mask = 64'h0010000000100000;
defparam \open[0][1] .shared_arith = "off";

arriaii_lcell_comb \Equal0~4 (
	.dataa(!to_bank_addr_r_2),
	.datab(!to_bank_addr_r_0),
	.datac(!to_bank_addr_r_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~4 .extended_lut = "off";
defparam \Equal0~4 .lut_mask = 64'h8080808080808080;
defparam \Equal0~4 .shared_arith = "off";

arriaii_lcell_comb \close[0][0] (
	.dataa(!always38),
	.datab(!always106),
	.datac(!\Equal0~4_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\close[0][0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \close[0][0] .extended_lut = "off";
defparam \close[0][0] .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \close[0][0] .shared_arith = "off";

arriaii_lcell_comb \open[0][0] (
	.dataa(!to_chip_r_0),
	.datab(!do_activate_r),
	.datac(!to_bank_addr_r_2),
	.datad(!to_bank_addr_r_0),
	.datae(!to_bank_addr_r_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\open[0][0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \open[0][0] .extended_lut = "off";
defparam \open[0][0] .lut_mask = 64'h1000000010000000;
defparam \open[0][0] .shared_arith = "off";

arriaii_lcell_comb \Equal0~5 (
	.dataa(!to_bank_addr_r_2),
	.datab(!to_bank_addr_r_0),
	.datac(!to_bank_addr_r_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~5 .extended_lut = "off";
defparam \Equal0~5 .lut_mask = 64'h4040404040404040;
defparam \Equal0~5 .shared_arith = "off";

arriaii_lcell_comb \close[0][4] (
	.dataa(!always38),
	.datab(!always106),
	.datac(!\Equal0~5_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\close[0][4]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \close[0][4] .extended_lut = "off";
defparam \close[0][4] .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \close[0][4] .shared_arith = "off";

arriaii_lcell_comb \open[0][4] (
	.dataa(!to_chip_r_0),
	.datab(!do_activate_r),
	.datac(!to_bank_addr_r_2),
	.datad(!to_bank_addr_r_0),
	.datae(!to_bank_addr_r_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\open[0][4]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \open[0][4] .extended_lut = "off";
defparam \open[0][4] .lut_mask = 64'h0100000001000000;
defparam \open[0][4] .shared_arith = "off";

arriaii_lcell_comb \Equal0~6 (
	.dataa(!to_bank_addr_r_2),
	.datab(!to_bank_addr_r_0),
	.datac(!to_bank_addr_r_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~6 .extended_lut = "off";
defparam \Equal0~6 .lut_mask = 64'h0808080808080808;
defparam \Equal0~6 .shared_arith = "off";

arriaii_lcell_comb \close[0][2] (
	.dataa(!always38),
	.datab(!always106),
	.datac(!\Equal0~6_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\close[0][2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \close[0][2] .extended_lut = "off";
defparam \close[0][2] .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \close[0][2] .shared_arith = "off";

arriaii_lcell_comb \open[0][2] (
	.dataa(!to_chip_r_0),
	.datab(!do_activate_r),
	.datac(!to_bank_addr_r_2),
	.datad(!to_bank_addr_r_0),
	.datae(!to_bank_addr_r_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\open[0][2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \open[0][2] .extended_lut = "off";
defparam \open[0][2] .lut_mask = 64'h0000100000001000;
defparam \open[0][2] .shared_arith = "off";

arriaii_lcell_comb \Equal0~7 (
	.dataa(!to_bank_addr_r_2),
	.datab(!to_bank_addr_r_0),
	.datac(!to_bank_addr_r_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~7 .extended_lut = "off";
defparam \Equal0~7 .lut_mask = 64'h0202020202020202;
defparam \Equal0~7 .shared_arith = "off";

arriaii_lcell_comb \close[0][3] (
	.dataa(!always38),
	.datab(!always106),
	.datac(!\Equal0~7_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\close[0][3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \close[0][3] .extended_lut = "off";
defparam \close[0][3] .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \close[0][3] .shared_arith = "off";

arriaii_lcell_comb \open[0][3] (
	.dataa(!to_chip_r_0),
	.datab(!do_activate_r),
	.datac(!to_bank_addr_r_2),
	.datad(!to_bank_addr_r_0),
	.datae(!to_bank_addr_r_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\open[0][3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \open[0][3] .extended_lut = "off";
defparam \open[0][3] .lut_mask = 64'h0000001000000010;
defparam \open[0][3] .shared_arith = "off";

arriaii_lcell_comb \Mux0~4 (
	.dataa(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[5].bank_timer_info_inst|current_state~q ),
	.datab(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[7].bank_timer_info_inst|current_state~q ),
	.datac(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[6].bank_timer_info_inst|current_state~q ),
	.datad(!current_bank_2),
	.datae(!current_bank_1),
	.dataf(!\Mux0~0_combout ),
	.datag(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[4].bank_timer_info_inst|current_state~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux0),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~4 .extended_lut = "on";
defparam \Mux0~4 .lut_mask = 64'h000F000FFF55FF33;
defparam \Mux0~4 .shared_arith = "off";

arriaii_lcell_comb \Mux25~4 (
	.dataa(!act_ready1),
	.datab(!act_ready),
	.datac(!act_ready2),
	.datad(!pipe_12_4),
	.datae(!pipe_11_4),
	.dataf(!\Mux25~0_combout ),
	.datag(!act_ready5),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux25),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux25~4 .extended_lut = "on";
defparam \Mux25~4 .lut_mask = 64'h000F000FFF55FF33;
defparam \Mux25~4 .shared_arith = "off";

arriaii_lcell_comb \Mux5~4 (
	.dataa(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[5].bank_timer_info_inst|current_state~q ),
	.datab(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[7].bank_timer_info_inst|current_state~q ),
	.datac(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[6].bank_timer_info_inst|current_state~q ),
	.datad(!pipe_12_4),
	.datae(!pipe_11_4),
	.dataf(!\Mux5~0_combout ),
	.datag(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[4].bank_timer_info_inst|current_state~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux5),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux5~4 .extended_lut = "on";
defparam \Mux5~4 .lut_mask = 64'h000F000FFF55FF33;
defparam \Mux5~4 .shared_arith = "off";

dffeas can_al_activate_write(
	.clk(clk_0),
	.d(can_al_activate_write2),
	.asdata(vcc),
	.clrn(reset_reg_8),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(can_al_activate_write1),
	.prn(vcc));
defparam can_al_activate_write.is_wysiwyg = "true";
defparam can_al_activate_write.power_up = "low";

dffeas can_al_activate_read(
	.clk(clk_0),
	.d(can_al_activate_read2),
	.asdata(vcc),
	.clrn(reset_reg_8),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(can_al_activate_read1),
	.prn(vcc));
defparam can_al_activate_read.is_wysiwyg = "true";
defparam can_al_activate_read.power_up = "low";

arriaii_lcell_comb \Mux10~2 (
	.dataa(!current_bank_2),
	.datab(!current_bank_0),
	.datac(!current_bank_1),
	.datad(!act_ready6),
	.datae(!\Mux10~0_combout ),
	.dataf(!\Mux10~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux10),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux10~2 .extended_lut = "off";
defparam \Mux10~2 .lut_mask = 64'h0008333BC4CCF7FF;
defparam \Mux10~2 .shared_arith = "off";

arriaii_lcell_comb \Mux13~2 (
	.dataa(!act_ready6),
	.datab(!pipe_10_0),
	.datac(!pipe_12_0),
	.datad(!pipe_11_0),
	.datae(!\Mux13~0_combout ),
	.dataf(!\Mux13~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux13),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux13~2 .extended_lut = "off";
defparam \Mux13~2 .lut_mask = 64'h00403373CC4CFF7F;
defparam \Mux13~2 .shared_arith = "off";

arriaii_lcell_comb \always106~0 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always106),
	.sumout(),
	.cout(),
	.shareout());
defparam \always106~0 .extended_lut = "off";
defparam \always106~0 .lut_mask = 64'h1111111111111111;
defparam \always106~0 .shared_arith = "off";

arriaii_lcell_comb \Mux1~2 (
	.dataa(!pipe_10_0),
	.datab(!\Mux1~0_combout ),
	.datac(!\Mux1~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux1),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~2 .extended_lut = "off";
defparam \Mux1~2 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \Mux1~2 .shared_arith = "off";

arriaii_lcell_comb \can_al_activate_write~0 (
	.dataa(!do_read_r),
	.datab(!more_than_3_wr_to_pch),
	.datac(!write_dqs_ready),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(can_al_activate_write2),
	.sumout(),
	.cout(),
	.shareout());
defparam \can_al_activate_write~0 .extended_lut = "off";
defparam \can_al_activate_write~0 .lut_mask = 64'h0E0E0E0E0E0E0E0E;
defparam \can_al_activate_write~0 .shared_arith = "off";

arriaii_lcell_comb \Mux12~0 (
	.dataa(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[1].bank_timer_info_inst|rdwr_ready~q ),
	.datab(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[5].bank_timer_info_inst|rdwr_ready~q ),
	.datac(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[3].bank_timer_info_inst|rdwr_ready~q ),
	.datad(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[7].bank_timer_info_inst|rdwr_ready~q ),
	.datae(!pipe_12_0),
	.dataf(!pipe_11_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux12),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux12~0 .extended_lut = "off";
defparam \Mux12~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux12~0 .shared_arith = "off";

arriaii_lcell_comb \Mux9~0 (
	.dataa(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[1].bank_timer_info_inst|rdwr_ready~q ),
	.datab(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[5].bank_timer_info_inst|rdwr_ready~q ),
	.datac(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[3].bank_timer_info_inst|rdwr_ready~q ),
	.datad(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[7].bank_timer_info_inst|rdwr_ready~q ),
	.datae(!current_bank_2),
	.dataf(!current_bank_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux9),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux9~0 .extended_lut = "off";
defparam \Mux9~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux9~0 .shared_arith = "off";

arriaii_lcell_comb \can_al_activate_read~0 (
	.dataa(!do_write_r),
	.datab(!more_than_3_wr_to_pch),
	.datac(!write_to_read_finish_twtr_0),
	.datad(!read_dqs_ready),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(can_al_activate_read2),
	.sumout(),
	.cout(),
	.shareout());
defparam \can_al_activate_read~0 .extended_lut = "off";
defparam \can_al_activate_read~0 .lut_mask = 64'h000E000E000E000E;
defparam \can_al_activate_read~0 .shared_arith = "off";

dffeas \cs_all_banks_closed[0] (
	.clk(clk_0),
	.d(\WideOr0~combout ),
	.asdata(vcc),
	.clrn(reset_reg_8),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(cs_all_banks_closed_0),
	.prn(vcc));
defparam \cs_all_banks_closed[0] .is_wysiwyg = "true";
defparam \cs_all_banks_closed[0] .power_up = "low";

arriaii_lcell_comb \Mux16~2 (
	.dataa(!act_ready6),
	.datab(!pipe_12_1),
	.datac(!pipe_10_1),
	.datad(!pipe_11_1),
	.datae(!\Mux16~0_combout ),
	.dataf(!\Mux16~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux16),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux16~2 .extended_lut = "off";
defparam \Mux16~2 .lut_mask = 64'h00400F4FF070FF7F;
defparam \Mux16~2 .shared_arith = "off";

arriaii_lcell_comb \Mux19~2 (
	.dataa(!act_ready6),
	.datab(!pipe_12_2),
	.datac(!pipe_10_2),
	.datad(!pipe_11_2),
	.datae(!\Mux19~0_combout ),
	.dataf(!\Mux19~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux19),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux19~2 .extended_lut = "off";
defparam \Mux19~2 .lut_mask = 64'h00400F4FF070FF7F;
defparam \Mux19~2 .shared_arith = "off";

arriaii_lcell_comb \Mux3~2 (
	.dataa(!pipe_10_2),
	.datab(!\Mux3~0_combout ),
	.datac(!\Mux3~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux3),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux3~2 .extended_lut = "off";
defparam \Mux3~2 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \Mux3~2 .shared_arith = "off";

arriaii_lcell_comb \Mux2~2 (
	.dataa(!pipe_10_1),
	.datab(!\Mux2~0_combout ),
	.datac(!\Mux2~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux2),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux2~2 .extended_lut = "off";
defparam \Mux2~2 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \Mux2~2 .shared_arith = "off";

arriaii_lcell_comb \Mux22~2 (
	.dataa(!act_ready6),
	.datab(!pipe_12_3),
	.datac(!pipe_10_3),
	.datad(!pipe_11_3),
	.datae(!\Mux22~0_combout ),
	.dataf(!\Mux22~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux22),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux22~2 .extended_lut = "off";
defparam \Mux22~2 .lut_mask = 64'h00400F4FF070FF7F;
defparam \Mux22~2 .shared_arith = "off";

arriaii_lcell_comb \Mux4~2 (
	.dataa(!pipe_10_3),
	.datab(!\Mux4~0_combout ),
	.datac(!\Mux4~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Mux4),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux4~2 .extended_lut = "off";
defparam \Mux4~2 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \Mux4~2 .shared_arith = "off";

arriaii_lcell_comb \Mux0~0 (
	.dataa(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[1].bank_timer_info_inst|current_state~q ),
	.datab(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[3].bank_timer_info_inst|current_state~q ),
	.datac(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[2].bank_timer_info_inst|current_state~q ),
	.datad(!current_bank_0),
	.datae(!current_bank_1),
	.dataf(!current_bank_2),
	.datag(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[0].bank_timer_info_inst|current_state~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~0 .extended_lut = "on";
defparam \Mux0~0 .lut_mask = 64'h0F550F3300FF00FF;
defparam \Mux0~0 .shared_arith = "off";

arriaii_lcell_comb \Mux25~0 (
	.dataa(!act_ready3),
	.datab(!act_ready7),
	.datac(!act_ready6),
	.datad(!pipe_10_4),
	.datae(!pipe_11_4),
	.dataf(!pipe_12_4),
	.datag(!act_ready4),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux25~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux25~0 .extended_lut = "on";
defparam \Mux25~0 .lut_mask = 64'h0F550F3300FF00FF;
defparam \Mux25~0 .shared_arith = "off";

arriaii_lcell_comb \Mux5~0 (
	.dataa(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[1].bank_timer_info_inst|current_state~q ),
	.datab(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[3].bank_timer_info_inst|current_state~q ),
	.datac(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[2].bank_timer_info_inst|current_state~q ),
	.datad(!pipe_10_4),
	.datae(!pipe_11_4),
	.dataf(!pipe_12_4),
	.datag(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[0].bank_timer_info_inst|current_state~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux5~0 .extended_lut = "on";
defparam \Mux5~0 .lut_mask = 64'h0F550F3300FF00FF;
defparam \Mux5~0 .shared_arith = "off";

arriaii_lcell_comb \Mux10~0 (
	.dataa(!act_ready3),
	.datab(!act_ready1),
	.datac(!act_ready7),
	.datad(!act_ready),
	.datae(!current_bank_2),
	.dataf(!current_bank_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux10~0 .extended_lut = "off";
defparam \Mux10~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux10~0 .shared_arith = "off";

arriaii_lcell_comb \Mux10~1 (
	.dataa(!current_bank_2),
	.datab(!current_bank_1),
	.datac(!act_ready2),
	.datad(!act_ready4),
	.datae(!act_ready5),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux10~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux10~1 .extended_lut = "off";
defparam \Mux10~1 .lut_mask = 64'h038B47CF038B47CF;
defparam \Mux10~1 .shared_arith = "off";

arriaii_lcell_comb \Mux13~0 (
	.dataa(!act_ready3),
	.datab(!act_ready1),
	.datac(!act_ready7),
	.datad(!act_ready),
	.datae(!pipe_12_0),
	.dataf(!pipe_11_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux13~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux13~0 .extended_lut = "off";
defparam \Mux13~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux13~0 .shared_arith = "off";

arriaii_lcell_comb \Mux13~1 (
	.dataa(!act_ready2),
	.datab(!act_ready4),
	.datac(!act_ready5),
	.datad(!pipe_12_0),
	.datae(!pipe_11_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux13~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux13~1 .extended_lut = "off";
defparam \Mux13~1 .lut_mask = 64'h330F5555330F5555;
defparam \Mux13~1 .shared_arith = "off";

arriaii_lcell_comb \Mux1~0 (
	.dataa(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[1].bank_timer_info_inst|current_state~q ),
	.datab(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[5].bank_timer_info_inst|current_state~q ),
	.datac(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[3].bank_timer_info_inst|current_state~q ),
	.datad(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[7].bank_timer_info_inst|current_state~q ),
	.datae(!pipe_12_0),
	.dataf(!pipe_11_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~0 .extended_lut = "off";
defparam \Mux1~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux1~0 .shared_arith = "off";

arriaii_lcell_comb \Mux1~1 (
	.dataa(!pipe_12_0),
	.datab(!pipe_11_0),
	.datac(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[4].bank_timer_info_inst|current_state~q ),
	.datad(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[0].bank_timer_info_inst|current_state~q ),
	.datae(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[2].bank_timer_info_inst|current_state~q ),
	.dataf(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[6].bank_timer_info_inst|current_state~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~1 .extended_lut = "off";
defparam \Mux1~1 .lut_mask = 64'h048C26AE159D37BF;
defparam \Mux1~1 .shared_arith = "off";

arriaii_lcell_comb \WideOr0~0 (
	.dataa(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[5].bank_timer_info_inst|current_state~q ),
	.datab(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[7].bank_timer_info_inst|current_state~q ),
	.datac(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[4].bank_timer_info_inst|current_state~q ),
	.datad(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[6].bank_timer_info_inst|current_state~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h8000800080008000;
defparam \WideOr0~0 .shared_arith = "off";

arriaii_lcell_comb WideOr0(
	.dataa(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[1].bank_timer_info_inst|current_state~q ),
	.datab(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[3].bank_timer_info_inst|current_state~q ),
	.datac(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[0].bank_timer_info_inst|current_state~q ),
	.datad(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[2].bank_timer_info_inst|current_state~q ),
	.datae(!\WideOr0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr0.extended_lut = "off";
defparam WideOr0.lut_mask = 64'h0000800000008000;
defparam WideOr0.shared_arith = "off";

arriaii_lcell_comb \Mux16~0 (
	.dataa(!act_ready3),
	.datab(!act_ready1),
	.datac(!act_ready7),
	.datad(!act_ready),
	.datae(!pipe_12_1),
	.dataf(!pipe_11_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux16~0 .extended_lut = "off";
defparam \Mux16~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux16~0 .shared_arith = "off";

arriaii_lcell_comb \Mux16~1 (
	.dataa(!act_ready2),
	.datab(!act_ready4),
	.datac(!act_ready5),
	.datad(!pipe_12_1),
	.datae(!pipe_11_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux16~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux16~1 .extended_lut = "off";
defparam \Mux16~1 .lut_mask = 64'h330F5555330F5555;
defparam \Mux16~1 .shared_arith = "off";

arriaii_lcell_comb \Mux19~0 (
	.dataa(!act_ready3),
	.datab(!act_ready1),
	.datac(!act_ready7),
	.datad(!act_ready),
	.datae(!pipe_12_2),
	.dataf(!pipe_11_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux19~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux19~0 .extended_lut = "off";
defparam \Mux19~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux19~0 .shared_arith = "off";

arriaii_lcell_comb \Mux19~1 (
	.dataa(!act_ready2),
	.datab(!act_ready4),
	.datac(!act_ready5),
	.datad(!pipe_12_2),
	.datae(!pipe_11_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux19~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux19~1 .extended_lut = "off";
defparam \Mux19~1 .lut_mask = 64'h330F5555330F5555;
defparam \Mux19~1 .shared_arith = "off";

arriaii_lcell_comb \Mux3~0 (
	.dataa(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[1].bank_timer_info_inst|current_state~q ),
	.datab(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[5].bank_timer_info_inst|current_state~q ),
	.datac(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[3].bank_timer_info_inst|current_state~q ),
	.datad(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[7].bank_timer_info_inst|current_state~q ),
	.datae(!pipe_12_2),
	.dataf(!pipe_11_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux3~0 .extended_lut = "off";
defparam \Mux3~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux3~0 .shared_arith = "off";

arriaii_lcell_comb \Mux3~1 (
	.dataa(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[4].bank_timer_info_inst|current_state~q ),
	.datab(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[0].bank_timer_info_inst|current_state~q ),
	.datac(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[2].bank_timer_info_inst|current_state~q ),
	.datad(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[6].bank_timer_info_inst|current_state~q ),
	.datae(!pipe_12_2),
	.dataf(!pipe_11_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux3~1 .extended_lut = "off";
defparam \Mux3~1 .lut_mask = 64'h333355550F0F00FF;
defparam \Mux3~1 .shared_arith = "off";

arriaii_lcell_comb \Mux2~0 (
	.dataa(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[1].bank_timer_info_inst|current_state~q ),
	.datab(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[5].bank_timer_info_inst|current_state~q ),
	.datac(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[3].bank_timer_info_inst|current_state~q ),
	.datad(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[7].bank_timer_info_inst|current_state~q ),
	.datae(!pipe_12_1),
	.dataf(!pipe_11_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux2~0 .extended_lut = "off";
defparam \Mux2~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux2~0 .shared_arith = "off";

arriaii_lcell_comb \Mux2~1 (
	.dataa(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[4].bank_timer_info_inst|current_state~q ),
	.datab(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[0].bank_timer_info_inst|current_state~q ),
	.datac(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[2].bank_timer_info_inst|current_state~q ),
	.datad(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[6].bank_timer_info_inst|current_state~q ),
	.datae(!pipe_12_1),
	.dataf(!pipe_11_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux2~1 .extended_lut = "off";
defparam \Mux2~1 .lut_mask = 64'h333355550F0F00FF;
defparam \Mux2~1 .shared_arith = "off";

arriaii_lcell_comb \Mux22~0 (
	.dataa(!act_ready3),
	.datab(!act_ready1),
	.datac(!act_ready7),
	.datad(!act_ready),
	.datae(!pipe_12_3),
	.dataf(!pipe_11_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux22~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux22~0 .extended_lut = "off";
defparam \Mux22~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux22~0 .shared_arith = "off";

arriaii_lcell_comb \Mux22~1 (
	.dataa(!act_ready2),
	.datab(!act_ready4),
	.datac(!act_ready5),
	.datad(!pipe_12_3),
	.datae(!pipe_11_3),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux22~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux22~1 .extended_lut = "off";
defparam \Mux22~1 .lut_mask = 64'h330F5555330F5555;
defparam \Mux22~1 .shared_arith = "off";

arriaii_lcell_comb \Mux4~0 (
	.dataa(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[1].bank_timer_info_inst|current_state~q ),
	.datab(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[5].bank_timer_info_inst|current_state~q ),
	.datac(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[3].bank_timer_info_inst|current_state~q ),
	.datad(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[7].bank_timer_info_inst|current_state~q ),
	.datae(!pipe_12_3),
	.dataf(!pipe_11_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux4~0 .extended_lut = "off";
defparam \Mux4~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux4~0 .shared_arith = "off";

arriaii_lcell_comb \Mux4~1 (
	.dataa(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[4].bank_timer_info_inst|current_state~q ),
	.datab(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[0].bank_timer_info_inst|current_state~q ),
	.datac(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[2].bank_timer_info_inst|current_state~q ),
	.datad(!\bank_timer_info_per_chip[0].bank_timer_info_per_bank[6].bank_timer_info_inst|current_state~q ),
	.datae(!pipe_12_3),
	.dataf(!pipe_11_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux4~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux4~1 .extended_lut = "off";
defparam \Mux4~1 .lut_mask = 64'h333355550F0F00FF;
defparam \Mux4~1 .shared_arith = "off";

endmodule

module ddr3_int_alt_ddrx_bank_timer_info (
	ctl_clk,
	do_read_r,
	do_auto_precharge_r,
	do_write_r,
	current_state1,
	do_precharge_all_r,
	to_chip_r_0,
	always38,
	act_ready1,
	act_to_rdwr_1,
	always106,
	always145,
	ctl_reset_n,
	rdwr_ready1,
	always140,
	Equal0,
	close_0_0,
	open_0_0,
	general_counter,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	ctl_clk;
input 	do_read_r;
input 	do_auto_precharge_r;
input 	do_write_r;
output 	current_state1;
input 	do_precharge_all_r;
input 	to_chip_r_0;
input 	always38;
output 	act_ready1;
input 	act_to_rdwr_1;
input 	always106;
input 	always145;
input 	ctl_reset_n;
output 	rdwr_ready1;
input 	always140;
input 	Equal0;
input 	close_0_0;
input 	open_0_0;
output 	general_counter;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \current_state~0_combout ;
wire \Add1~1_sumout ;
wire \general_counter~2_combout ;
wire \general_counter[0]~q ;
wire \Add1~10 ;
wire \Add1~13_sumout ;
wire \general_counter~4_combout ;
wire \general_counter[3]~q ;
wire \Add1~14 ;
wire \Add1~17_sumout ;
wire \general_counter~6_combout ;
wire \general_counter[4]~q ;
wire \Add1~18 ;
wire \Add1~21_sumout ;
wire \general_counter~5_combout ;
wire \general_counter[5]~q ;
wire \Equal1~0_combout ;
wire \Add1~2 ;
wire \Add1~5_sumout ;
wire \general_counter~3_combout ;
wire \general_counter[1]~q ;
wire \Add1~6 ;
wire \Add1~9_sumout ;
wire \general_counter~1_combout ;
wire \general_counter[2]~q ;
wire \doing_auto_precharge~0_combout ;
wire \doing_precharge~0_combout ;
wire \doing_auto_precharge~q ;
wire \doing_precharge~1_combout ;
wire \doing_precharge~q ;
wire \int_rdwr_to_valid_ready~0_combout ;
wire \int_rdwr_to_valid_ready~1_combout ;
wire \doing_read~0_combout ;
wire \doing_read~q ;
wire \int_rdwr_to_valid_ready~2_combout ;
wire \int_rdwr_to_valid_ready~3_combout ;
wire \int_rdwr_to_valid_ready~q ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \act_counter[4]~q ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \act_counter[5]~q ;
wire \Add0~1_sumout ;
wire \act_counter[0]~q ;
wire \Equal0~0_combout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \act_counter[1]~q ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \act_counter[2]~q ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \act_counter[3]~q ;
wire \LessThan0~0_combout ;
wire \int_act_to_act_ready~q ;
wire \rdwr_ready~0_combout ;
wire \rdwr_ready~1_combout ;


dffeas current_state(
	.clk(ctl_clk),
	.d(\current_state~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_0_0),
	.ena(vcc),
	.q(current_state1),
	.prn(vcc));
defparam current_state.is_wysiwyg = "true";
defparam current_state.power_up = "low";

arriaii_lcell_comb act_ready(
	.dataa(!\int_rdwr_to_valid_ready~q ),
	.datab(!\int_act_to_act_ready~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(act_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam act_ready.extended_lut = "off";
defparam act_ready.lut_mask = 64'h4444444444444444;
defparam act_ready.shared_arith = "off";

dffeas rdwr_ready(
	.clk(ctl_clk),
	.d(\rdwr_ready~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rdwr_ready1),
	.prn(vcc));
defparam rdwr_ready.is_wysiwyg = "true";
defparam rdwr_ready.power_up = "low";

arriaii_lcell_comb \general_counter~0 (
	.dataa(!do_read_r),
	.datab(!do_auto_precharge_r),
	.datac(!do_write_r),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(general_counter),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~0 .extended_lut = "off";
defparam \general_counter~0 .lut_mask = 64'h8080808080808080;
defparam \general_counter~0 .shared_arith = "off";

arriaii_lcell_comb \current_state~0 (
	.dataa(!always38),
	.datab(!always106),
	.datac(!current_state1),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\current_state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \current_state~0 .extended_lut = "off";
defparam \current_state~0 .lut_mask = 64'h0C080C080C080C08;
defparam \current_state~0 .shared_arith = "off";

arriaii_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Equal1~0_combout ),
	.datae(gnd),
	.dataf(!\general_counter[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(\Add1~2 ),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h0000FF000000FF00;
defparam \Add1~1 .shared_arith = "off";

arriaii_lcell_comb \general_counter~2 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~1_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~2 .extended_lut = "off";
defparam \general_counter~2 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~2 .shared_arith = "off";

dffeas \general_counter[0] (
	.clk(ctl_clk),
	.d(\general_counter~2_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[0]~q ),
	.prn(vcc));
defparam \general_counter[0] .is_wysiwyg = "true";
defparam \general_counter[0] .power_up = "low";

arriaii_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~9 .shared_arith = "off";

arriaii_lcell_comb \Add1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~13 .shared_arith = "off";

arriaii_lcell_comb \general_counter~4 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~13_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~4 .extended_lut = "off";
defparam \general_counter~4 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~4 .shared_arith = "off";

dffeas \general_counter[3] (
	.clk(ctl_clk),
	.d(\general_counter~4_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[3]~q ),
	.prn(vcc));
defparam \general_counter[3] .is_wysiwyg = "true";
defparam \general_counter[3] .power_up = "low";

arriaii_lcell_comb \Add1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~17 .shared_arith = "off";

arriaii_lcell_comb \general_counter~6 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~17_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~6 .extended_lut = "off";
defparam \general_counter~6 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~6 .shared_arith = "off";

dffeas \general_counter[4] (
	.clk(ctl_clk),
	.d(\general_counter~6_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[4]~q ),
	.prn(vcc));
defparam \general_counter[4] .is_wysiwyg = "true";
defparam \general_counter[4] .power_up = "low";

arriaii_lcell_comb \Add1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~21_sumout ),
	.cout(),
	.shareout());
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~21 .shared_arith = "off";

arriaii_lcell_comb \general_counter~5 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~21_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~5 .extended_lut = "off";
defparam \general_counter~5 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~5 .shared_arith = "off";

dffeas \general_counter[5] (
	.clk(ctl_clk),
	.d(\general_counter~5_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[5]~q ),
	.prn(vcc));
defparam \general_counter[5] .is_wysiwyg = "true";
defparam \general_counter[5] .power_up = "low";

arriaii_lcell_comb \Equal1~0 (
	.dataa(!\general_counter[2]~q ),
	.datab(!\general_counter[0]~q ),
	.datac(!\general_counter[1]~q ),
	.datad(!\general_counter[3]~q ),
	.datae(!\general_counter[5]~q ),
	.dataf(!\general_counter[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'h0000000000000001;
defparam \Equal1~0 .shared_arith = "off";

arriaii_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~5 .shared_arith = "off";

arriaii_lcell_comb \general_counter~3 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~5_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~3 .extended_lut = "off";
defparam \general_counter~3 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~3 .shared_arith = "off";

dffeas \general_counter[1] (
	.clk(ctl_clk),
	.d(\general_counter~3_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[1]~q ),
	.prn(vcc));
defparam \general_counter[1] .is_wysiwyg = "true";
defparam \general_counter[1] .power_up = "low";

arriaii_lcell_comb \general_counter~1 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~9_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~1 .extended_lut = "off";
defparam \general_counter~1 .lut_mask = 64'h1311FFFF1311FFFF;
defparam \general_counter~1 .shared_arith = "off";

dffeas \general_counter[2] (
	.clk(ctl_clk),
	.d(\general_counter~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[2]~q ),
	.prn(vcc));
defparam \general_counter[2] .is_wysiwyg = "true";
defparam \general_counter[2] .power_up = "low";

arriaii_lcell_comb \doing_auto_precharge~0 (
	.dataa(!always38),
	.datab(!always106),
	.datac(!always140),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_auto_precharge~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_auto_precharge~0 .extended_lut = "off";
defparam \doing_auto_precharge~0 .lut_mask = 64'h0007000700070007;
defparam \doing_auto_precharge~0 .shared_arith = "off";

arriaii_lcell_comb \doing_precharge~0 (
	.dataa(!always38),
	.datab(!always145),
	.datac(!always106),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_precharge~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_precharge~0 .extended_lut = "off";
defparam \doing_precharge~0 .lut_mask = 64'h0F7F0F7F0F7F0F7F;
defparam \doing_precharge~0 .shared_arith = "off";

dffeas doing_auto_precharge(
	.clk(ctl_clk),
	.d(\doing_auto_precharge~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\doing_precharge~0_combout ),
	.q(\doing_auto_precharge~q ),
	.prn(vcc));
defparam doing_auto_precharge.is_wysiwyg = "true";
defparam doing_auto_precharge.power_up = "low";

arriaii_lcell_comb \doing_precharge~1 (
	.dataa(!always38),
	.datab(!always106),
	.datac(!always140),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_precharge~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_precharge~1 .extended_lut = "off";
defparam \doing_precharge~1 .lut_mask = 64'h3370337033703370;
defparam \doing_precharge~1 .shared_arith = "off";

dffeas doing_precharge(
	.clk(ctl_clk),
	.d(\doing_precharge~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\doing_precharge~0_combout ),
	.q(\doing_precharge~q ),
	.prn(vcc));
defparam doing_precharge.is_wysiwyg = "true";
defparam doing_precharge.power_up = "low";

arriaii_lcell_comb \int_rdwr_to_valid_ready~0 (
	.dataa(!\doing_read~q ),
	.datab(!\general_counter[0]~q ),
	.datac(!\general_counter[1]~q ),
	.datad(!\doing_auto_precharge~q ),
	.datae(!\general_counter[3]~q ),
	.dataf(!\doing_precharge~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_rdwr_to_valid_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_rdwr_to_valid_ready~0 .extended_lut = "off";
defparam \int_rdwr_to_valid_ready~0 .lut_mask = 64'hA8EA000000000000;
defparam \int_rdwr_to_valid_ready~0 .shared_arith = "off";

arriaii_lcell_comb \int_rdwr_to_valid_ready~1 (
	.dataa(!\general_counter[0]~q ),
	.datab(!\general_counter[1]~q ),
	.datac(!\doing_precharge~q ),
	.datad(!\general_counter[5]~q ),
	.datae(!\general_counter[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_rdwr_to_valid_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_rdwr_to_valid_ready~1 .extended_lut = "off";
defparam \int_rdwr_to_valid_ready~1 .lut_mask = 64'hFE000000FE000000;
defparam \int_rdwr_to_valid_ready~1 .shared_arith = "off";

arriaii_lcell_comb \doing_read~0 (
	.dataa(!do_read_r),
	.datab(!to_chip_r_0),
	.datac(!do_write_r),
	.datad(!Equal0),
	.datae(!\doing_read~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_read~0 .extended_lut = "off";
defparam \doing_read~0 .lut_mask = 64'h0010FFFC0010FFFC;
defparam \doing_read~0 .shared_arith = "off";

dffeas doing_read(
	.clk(ctl_clk),
	.d(\doing_read~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_read~q ),
	.prn(vcc));
defparam doing_read.is_wysiwyg = "true";
defparam doing_read.power_up = "low";

arriaii_lcell_comb \int_rdwr_to_valid_ready~2 (
	.dataa(!act_to_rdwr_1),
	.datab(!\doing_read~q ),
	.datac(!\general_counter[1]~q ),
	.datad(!\doing_auto_precharge~q ),
	.datae(!\general_counter[3]~q ),
	.dataf(!\doing_precharge~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_rdwr_to_valid_ready~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_rdwr_to_valid_ready~2 .extended_lut = "off";
defparam \int_rdwr_to_valid_ready~2 .lut_mask = 64'h54550040FFFF0000;
defparam \int_rdwr_to_valid_ready~2 .shared_arith = "off";

arriaii_lcell_comb \int_rdwr_to_valid_ready~3 (
	.dataa(!close_0_0),
	.datab(!\general_counter[2]~q ),
	.datac(!\int_rdwr_to_valid_ready~0_combout ),
	.datad(!\int_rdwr_to_valid_ready~1_combout ),
	.datae(!\int_rdwr_to_valid_ready~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_rdwr_to_valid_ready~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_rdwr_to_valid_ready~3 .extended_lut = "off";
defparam \int_rdwr_to_valid_ready~3 .lut_mask = 64'h5555551055555510;
defparam \int_rdwr_to_valid_ready~3 .shared_arith = "off";

dffeas int_rdwr_to_valid_ready(
	.clk(ctl_clk),
	.d(\int_rdwr_to_valid_ready~3_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\int_rdwr_to_valid_ready~q ),
	.prn(vcc));
defparam int_rdwr_to_valid_ready.is_wysiwyg = "true";
defparam int_rdwr_to_valid_ready.power_up = "low";

arriaii_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~13 .shared_arith = "off";

arriaii_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \act_counter[4] (
	.clk(ctl_clk),
	.d(\Add0~17_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_0_0),
	.ena(vcc),
	.q(\act_counter[4]~q ),
	.prn(vcc));
defparam \act_counter[4] .is_wysiwyg = "true";
defparam \act_counter[4] .power_up = "low";

arriaii_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \act_counter[5] (
	.clk(ctl_clk),
	.d(\Add0~21_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_0_0),
	.ena(vcc),
	.q(\act_counter[5]~q ),
	.prn(vcc));
defparam \act_counter[5] .is_wysiwyg = "true";
defparam \act_counter[5] .power_up = "low";

arriaii_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Equal0~0_combout ),
	.datae(gnd),
	.dataf(!\act_counter[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF000000FF00;
defparam \Add0~1 .shared_arith = "off";

dffeas \act_counter[0] (
	.clk(ctl_clk),
	.d(\Add0~1_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_0_0),
	.ena(vcc),
	.q(\act_counter[0]~q ),
	.prn(vcc));
defparam \act_counter[0] .is_wysiwyg = "true";
defparam \act_counter[0] .power_up = "low";

arriaii_lcell_comb \Equal0~0 (
	.dataa(!\act_counter[3]~q ),
	.datab(!\act_counter[4]~q ),
	.datac(!\act_counter[5]~q ),
	.datad(!\act_counter[2]~q ),
	.datae(!\act_counter[1]~q ),
	.dataf(!\act_counter[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h0000000000000001;
defparam \Equal0~0 .shared_arith = "off";

arriaii_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \act_counter[1] (
	.clk(ctl_clk),
	.d(\Add0~5_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_0_0),
	.ena(vcc),
	.q(\act_counter[1]~q ),
	.prn(vcc));
defparam \act_counter[1] .is_wysiwyg = "true";
defparam \act_counter[1] .power_up = "low";

arriaii_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \act_counter[2] (
	.clk(ctl_clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_0_0),
	.ena(vcc),
	.q(\act_counter[2]~q ),
	.prn(vcc));
defparam \act_counter[2] .is_wysiwyg = "true";
defparam \act_counter[2] .power_up = "low";

dffeas \act_counter[3] (
	.clk(ctl_clk),
	.d(\Add0~13_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_0_0),
	.ena(vcc),
	.q(\act_counter[3]~q ),
	.prn(vcc));
defparam \act_counter[3] .is_wysiwyg = "true";
defparam \act_counter[3] .power_up = "low";

arriaii_lcell_comb \LessThan0~0 (
	.dataa(!act_to_rdwr_1),
	.datab(!\act_counter[3]~q ),
	.datac(!\act_counter[4]~q ),
	.datad(!\act_counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h4000400040004000;
defparam \LessThan0~0 .shared_arith = "off";

dffeas int_act_to_act_ready(
	.clk(ctl_clk),
	.d(\LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_0_0),
	.ena(vcc),
	.q(\int_act_to_act_ready~q ),
	.prn(vcc));
defparam int_act_to_act_ready.is_wysiwyg = "true";
defparam int_act_to_act_ready.power_up = "low";

arriaii_lcell_comb \rdwr_ready~0 (
	.dataa(!current_state1),
	.datab(!\LessThan0~0_combout ),
	.datac(!\act_counter[2]~q ),
	.datad(!\act_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdwr_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdwr_ready~0 .extended_lut = "off";
defparam \rdwr_ready~0 .lut_mask = 64'h4555455545554555;
defparam \rdwr_ready~0 .shared_arith = "off";

arriaii_lcell_comb \rdwr_ready~1 (
	.dataa(!act_to_rdwr_1),
	.datab(!close_0_0),
	.datac(!open_0_0),
	.datad(!\rdwr_ready~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdwr_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdwr_ready~1 .extended_lut = "off";
defparam \rdwr_ready~1 .lut_mask = 64'h0133013301330133;
defparam \rdwr_ready~1 .shared_arith = "off";

endmodule

module ddr3_int_alt_ddrx_bank_timer_info_1 (
	ctl_clk,
	do_read_r,
	do_write_r,
	current_state1,
	do_precharge_all_r,
	to_chip_r_0,
	always38,
	act_ready1,
	act_to_rdwr_1,
	always106,
	always145,
	ctl_reset_n,
	rdwr_ready1,
	always140,
	Equal0,
	close_1_0,
	open_1_0,
	general_counter,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	ctl_clk;
input 	do_read_r;
input 	do_write_r;
output 	current_state1;
input 	do_precharge_all_r;
input 	to_chip_r_0;
input 	always38;
output 	act_ready1;
input 	act_to_rdwr_1;
input 	always106;
input 	always145;
input 	ctl_reset_n;
output 	rdwr_ready1;
input 	always140;
input 	Equal0;
input 	close_1_0;
input 	open_1_0;
input 	general_counter;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \current_state~0_combout ;
wire \Add1~1_sumout ;
wire \general_counter~1_combout ;
wire \general_counter[0]~q ;
wire \Add1~10 ;
wire \Add1~13_sumout ;
wire \general_counter~3_combout ;
wire \general_counter[3]~q ;
wire \Add1~14 ;
wire \Add1~17_sumout ;
wire \general_counter~5_combout ;
wire \general_counter[4]~q ;
wire \Add1~18 ;
wire \Add1~21_sumout ;
wire \general_counter~4_combout ;
wire \general_counter[5]~q ;
wire \Equal1~0_combout ;
wire \Add1~2 ;
wire \Add1~5_sumout ;
wire \general_counter~2_combout ;
wire \general_counter[1]~q ;
wire \Add1~6 ;
wire \Add1~9_sumout ;
wire \general_counter~0_combout ;
wire \general_counter[2]~q ;
wire \doing_auto_precharge~0_combout ;
wire \doing_precharge~0_combout ;
wire \doing_auto_precharge~q ;
wire \doing_precharge~1_combout ;
wire \doing_precharge~q ;
wire \int_rdwr_to_valid_ready~0_combout ;
wire \int_rdwr_to_valid_ready~1_combout ;
wire \doing_read~0_combout ;
wire \doing_read~q ;
wire \int_rdwr_to_valid_ready~2_combout ;
wire \int_rdwr_to_valid_ready~3_combout ;
wire \int_rdwr_to_valid_ready~q ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \act_counter[4]~q ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \act_counter[5]~q ;
wire \Add0~1_sumout ;
wire \act_counter[0]~q ;
wire \Equal0~0_combout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \act_counter[1]~q ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \act_counter[2]~q ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \act_counter[3]~q ;
wire \LessThan0~0_combout ;
wire \int_act_to_act_ready~q ;
wire \rdwr_ready~0_combout ;
wire \rdwr_ready~1_combout ;


dffeas current_state(
	.clk(ctl_clk),
	.d(\current_state~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_1_0),
	.ena(vcc),
	.q(current_state1),
	.prn(vcc));
defparam current_state.is_wysiwyg = "true";
defparam current_state.power_up = "low";

arriaii_lcell_comb act_ready(
	.dataa(!\int_rdwr_to_valid_ready~q ),
	.datab(!\int_act_to_act_ready~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(act_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam act_ready.extended_lut = "off";
defparam act_ready.lut_mask = 64'h4444444444444444;
defparam act_ready.shared_arith = "off";

dffeas rdwr_ready(
	.clk(ctl_clk),
	.d(\rdwr_ready~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rdwr_ready1),
	.prn(vcc));
defparam rdwr_ready.is_wysiwyg = "true";
defparam rdwr_ready.power_up = "low";

arriaii_lcell_comb \current_state~0 (
	.dataa(!always38),
	.datab(!always106),
	.datac(!current_state1),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\current_state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \current_state~0 .extended_lut = "off";
defparam \current_state~0 .lut_mask = 64'h0C080C080C080C08;
defparam \current_state~0 .shared_arith = "off";

arriaii_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Equal1~0_combout ),
	.datae(gnd),
	.dataf(!\general_counter[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(\Add1~2 ),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h0000FF000000FF00;
defparam \Add1~1 .shared_arith = "off";

arriaii_lcell_comb \general_counter~1 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~1_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~1 .extended_lut = "off";
defparam \general_counter~1 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~1 .shared_arith = "off";

dffeas \general_counter[0] (
	.clk(ctl_clk),
	.d(\general_counter~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[0]~q ),
	.prn(vcc));
defparam \general_counter[0] .is_wysiwyg = "true";
defparam \general_counter[0] .power_up = "low";

arriaii_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~9 .shared_arith = "off";

arriaii_lcell_comb \Add1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~13 .shared_arith = "off";

arriaii_lcell_comb \general_counter~3 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~13_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~3 .extended_lut = "off";
defparam \general_counter~3 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~3 .shared_arith = "off";

dffeas \general_counter[3] (
	.clk(ctl_clk),
	.d(\general_counter~3_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[3]~q ),
	.prn(vcc));
defparam \general_counter[3] .is_wysiwyg = "true";
defparam \general_counter[3] .power_up = "low";

arriaii_lcell_comb \Add1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~17 .shared_arith = "off";

arriaii_lcell_comb \general_counter~5 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~17_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~5 .extended_lut = "off";
defparam \general_counter~5 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~5 .shared_arith = "off";

dffeas \general_counter[4] (
	.clk(ctl_clk),
	.d(\general_counter~5_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[4]~q ),
	.prn(vcc));
defparam \general_counter[4] .is_wysiwyg = "true";
defparam \general_counter[4] .power_up = "low";

arriaii_lcell_comb \Add1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~21_sumout ),
	.cout(),
	.shareout());
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~21 .shared_arith = "off";

arriaii_lcell_comb \general_counter~4 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~21_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~4 .extended_lut = "off";
defparam \general_counter~4 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~4 .shared_arith = "off";

dffeas \general_counter[5] (
	.clk(ctl_clk),
	.d(\general_counter~4_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[5]~q ),
	.prn(vcc));
defparam \general_counter[5] .is_wysiwyg = "true";
defparam \general_counter[5] .power_up = "low";

arriaii_lcell_comb \Equal1~0 (
	.dataa(!\general_counter[2]~q ),
	.datab(!\general_counter[0]~q ),
	.datac(!\general_counter[1]~q ),
	.datad(!\general_counter[3]~q ),
	.datae(!\general_counter[5]~q ),
	.dataf(!\general_counter[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'h0000000000000001;
defparam \Equal1~0 .shared_arith = "off";

arriaii_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~5 .shared_arith = "off";

arriaii_lcell_comb \general_counter~2 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~5_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~2 .extended_lut = "off";
defparam \general_counter~2 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~2 .shared_arith = "off";

dffeas \general_counter[1] (
	.clk(ctl_clk),
	.d(\general_counter~2_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[1]~q ),
	.prn(vcc));
defparam \general_counter[1] .is_wysiwyg = "true";
defparam \general_counter[1] .power_up = "low";

arriaii_lcell_comb \general_counter~0 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~9_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~0 .extended_lut = "off";
defparam \general_counter~0 .lut_mask = 64'h1311FFFF1311FFFF;
defparam \general_counter~0 .shared_arith = "off";

dffeas \general_counter[2] (
	.clk(ctl_clk),
	.d(\general_counter~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[2]~q ),
	.prn(vcc));
defparam \general_counter[2] .is_wysiwyg = "true";
defparam \general_counter[2] .power_up = "low";

arriaii_lcell_comb \doing_auto_precharge~0 (
	.dataa(!always38),
	.datab(!always106),
	.datac(!always140),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_auto_precharge~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_auto_precharge~0 .extended_lut = "off";
defparam \doing_auto_precharge~0 .lut_mask = 64'h0007000700070007;
defparam \doing_auto_precharge~0 .shared_arith = "off";

arriaii_lcell_comb \doing_precharge~0 (
	.dataa(!always38),
	.datab(!always145),
	.datac(!always106),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_precharge~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_precharge~0 .extended_lut = "off";
defparam \doing_precharge~0 .lut_mask = 64'h0F7F0F7F0F7F0F7F;
defparam \doing_precharge~0 .shared_arith = "off";

dffeas doing_auto_precharge(
	.clk(ctl_clk),
	.d(\doing_auto_precharge~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\doing_precharge~0_combout ),
	.q(\doing_auto_precharge~q ),
	.prn(vcc));
defparam doing_auto_precharge.is_wysiwyg = "true";
defparam doing_auto_precharge.power_up = "low";

arriaii_lcell_comb \doing_precharge~1 (
	.dataa(!always38),
	.datab(!always106),
	.datac(!always140),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_precharge~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_precharge~1 .extended_lut = "off";
defparam \doing_precharge~1 .lut_mask = 64'h3370337033703370;
defparam \doing_precharge~1 .shared_arith = "off";

dffeas doing_precharge(
	.clk(ctl_clk),
	.d(\doing_precharge~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\doing_precharge~0_combout ),
	.q(\doing_precharge~q ),
	.prn(vcc));
defparam doing_precharge.is_wysiwyg = "true";
defparam doing_precharge.power_up = "low";

arriaii_lcell_comb \int_rdwr_to_valid_ready~0 (
	.dataa(!\doing_read~q ),
	.datab(!\general_counter[0]~q ),
	.datac(!\general_counter[1]~q ),
	.datad(!\doing_auto_precharge~q ),
	.datae(!\general_counter[3]~q ),
	.dataf(!\doing_precharge~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_rdwr_to_valid_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_rdwr_to_valid_ready~0 .extended_lut = "off";
defparam \int_rdwr_to_valid_ready~0 .lut_mask = 64'hA8EA000000000000;
defparam \int_rdwr_to_valid_ready~0 .shared_arith = "off";

arriaii_lcell_comb \int_rdwr_to_valid_ready~1 (
	.dataa(!\general_counter[0]~q ),
	.datab(!\general_counter[1]~q ),
	.datac(!\doing_precharge~q ),
	.datad(!\general_counter[5]~q ),
	.datae(!\general_counter[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_rdwr_to_valid_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_rdwr_to_valid_ready~1 .extended_lut = "off";
defparam \int_rdwr_to_valid_ready~1 .lut_mask = 64'hFE000000FE000000;
defparam \int_rdwr_to_valid_ready~1 .shared_arith = "off";

arriaii_lcell_comb \doing_read~0 (
	.dataa(!do_read_r),
	.datab(!to_chip_r_0),
	.datac(!do_write_r),
	.datad(!Equal0),
	.datae(!\doing_read~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_read~0 .extended_lut = "off";
defparam \doing_read~0 .lut_mask = 64'h0010FFFC0010FFFC;
defparam \doing_read~0 .shared_arith = "off";

dffeas doing_read(
	.clk(ctl_clk),
	.d(\doing_read~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_read~q ),
	.prn(vcc));
defparam doing_read.is_wysiwyg = "true";
defparam doing_read.power_up = "low";

arriaii_lcell_comb \int_rdwr_to_valid_ready~2 (
	.dataa(!act_to_rdwr_1),
	.datab(!\doing_read~q ),
	.datac(!\general_counter[1]~q ),
	.datad(!\doing_auto_precharge~q ),
	.datae(!\general_counter[3]~q ),
	.dataf(!\doing_precharge~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_rdwr_to_valid_ready~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_rdwr_to_valid_ready~2 .extended_lut = "off";
defparam \int_rdwr_to_valid_ready~2 .lut_mask = 64'h54550040FFFF0000;
defparam \int_rdwr_to_valid_ready~2 .shared_arith = "off";

arriaii_lcell_comb \int_rdwr_to_valid_ready~3 (
	.dataa(!close_1_0),
	.datab(!\general_counter[2]~q ),
	.datac(!\int_rdwr_to_valid_ready~0_combout ),
	.datad(!\int_rdwr_to_valid_ready~1_combout ),
	.datae(!\int_rdwr_to_valid_ready~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_rdwr_to_valid_ready~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_rdwr_to_valid_ready~3 .extended_lut = "off";
defparam \int_rdwr_to_valid_ready~3 .lut_mask = 64'h5555551055555510;
defparam \int_rdwr_to_valid_ready~3 .shared_arith = "off";

dffeas int_rdwr_to_valid_ready(
	.clk(ctl_clk),
	.d(\int_rdwr_to_valid_ready~3_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\int_rdwr_to_valid_ready~q ),
	.prn(vcc));
defparam int_rdwr_to_valid_ready.is_wysiwyg = "true";
defparam int_rdwr_to_valid_ready.power_up = "low";

arriaii_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~13 .shared_arith = "off";

arriaii_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \act_counter[4] (
	.clk(ctl_clk),
	.d(\Add0~17_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_1_0),
	.ena(vcc),
	.q(\act_counter[4]~q ),
	.prn(vcc));
defparam \act_counter[4] .is_wysiwyg = "true";
defparam \act_counter[4] .power_up = "low";

arriaii_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \act_counter[5] (
	.clk(ctl_clk),
	.d(\Add0~21_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_1_0),
	.ena(vcc),
	.q(\act_counter[5]~q ),
	.prn(vcc));
defparam \act_counter[5] .is_wysiwyg = "true";
defparam \act_counter[5] .power_up = "low";

arriaii_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Equal0~0_combout ),
	.datae(gnd),
	.dataf(!\act_counter[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF000000FF00;
defparam \Add0~1 .shared_arith = "off";

dffeas \act_counter[0] (
	.clk(ctl_clk),
	.d(\Add0~1_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_1_0),
	.ena(vcc),
	.q(\act_counter[0]~q ),
	.prn(vcc));
defparam \act_counter[0] .is_wysiwyg = "true";
defparam \act_counter[0] .power_up = "low";

arriaii_lcell_comb \Equal0~0 (
	.dataa(!\act_counter[3]~q ),
	.datab(!\act_counter[4]~q ),
	.datac(!\act_counter[5]~q ),
	.datad(!\act_counter[2]~q ),
	.datae(!\act_counter[1]~q ),
	.dataf(!\act_counter[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h0000000000000001;
defparam \Equal0~0 .shared_arith = "off";

arriaii_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \act_counter[1] (
	.clk(ctl_clk),
	.d(\Add0~5_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_1_0),
	.ena(vcc),
	.q(\act_counter[1]~q ),
	.prn(vcc));
defparam \act_counter[1] .is_wysiwyg = "true";
defparam \act_counter[1] .power_up = "low";

arriaii_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \act_counter[2] (
	.clk(ctl_clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_1_0),
	.ena(vcc),
	.q(\act_counter[2]~q ),
	.prn(vcc));
defparam \act_counter[2] .is_wysiwyg = "true";
defparam \act_counter[2] .power_up = "low";

dffeas \act_counter[3] (
	.clk(ctl_clk),
	.d(\Add0~13_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_1_0),
	.ena(vcc),
	.q(\act_counter[3]~q ),
	.prn(vcc));
defparam \act_counter[3] .is_wysiwyg = "true";
defparam \act_counter[3] .power_up = "low";

arriaii_lcell_comb \LessThan0~0 (
	.dataa(!act_to_rdwr_1),
	.datab(!\act_counter[3]~q ),
	.datac(!\act_counter[4]~q ),
	.datad(!\act_counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h4000400040004000;
defparam \LessThan0~0 .shared_arith = "off";

dffeas int_act_to_act_ready(
	.clk(ctl_clk),
	.d(\LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_1_0),
	.ena(vcc),
	.q(\int_act_to_act_ready~q ),
	.prn(vcc));
defparam int_act_to_act_ready.is_wysiwyg = "true";
defparam int_act_to_act_ready.power_up = "low";

arriaii_lcell_comb \rdwr_ready~0 (
	.dataa(!current_state1),
	.datab(!\LessThan0~0_combout ),
	.datac(!\act_counter[2]~q ),
	.datad(!\act_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdwr_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdwr_ready~0 .extended_lut = "off";
defparam \rdwr_ready~0 .lut_mask = 64'h4555455545554555;
defparam \rdwr_ready~0 .shared_arith = "off";

arriaii_lcell_comb \rdwr_ready~1 (
	.dataa(!act_to_rdwr_1),
	.datab(!close_1_0),
	.datac(!open_1_0),
	.datad(!\rdwr_ready~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdwr_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdwr_ready~1 .extended_lut = "off";
defparam \rdwr_ready~1 .lut_mask = 64'h0133013301330133;
defparam \rdwr_ready~1 .shared_arith = "off";

endmodule

module ddr3_int_alt_ddrx_bank_timer_info_2 (
	ctl_clk,
	do_read_r,
	do_write_r,
	current_state1,
	do_precharge_all_r,
	to_chip_r_0,
	always38,
	act_ready1,
	act_to_rdwr_1,
	always106,
	always145,
	ctl_reset_n,
	rdwr_ready1,
	always140,
	Equal0,
	close_2_0,
	open_2_0,
	general_counter,
	always1,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	ctl_clk;
input 	do_read_r;
input 	do_write_r;
output 	current_state1;
input 	do_precharge_all_r;
input 	to_chip_r_0;
input 	always38;
output 	act_ready1;
input 	act_to_rdwr_1;
input 	always106;
input 	always145;
input 	ctl_reset_n;
output 	rdwr_ready1;
input 	always140;
input 	Equal0;
input 	close_2_0;
input 	open_2_0;
input 	general_counter;
output 	always1;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \current_state~0_combout ;
wire \Add1~1_sumout ;
wire \general_counter~1_combout ;
wire \general_counter[0]~q ;
wire \Add1~10 ;
wire \Add1~13_sumout ;
wire \general_counter~3_combout ;
wire \general_counter[3]~q ;
wire \Add1~14 ;
wire \Add1~17_sumout ;
wire \general_counter~5_combout ;
wire \general_counter[4]~q ;
wire \Add1~18 ;
wire \Add1~21_sumout ;
wire \general_counter~4_combout ;
wire \general_counter[5]~q ;
wire \Equal1~0_combout ;
wire \Add1~2 ;
wire \Add1~5_sumout ;
wire \general_counter~2_combout ;
wire \general_counter[1]~q ;
wire \Add1~6 ;
wire \Add1~9_sumout ;
wire \general_counter~0_combout ;
wire \general_counter[2]~q ;
wire \doing_auto_precharge~0_combout ;
wire \doing_precharge~0_combout ;
wire \doing_auto_precharge~q ;
wire \doing_precharge~1_combout ;
wire \doing_precharge~q ;
wire \int_rdwr_to_valid_ready~0_combout ;
wire \int_rdwr_to_valid_ready~1_combout ;
wire \doing_read~0_combout ;
wire \doing_read~q ;
wire \int_rdwr_to_valid_ready~2_combout ;
wire \int_rdwr_to_valid_ready~3_combout ;
wire \int_rdwr_to_valid_ready~q ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \act_counter[4]~q ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \act_counter[5]~q ;
wire \Add0~1_sumout ;
wire \act_counter[0]~q ;
wire \Equal0~0_combout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \act_counter[1]~q ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \act_counter[2]~q ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \act_counter[3]~q ;
wire \LessThan0~0_combout ;
wire \int_act_to_act_ready~q ;
wire \rdwr_ready~0_combout ;
wire \rdwr_ready~1_combout ;


dffeas current_state(
	.clk(ctl_clk),
	.d(\current_state~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_2_0),
	.ena(vcc),
	.q(current_state1),
	.prn(vcc));
defparam current_state.is_wysiwyg = "true";
defparam current_state.power_up = "low";

arriaii_lcell_comb act_ready(
	.dataa(!\int_rdwr_to_valid_ready~q ),
	.datab(!\int_act_to_act_ready~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(act_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam act_ready.extended_lut = "off";
defparam act_ready.lut_mask = 64'h4444444444444444;
defparam act_ready.shared_arith = "off";

dffeas rdwr_ready(
	.clk(ctl_clk),
	.d(\rdwr_ready~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rdwr_ready1),
	.prn(vcc));
defparam rdwr_ready.is_wysiwyg = "true";
defparam rdwr_ready.power_up = "low";

arriaii_lcell_comb \always1~0 (
	.dataa(!do_read_r),
	.datab(!do_write_r),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always1),
	.sumout(),
	.cout(),
	.shareout());
defparam \always1~0 .extended_lut = "off";
defparam \always1~0 .lut_mask = 64'h7777777777777777;
defparam \always1~0 .shared_arith = "off";

arriaii_lcell_comb \current_state~0 (
	.dataa(!always38),
	.datab(!always106),
	.datac(!current_state1),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\current_state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \current_state~0 .extended_lut = "off";
defparam \current_state~0 .lut_mask = 64'h0C080C080C080C08;
defparam \current_state~0 .shared_arith = "off";

arriaii_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Equal1~0_combout ),
	.datae(gnd),
	.dataf(!\general_counter[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(\Add1~2 ),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h0000FF000000FF00;
defparam \Add1~1 .shared_arith = "off";

arriaii_lcell_comb \general_counter~1 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~1_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~1 .extended_lut = "off";
defparam \general_counter~1 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~1 .shared_arith = "off";

dffeas \general_counter[0] (
	.clk(ctl_clk),
	.d(\general_counter~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[0]~q ),
	.prn(vcc));
defparam \general_counter[0] .is_wysiwyg = "true";
defparam \general_counter[0] .power_up = "low";

arriaii_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~9 .shared_arith = "off";

arriaii_lcell_comb \Add1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~13 .shared_arith = "off";

arriaii_lcell_comb \general_counter~3 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~13_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~3 .extended_lut = "off";
defparam \general_counter~3 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~3 .shared_arith = "off";

dffeas \general_counter[3] (
	.clk(ctl_clk),
	.d(\general_counter~3_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[3]~q ),
	.prn(vcc));
defparam \general_counter[3] .is_wysiwyg = "true";
defparam \general_counter[3] .power_up = "low";

arriaii_lcell_comb \Add1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~17 .shared_arith = "off";

arriaii_lcell_comb \general_counter~5 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~17_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~5 .extended_lut = "off";
defparam \general_counter~5 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~5 .shared_arith = "off";

dffeas \general_counter[4] (
	.clk(ctl_clk),
	.d(\general_counter~5_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[4]~q ),
	.prn(vcc));
defparam \general_counter[4] .is_wysiwyg = "true";
defparam \general_counter[4] .power_up = "low";

arriaii_lcell_comb \Add1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~21_sumout ),
	.cout(),
	.shareout());
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~21 .shared_arith = "off";

arriaii_lcell_comb \general_counter~4 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~21_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~4 .extended_lut = "off";
defparam \general_counter~4 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~4 .shared_arith = "off";

dffeas \general_counter[5] (
	.clk(ctl_clk),
	.d(\general_counter~4_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[5]~q ),
	.prn(vcc));
defparam \general_counter[5] .is_wysiwyg = "true";
defparam \general_counter[5] .power_up = "low";

arriaii_lcell_comb \Equal1~0 (
	.dataa(!\general_counter[2]~q ),
	.datab(!\general_counter[0]~q ),
	.datac(!\general_counter[1]~q ),
	.datad(!\general_counter[3]~q ),
	.datae(!\general_counter[5]~q ),
	.dataf(!\general_counter[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'h0000000000000001;
defparam \Equal1~0 .shared_arith = "off";

arriaii_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~5 .shared_arith = "off";

arriaii_lcell_comb \general_counter~2 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~5_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~2 .extended_lut = "off";
defparam \general_counter~2 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~2 .shared_arith = "off";

dffeas \general_counter[1] (
	.clk(ctl_clk),
	.d(\general_counter~2_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[1]~q ),
	.prn(vcc));
defparam \general_counter[1] .is_wysiwyg = "true";
defparam \general_counter[1] .power_up = "low";

arriaii_lcell_comb \general_counter~0 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~9_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~0 .extended_lut = "off";
defparam \general_counter~0 .lut_mask = 64'h1311FFFF1311FFFF;
defparam \general_counter~0 .shared_arith = "off";

dffeas \general_counter[2] (
	.clk(ctl_clk),
	.d(\general_counter~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[2]~q ),
	.prn(vcc));
defparam \general_counter[2] .is_wysiwyg = "true";
defparam \general_counter[2] .power_up = "low";

arriaii_lcell_comb \doing_auto_precharge~0 (
	.dataa(!always38),
	.datab(!always106),
	.datac(!always140),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_auto_precharge~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_auto_precharge~0 .extended_lut = "off";
defparam \doing_auto_precharge~0 .lut_mask = 64'h0007000700070007;
defparam \doing_auto_precharge~0 .shared_arith = "off";

arriaii_lcell_comb \doing_precharge~0 (
	.dataa(!always38),
	.datab(!always145),
	.datac(!always106),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_precharge~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_precharge~0 .extended_lut = "off";
defparam \doing_precharge~0 .lut_mask = 64'h0F7F0F7F0F7F0F7F;
defparam \doing_precharge~0 .shared_arith = "off";

dffeas doing_auto_precharge(
	.clk(ctl_clk),
	.d(\doing_auto_precharge~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\doing_precharge~0_combout ),
	.q(\doing_auto_precharge~q ),
	.prn(vcc));
defparam doing_auto_precharge.is_wysiwyg = "true";
defparam doing_auto_precharge.power_up = "low";

arriaii_lcell_comb \doing_precharge~1 (
	.dataa(!always38),
	.datab(!always106),
	.datac(!always140),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_precharge~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_precharge~1 .extended_lut = "off";
defparam \doing_precharge~1 .lut_mask = 64'h3370337033703370;
defparam \doing_precharge~1 .shared_arith = "off";

dffeas doing_precharge(
	.clk(ctl_clk),
	.d(\doing_precharge~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\doing_precharge~0_combout ),
	.q(\doing_precharge~q ),
	.prn(vcc));
defparam doing_precharge.is_wysiwyg = "true";
defparam doing_precharge.power_up = "low";

arriaii_lcell_comb \int_rdwr_to_valid_ready~0 (
	.dataa(!\doing_read~q ),
	.datab(!\general_counter[0]~q ),
	.datac(!\general_counter[1]~q ),
	.datad(!\doing_auto_precharge~q ),
	.datae(!\general_counter[3]~q ),
	.dataf(!\doing_precharge~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_rdwr_to_valid_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_rdwr_to_valid_ready~0 .extended_lut = "off";
defparam \int_rdwr_to_valid_ready~0 .lut_mask = 64'hA8EA000000000000;
defparam \int_rdwr_to_valid_ready~0 .shared_arith = "off";

arriaii_lcell_comb \int_rdwr_to_valid_ready~1 (
	.dataa(!\general_counter[0]~q ),
	.datab(!\general_counter[1]~q ),
	.datac(!\doing_precharge~q ),
	.datad(!\general_counter[5]~q ),
	.datae(!\general_counter[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_rdwr_to_valid_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_rdwr_to_valid_ready~1 .extended_lut = "off";
defparam \int_rdwr_to_valid_ready~1 .lut_mask = 64'hFE000000FE000000;
defparam \int_rdwr_to_valid_ready~1 .shared_arith = "off";

arriaii_lcell_comb \doing_read~0 (
	.dataa(!do_read_r),
	.datab(!to_chip_r_0),
	.datac(!do_write_r),
	.datad(!Equal0),
	.datae(!\doing_read~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_read~0 .extended_lut = "off";
defparam \doing_read~0 .lut_mask = 64'h0010FFFC0010FFFC;
defparam \doing_read~0 .shared_arith = "off";

dffeas doing_read(
	.clk(ctl_clk),
	.d(\doing_read~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_read~q ),
	.prn(vcc));
defparam doing_read.is_wysiwyg = "true";
defparam doing_read.power_up = "low";

arriaii_lcell_comb \int_rdwr_to_valid_ready~2 (
	.dataa(!act_to_rdwr_1),
	.datab(!\doing_read~q ),
	.datac(!\general_counter[1]~q ),
	.datad(!\doing_auto_precharge~q ),
	.datae(!\general_counter[3]~q ),
	.dataf(!\doing_precharge~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_rdwr_to_valid_ready~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_rdwr_to_valid_ready~2 .extended_lut = "off";
defparam \int_rdwr_to_valid_ready~2 .lut_mask = 64'h54550040FFFF0000;
defparam \int_rdwr_to_valid_ready~2 .shared_arith = "off";

arriaii_lcell_comb \int_rdwr_to_valid_ready~3 (
	.dataa(!close_2_0),
	.datab(!\general_counter[2]~q ),
	.datac(!\int_rdwr_to_valid_ready~0_combout ),
	.datad(!\int_rdwr_to_valid_ready~1_combout ),
	.datae(!\int_rdwr_to_valid_ready~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_rdwr_to_valid_ready~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_rdwr_to_valid_ready~3 .extended_lut = "off";
defparam \int_rdwr_to_valid_ready~3 .lut_mask = 64'h5555551055555510;
defparam \int_rdwr_to_valid_ready~3 .shared_arith = "off";

dffeas int_rdwr_to_valid_ready(
	.clk(ctl_clk),
	.d(\int_rdwr_to_valid_ready~3_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\int_rdwr_to_valid_ready~q ),
	.prn(vcc));
defparam int_rdwr_to_valid_ready.is_wysiwyg = "true";
defparam int_rdwr_to_valid_ready.power_up = "low";

arriaii_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~13 .shared_arith = "off";

arriaii_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \act_counter[4] (
	.clk(ctl_clk),
	.d(\Add0~17_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_2_0),
	.ena(vcc),
	.q(\act_counter[4]~q ),
	.prn(vcc));
defparam \act_counter[4] .is_wysiwyg = "true";
defparam \act_counter[4] .power_up = "low";

arriaii_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \act_counter[5] (
	.clk(ctl_clk),
	.d(\Add0~21_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_2_0),
	.ena(vcc),
	.q(\act_counter[5]~q ),
	.prn(vcc));
defparam \act_counter[5] .is_wysiwyg = "true";
defparam \act_counter[5] .power_up = "low";

arriaii_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Equal0~0_combout ),
	.datae(gnd),
	.dataf(!\act_counter[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF000000FF00;
defparam \Add0~1 .shared_arith = "off";

dffeas \act_counter[0] (
	.clk(ctl_clk),
	.d(\Add0~1_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_2_0),
	.ena(vcc),
	.q(\act_counter[0]~q ),
	.prn(vcc));
defparam \act_counter[0] .is_wysiwyg = "true";
defparam \act_counter[0] .power_up = "low";

arriaii_lcell_comb \Equal0~0 (
	.dataa(!\act_counter[3]~q ),
	.datab(!\act_counter[4]~q ),
	.datac(!\act_counter[5]~q ),
	.datad(!\act_counter[2]~q ),
	.datae(!\act_counter[1]~q ),
	.dataf(!\act_counter[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h0000000000000001;
defparam \Equal0~0 .shared_arith = "off";

arriaii_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \act_counter[1] (
	.clk(ctl_clk),
	.d(\Add0~5_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_2_0),
	.ena(vcc),
	.q(\act_counter[1]~q ),
	.prn(vcc));
defparam \act_counter[1] .is_wysiwyg = "true";
defparam \act_counter[1] .power_up = "low";

arriaii_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \act_counter[2] (
	.clk(ctl_clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_2_0),
	.ena(vcc),
	.q(\act_counter[2]~q ),
	.prn(vcc));
defparam \act_counter[2] .is_wysiwyg = "true";
defparam \act_counter[2] .power_up = "low";

dffeas \act_counter[3] (
	.clk(ctl_clk),
	.d(\Add0~13_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_2_0),
	.ena(vcc),
	.q(\act_counter[3]~q ),
	.prn(vcc));
defparam \act_counter[3] .is_wysiwyg = "true";
defparam \act_counter[3] .power_up = "low";

arriaii_lcell_comb \LessThan0~0 (
	.dataa(!act_to_rdwr_1),
	.datab(!\act_counter[3]~q ),
	.datac(!\act_counter[4]~q ),
	.datad(!\act_counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h4000400040004000;
defparam \LessThan0~0 .shared_arith = "off";

dffeas int_act_to_act_ready(
	.clk(ctl_clk),
	.d(\LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_2_0),
	.ena(vcc),
	.q(\int_act_to_act_ready~q ),
	.prn(vcc));
defparam int_act_to_act_ready.is_wysiwyg = "true";
defparam int_act_to_act_ready.power_up = "low";

arriaii_lcell_comb \rdwr_ready~0 (
	.dataa(!current_state1),
	.datab(!\LessThan0~0_combout ),
	.datac(!\act_counter[2]~q ),
	.datad(!\act_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdwr_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdwr_ready~0 .extended_lut = "off";
defparam \rdwr_ready~0 .lut_mask = 64'h4555455545554555;
defparam \rdwr_ready~0 .shared_arith = "off";

arriaii_lcell_comb \rdwr_ready~1 (
	.dataa(!act_to_rdwr_1),
	.datab(!close_2_0),
	.datac(!open_2_0),
	.datad(!\rdwr_ready~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdwr_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdwr_ready~1 .extended_lut = "off";
defparam \rdwr_ready~1 .lut_mask = 64'h0133013301330133;
defparam \rdwr_ready~1 .shared_arith = "off";

endmodule

module ddr3_int_alt_ddrx_bank_timer_info_3 (
	ctl_clk,
	do_read_r,
	do_write_r,
	current_state1,
	do_precharge_all_r,
	to_chip_r_0,
	always38,
	act_ready1,
	act_to_rdwr_1,
	always106,
	always145,
	ctl_reset_n,
	rdwr_ready1,
	always140,
	Equal0,
	close_3_0,
	open_3_0,
	general_counter,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	ctl_clk;
input 	do_read_r;
input 	do_write_r;
output 	current_state1;
input 	do_precharge_all_r;
input 	to_chip_r_0;
input 	always38;
output 	act_ready1;
input 	act_to_rdwr_1;
input 	always106;
input 	always145;
input 	ctl_reset_n;
output 	rdwr_ready1;
input 	always140;
input 	Equal0;
input 	close_3_0;
input 	open_3_0;
input 	general_counter;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \current_state~0_combout ;
wire \Add1~1_sumout ;
wire \general_counter~1_combout ;
wire \general_counter[0]~q ;
wire \Add1~10 ;
wire \Add1~13_sumout ;
wire \general_counter~3_combout ;
wire \general_counter[3]~q ;
wire \Add1~14 ;
wire \Add1~17_sumout ;
wire \general_counter~5_combout ;
wire \general_counter[4]~q ;
wire \Add1~18 ;
wire \Add1~21_sumout ;
wire \general_counter~4_combout ;
wire \general_counter[5]~q ;
wire \Equal1~0_combout ;
wire \Add1~2 ;
wire \Add1~5_sumout ;
wire \general_counter~2_combout ;
wire \general_counter[1]~q ;
wire \Add1~6 ;
wire \Add1~9_sumout ;
wire \general_counter~0_combout ;
wire \general_counter[2]~q ;
wire \doing_auto_precharge~0_combout ;
wire \doing_precharge~0_combout ;
wire \doing_auto_precharge~q ;
wire \doing_precharge~1_combout ;
wire \doing_precharge~q ;
wire \int_rdwr_to_valid_ready~0_combout ;
wire \int_rdwr_to_valid_ready~1_combout ;
wire \doing_read~0_combout ;
wire \doing_read~q ;
wire \int_rdwr_to_valid_ready~2_combout ;
wire \int_rdwr_to_valid_ready~3_combout ;
wire \int_rdwr_to_valid_ready~q ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \act_counter[4]~q ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \act_counter[5]~q ;
wire \Add0~1_sumout ;
wire \act_counter[0]~q ;
wire \Equal0~0_combout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \act_counter[1]~q ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \act_counter[2]~q ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \act_counter[3]~q ;
wire \LessThan0~0_combout ;
wire \int_act_to_act_ready~q ;
wire \rdwr_ready~0_combout ;
wire \rdwr_ready~1_combout ;


dffeas current_state(
	.clk(ctl_clk),
	.d(\current_state~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_3_0),
	.ena(vcc),
	.q(current_state1),
	.prn(vcc));
defparam current_state.is_wysiwyg = "true";
defparam current_state.power_up = "low";

arriaii_lcell_comb act_ready(
	.dataa(!\int_rdwr_to_valid_ready~q ),
	.datab(!\int_act_to_act_ready~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(act_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam act_ready.extended_lut = "off";
defparam act_ready.lut_mask = 64'h4444444444444444;
defparam act_ready.shared_arith = "off";

dffeas rdwr_ready(
	.clk(ctl_clk),
	.d(\rdwr_ready~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rdwr_ready1),
	.prn(vcc));
defparam rdwr_ready.is_wysiwyg = "true";
defparam rdwr_ready.power_up = "low";

arriaii_lcell_comb \current_state~0 (
	.dataa(!always38),
	.datab(!always106),
	.datac(!current_state1),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\current_state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \current_state~0 .extended_lut = "off";
defparam \current_state~0 .lut_mask = 64'h0C080C080C080C08;
defparam \current_state~0 .shared_arith = "off";

arriaii_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Equal1~0_combout ),
	.datae(gnd),
	.dataf(!\general_counter[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(\Add1~2 ),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h0000FF000000FF00;
defparam \Add1~1 .shared_arith = "off";

arriaii_lcell_comb \general_counter~1 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~1_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~1 .extended_lut = "off";
defparam \general_counter~1 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~1 .shared_arith = "off";

dffeas \general_counter[0] (
	.clk(ctl_clk),
	.d(\general_counter~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[0]~q ),
	.prn(vcc));
defparam \general_counter[0] .is_wysiwyg = "true";
defparam \general_counter[0] .power_up = "low";

arriaii_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~9 .shared_arith = "off";

arriaii_lcell_comb \Add1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~13 .shared_arith = "off";

arriaii_lcell_comb \general_counter~3 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~13_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~3 .extended_lut = "off";
defparam \general_counter~3 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~3 .shared_arith = "off";

dffeas \general_counter[3] (
	.clk(ctl_clk),
	.d(\general_counter~3_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[3]~q ),
	.prn(vcc));
defparam \general_counter[3] .is_wysiwyg = "true";
defparam \general_counter[3] .power_up = "low";

arriaii_lcell_comb \Add1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~17 .shared_arith = "off";

arriaii_lcell_comb \general_counter~5 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~17_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~5 .extended_lut = "off";
defparam \general_counter~5 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~5 .shared_arith = "off";

dffeas \general_counter[4] (
	.clk(ctl_clk),
	.d(\general_counter~5_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[4]~q ),
	.prn(vcc));
defparam \general_counter[4] .is_wysiwyg = "true";
defparam \general_counter[4] .power_up = "low";

arriaii_lcell_comb \Add1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~21_sumout ),
	.cout(),
	.shareout());
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~21 .shared_arith = "off";

arriaii_lcell_comb \general_counter~4 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~21_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~4 .extended_lut = "off";
defparam \general_counter~4 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~4 .shared_arith = "off";

dffeas \general_counter[5] (
	.clk(ctl_clk),
	.d(\general_counter~4_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[5]~q ),
	.prn(vcc));
defparam \general_counter[5] .is_wysiwyg = "true";
defparam \general_counter[5] .power_up = "low";

arriaii_lcell_comb \Equal1~0 (
	.dataa(!\general_counter[2]~q ),
	.datab(!\general_counter[0]~q ),
	.datac(!\general_counter[1]~q ),
	.datad(!\general_counter[3]~q ),
	.datae(!\general_counter[5]~q ),
	.dataf(!\general_counter[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'h0000000000000001;
defparam \Equal1~0 .shared_arith = "off";

arriaii_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~5 .shared_arith = "off";

arriaii_lcell_comb \general_counter~2 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~5_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~2 .extended_lut = "off";
defparam \general_counter~2 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~2 .shared_arith = "off";

dffeas \general_counter[1] (
	.clk(ctl_clk),
	.d(\general_counter~2_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[1]~q ),
	.prn(vcc));
defparam \general_counter[1] .is_wysiwyg = "true";
defparam \general_counter[1] .power_up = "low";

arriaii_lcell_comb \general_counter~0 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~9_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~0 .extended_lut = "off";
defparam \general_counter~0 .lut_mask = 64'h1311FFFF1311FFFF;
defparam \general_counter~0 .shared_arith = "off";

dffeas \general_counter[2] (
	.clk(ctl_clk),
	.d(\general_counter~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[2]~q ),
	.prn(vcc));
defparam \general_counter[2] .is_wysiwyg = "true";
defparam \general_counter[2] .power_up = "low";

arriaii_lcell_comb \doing_auto_precharge~0 (
	.dataa(!always38),
	.datab(!always106),
	.datac(!always140),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_auto_precharge~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_auto_precharge~0 .extended_lut = "off";
defparam \doing_auto_precharge~0 .lut_mask = 64'h0007000700070007;
defparam \doing_auto_precharge~0 .shared_arith = "off";

arriaii_lcell_comb \doing_precharge~0 (
	.dataa(!always38),
	.datab(!always145),
	.datac(!always106),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_precharge~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_precharge~0 .extended_lut = "off";
defparam \doing_precharge~0 .lut_mask = 64'h0F7F0F7F0F7F0F7F;
defparam \doing_precharge~0 .shared_arith = "off";

dffeas doing_auto_precharge(
	.clk(ctl_clk),
	.d(\doing_auto_precharge~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\doing_precharge~0_combout ),
	.q(\doing_auto_precharge~q ),
	.prn(vcc));
defparam doing_auto_precharge.is_wysiwyg = "true";
defparam doing_auto_precharge.power_up = "low";

arriaii_lcell_comb \doing_precharge~1 (
	.dataa(!always38),
	.datab(!always106),
	.datac(!always140),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_precharge~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_precharge~1 .extended_lut = "off";
defparam \doing_precharge~1 .lut_mask = 64'h3370337033703370;
defparam \doing_precharge~1 .shared_arith = "off";

dffeas doing_precharge(
	.clk(ctl_clk),
	.d(\doing_precharge~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\doing_precharge~0_combout ),
	.q(\doing_precharge~q ),
	.prn(vcc));
defparam doing_precharge.is_wysiwyg = "true";
defparam doing_precharge.power_up = "low";

arriaii_lcell_comb \int_rdwr_to_valid_ready~0 (
	.dataa(!\doing_read~q ),
	.datab(!\general_counter[0]~q ),
	.datac(!\general_counter[1]~q ),
	.datad(!\doing_auto_precharge~q ),
	.datae(!\general_counter[3]~q ),
	.dataf(!\doing_precharge~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_rdwr_to_valid_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_rdwr_to_valid_ready~0 .extended_lut = "off";
defparam \int_rdwr_to_valid_ready~0 .lut_mask = 64'hA8EA000000000000;
defparam \int_rdwr_to_valid_ready~0 .shared_arith = "off";

arriaii_lcell_comb \int_rdwr_to_valid_ready~1 (
	.dataa(!\general_counter[0]~q ),
	.datab(!\general_counter[1]~q ),
	.datac(!\doing_precharge~q ),
	.datad(!\general_counter[5]~q ),
	.datae(!\general_counter[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_rdwr_to_valid_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_rdwr_to_valid_ready~1 .extended_lut = "off";
defparam \int_rdwr_to_valid_ready~1 .lut_mask = 64'hFE000000FE000000;
defparam \int_rdwr_to_valid_ready~1 .shared_arith = "off";

arriaii_lcell_comb \doing_read~0 (
	.dataa(!do_read_r),
	.datab(!to_chip_r_0),
	.datac(!do_write_r),
	.datad(!Equal0),
	.datae(!\doing_read~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_read~0 .extended_lut = "off";
defparam \doing_read~0 .lut_mask = 64'h0010FFFC0010FFFC;
defparam \doing_read~0 .shared_arith = "off";

dffeas doing_read(
	.clk(ctl_clk),
	.d(\doing_read~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_read~q ),
	.prn(vcc));
defparam doing_read.is_wysiwyg = "true";
defparam doing_read.power_up = "low";

arriaii_lcell_comb \int_rdwr_to_valid_ready~2 (
	.dataa(!act_to_rdwr_1),
	.datab(!\doing_read~q ),
	.datac(!\general_counter[1]~q ),
	.datad(!\doing_auto_precharge~q ),
	.datae(!\general_counter[3]~q ),
	.dataf(!\doing_precharge~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_rdwr_to_valid_ready~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_rdwr_to_valid_ready~2 .extended_lut = "off";
defparam \int_rdwr_to_valid_ready~2 .lut_mask = 64'h54550040FFFF0000;
defparam \int_rdwr_to_valid_ready~2 .shared_arith = "off";

arriaii_lcell_comb \int_rdwr_to_valid_ready~3 (
	.dataa(!close_3_0),
	.datab(!\general_counter[2]~q ),
	.datac(!\int_rdwr_to_valid_ready~0_combout ),
	.datad(!\int_rdwr_to_valid_ready~1_combout ),
	.datae(!\int_rdwr_to_valid_ready~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_rdwr_to_valid_ready~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_rdwr_to_valid_ready~3 .extended_lut = "off";
defparam \int_rdwr_to_valid_ready~3 .lut_mask = 64'h5555551055555510;
defparam \int_rdwr_to_valid_ready~3 .shared_arith = "off";

dffeas int_rdwr_to_valid_ready(
	.clk(ctl_clk),
	.d(\int_rdwr_to_valid_ready~3_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\int_rdwr_to_valid_ready~q ),
	.prn(vcc));
defparam int_rdwr_to_valid_ready.is_wysiwyg = "true";
defparam int_rdwr_to_valid_ready.power_up = "low";

arriaii_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~13 .shared_arith = "off";

arriaii_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \act_counter[4] (
	.clk(ctl_clk),
	.d(\Add0~17_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_3_0),
	.ena(vcc),
	.q(\act_counter[4]~q ),
	.prn(vcc));
defparam \act_counter[4] .is_wysiwyg = "true";
defparam \act_counter[4] .power_up = "low";

arriaii_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \act_counter[5] (
	.clk(ctl_clk),
	.d(\Add0~21_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_3_0),
	.ena(vcc),
	.q(\act_counter[5]~q ),
	.prn(vcc));
defparam \act_counter[5] .is_wysiwyg = "true";
defparam \act_counter[5] .power_up = "low";

arriaii_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Equal0~0_combout ),
	.datae(gnd),
	.dataf(!\act_counter[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF000000FF00;
defparam \Add0~1 .shared_arith = "off";

dffeas \act_counter[0] (
	.clk(ctl_clk),
	.d(\Add0~1_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_3_0),
	.ena(vcc),
	.q(\act_counter[0]~q ),
	.prn(vcc));
defparam \act_counter[0] .is_wysiwyg = "true";
defparam \act_counter[0] .power_up = "low";

arriaii_lcell_comb \Equal0~0 (
	.dataa(!\act_counter[3]~q ),
	.datab(!\act_counter[4]~q ),
	.datac(!\act_counter[5]~q ),
	.datad(!\act_counter[2]~q ),
	.datae(!\act_counter[1]~q ),
	.dataf(!\act_counter[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h0000000000000001;
defparam \Equal0~0 .shared_arith = "off";

arriaii_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \act_counter[1] (
	.clk(ctl_clk),
	.d(\Add0~5_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_3_0),
	.ena(vcc),
	.q(\act_counter[1]~q ),
	.prn(vcc));
defparam \act_counter[1] .is_wysiwyg = "true";
defparam \act_counter[1] .power_up = "low";

arriaii_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \act_counter[2] (
	.clk(ctl_clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_3_0),
	.ena(vcc),
	.q(\act_counter[2]~q ),
	.prn(vcc));
defparam \act_counter[2] .is_wysiwyg = "true";
defparam \act_counter[2] .power_up = "low";

dffeas \act_counter[3] (
	.clk(ctl_clk),
	.d(\Add0~13_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_3_0),
	.ena(vcc),
	.q(\act_counter[3]~q ),
	.prn(vcc));
defparam \act_counter[3] .is_wysiwyg = "true";
defparam \act_counter[3] .power_up = "low";

arriaii_lcell_comb \LessThan0~0 (
	.dataa(!act_to_rdwr_1),
	.datab(!\act_counter[3]~q ),
	.datac(!\act_counter[4]~q ),
	.datad(!\act_counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h4000400040004000;
defparam \LessThan0~0 .shared_arith = "off";

dffeas int_act_to_act_ready(
	.clk(ctl_clk),
	.d(\LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_3_0),
	.ena(vcc),
	.q(\int_act_to_act_ready~q ),
	.prn(vcc));
defparam int_act_to_act_ready.is_wysiwyg = "true";
defparam int_act_to_act_ready.power_up = "low";

arriaii_lcell_comb \rdwr_ready~0 (
	.dataa(!current_state1),
	.datab(!\LessThan0~0_combout ),
	.datac(!\act_counter[2]~q ),
	.datad(!\act_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdwr_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdwr_ready~0 .extended_lut = "off";
defparam \rdwr_ready~0 .lut_mask = 64'h4555455545554555;
defparam \rdwr_ready~0 .shared_arith = "off";

arriaii_lcell_comb \rdwr_ready~1 (
	.dataa(!act_to_rdwr_1),
	.datab(!close_3_0),
	.datac(!open_3_0),
	.datad(!\rdwr_ready~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdwr_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdwr_ready~1 .extended_lut = "off";
defparam \rdwr_ready~1 .lut_mask = 64'h0133013301330133;
defparam \rdwr_ready~1 .shared_arith = "off";

endmodule

module ddr3_int_alt_ddrx_bank_timer_info_4 (
	ctl_clk,
	do_read_r,
	do_write_r,
	current_state1,
	do_precharge_all_r,
	to_chip_r_0,
	always38,
	act_ready1,
	act_to_rdwr_1,
	always106,
	always145,
	ctl_reset_n,
	rdwr_ready1,
	always140,
	Equal0,
	close_4_0,
	open_4_0,
	general_counter,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	ctl_clk;
input 	do_read_r;
input 	do_write_r;
output 	current_state1;
input 	do_precharge_all_r;
input 	to_chip_r_0;
input 	always38;
output 	act_ready1;
input 	act_to_rdwr_1;
input 	always106;
input 	always145;
input 	ctl_reset_n;
output 	rdwr_ready1;
input 	always140;
input 	Equal0;
input 	close_4_0;
input 	open_4_0;
input 	general_counter;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \current_state~0_combout ;
wire \Add1~1_sumout ;
wire \general_counter~1_combout ;
wire \general_counter[0]~q ;
wire \Add1~10 ;
wire \Add1~13_sumout ;
wire \general_counter~3_combout ;
wire \general_counter[3]~q ;
wire \Add1~14 ;
wire \Add1~17_sumout ;
wire \general_counter~5_combout ;
wire \general_counter[4]~q ;
wire \Add1~18 ;
wire \Add1~21_sumout ;
wire \general_counter~4_combout ;
wire \general_counter[5]~q ;
wire \Equal1~0_combout ;
wire \Add1~2 ;
wire \Add1~5_sumout ;
wire \general_counter~2_combout ;
wire \general_counter[1]~q ;
wire \Add1~6 ;
wire \Add1~9_sumout ;
wire \general_counter~0_combout ;
wire \general_counter[2]~q ;
wire \doing_auto_precharge~0_combout ;
wire \doing_precharge~0_combout ;
wire \doing_auto_precharge~q ;
wire \doing_precharge~1_combout ;
wire \doing_precharge~q ;
wire \int_rdwr_to_valid_ready~0_combout ;
wire \int_rdwr_to_valid_ready~1_combout ;
wire \doing_read~0_combout ;
wire \doing_read~q ;
wire \int_rdwr_to_valid_ready~2_combout ;
wire \int_rdwr_to_valid_ready~3_combout ;
wire \int_rdwr_to_valid_ready~q ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \act_counter[4]~q ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \act_counter[5]~q ;
wire \Add0~1_sumout ;
wire \act_counter[0]~q ;
wire \Equal0~0_combout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \act_counter[1]~q ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \act_counter[2]~q ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \act_counter[3]~q ;
wire \LessThan0~0_combout ;
wire \int_act_to_act_ready~q ;
wire \rdwr_ready~0_combout ;
wire \rdwr_ready~1_combout ;


dffeas current_state(
	.clk(ctl_clk),
	.d(\current_state~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_4_0),
	.ena(vcc),
	.q(current_state1),
	.prn(vcc));
defparam current_state.is_wysiwyg = "true";
defparam current_state.power_up = "low";

arriaii_lcell_comb act_ready(
	.dataa(!\int_rdwr_to_valid_ready~q ),
	.datab(!\int_act_to_act_ready~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(act_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam act_ready.extended_lut = "off";
defparam act_ready.lut_mask = 64'h4444444444444444;
defparam act_ready.shared_arith = "off";

dffeas rdwr_ready(
	.clk(ctl_clk),
	.d(\rdwr_ready~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rdwr_ready1),
	.prn(vcc));
defparam rdwr_ready.is_wysiwyg = "true";
defparam rdwr_ready.power_up = "low";

arriaii_lcell_comb \current_state~0 (
	.dataa(!always38),
	.datab(!always106),
	.datac(!current_state1),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\current_state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \current_state~0 .extended_lut = "off";
defparam \current_state~0 .lut_mask = 64'h0C080C080C080C08;
defparam \current_state~0 .shared_arith = "off";

arriaii_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Equal1~0_combout ),
	.datae(gnd),
	.dataf(!\general_counter[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(\Add1~2 ),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h0000FF000000FF00;
defparam \Add1~1 .shared_arith = "off";

arriaii_lcell_comb \general_counter~1 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~1_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~1 .extended_lut = "off";
defparam \general_counter~1 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~1 .shared_arith = "off";

dffeas \general_counter[0] (
	.clk(ctl_clk),
	.d(\general_counter~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[0]~q ),
	.prn(vcc));
defparam \general_counter[0] .is_wysiwyg = "true";
defparam \general_counter[0] .power_up = "low";

arriaii_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~9 .shared_arith = "off";

arriaii_lcell_comb \Add1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~13 .shared_arith = "off";

arriaii_lcell_comb \general_counter~3 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~13_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~3 .extended_lut = "off";
defparam \general_counter~3 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~3 .shared_arith = "off";

dffeas \general_counter[3] (
	.clk(ctl_clk),
	.d(\general_counter~3_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[3]~q ),
	.prn(vcc));
defparam \general_counter[3] .is_wysiwyg = "true";
defparam \general_counter[3] .power_up = "low";

arriaii_lcell_comb \Add1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~17 .shared_arith = "off";

arriaii_lcell_comb \general_counter~5 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~17_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~5 .extended_lut = "off";
defparam \general_counter~5 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~5 .shared_arith = "off";

dffeas \general_counter[4] (
	.clk(ctl_clk),
	.d(\general_counter~5_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[4]~q ),
	.prn(vcc));
defparam \general_counter[4] .is_wysiwyg = "true";
defparam \general_counter[4] .power_up = "low";

arriaii_lcell_comb \Add1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~21_sumout ),
	.cout(),
	.shareout());
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~21 .shared_arith = "off";

arriaii_lcell_comb \general_counter~4 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~21_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~4 .extended_lut = "off";
defparam \general_counter~4 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~4 .shared_arith = "off";

dffeas \general_counter[5] (
	.clk(ctl_clk),
	.d(\general_counter~4_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[5]~q ),
	.prn(vcc));
defparam \general_counter[5] .is_wysiwyg = "true";
defparam \general_counter[5] .power_up = "low";

arriaii_lcell_comb \Equal1~0 (
	.dataa(!\general_counter[2]~q ),
	.datab(!\general_counter[0]~q ),
	.datac(!\general_counter[1]~q ),
	.datad(!\general_counter[3]~q ),
	.datae(!\general_counter[5]~q ),
	.dataf(!\general_counter[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'h0000000000000001;
defparam \Equal1~0 .shared_arith = "off";

arriaii_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~5 .shared_arith = "off";

arriaii_lcell_comb \general_counter~2 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~5_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~2 .extended_lut = "off";
defparam \general_counter~2 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~2 .shared_arith = "off";

dffeas \general_counter[1] (
	.clk(ctl_clk),
	.d(\general_counter~2_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[1]~q ),
	.prn(vcc));
defparam \general_counter[1] .is_wysiwyg = "true";
defparam \general_counter[1] .power_up = "low";

arriaii_lcell_comb \general_counter~0 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~9_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~0 .extended_lut = "off";
defparam \general_counter~0 .lut_mask = 64'h1311FFFF1311FFFF;
defparam \general_counter~0 .shared_arith = "off";

dffeas \general_counter[2] (
	.clk(ctl_clk),
	.d(\general_counter~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[2]~q ),
	.prn(vcc));
defparam \general_counter[2] .is_wysiwyg = "true";
defparam \general_counter[2] .power_up = "low";

arriaii_lcell_comb \doing_auto_precharge~0 (
	.dataa(!always38),
	.datab(!always106),
	.datac(!always140),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_auto_precharge~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_auto_precharge~0 .extended_lut = "off";
defparam \doing_auto_precharge~0 .lut_mask = 64'h0007000700070007;
defparam \doing_auto_precharge~0 .shared_arith = "off";

arriaii_lcell_comb \doing_precharge~0 (
	.dataa(!always38),
	.datab(!always145),
	.datac(!always106),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_precharge~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_precharge~0 .extended_lut = "off";
defparam \doing_precharge~0 .lut_mask = 64'h0F7F0F7F0F7F0F7F;
defparam \doing_precharge~0 .shared_arith = "off";

dffeas doing_auto_precharge(
	.clk(ctl_clk),
	.d(\doing_auto_precharge~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\doing_precharge~0_combout ),
	.q(\doing_auto_precharge~q ),
	.prn(vcc));
defparam doing_auto_precharge.is_wysiwyg = "true";
defparam doing_auto_precharge.power_up = "low";

arriaii_lcell_comb \doing_precharge~1 (
	.dataa(!always38),
	.datab(!always106),
	.datac(!always140),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_precharge~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_precharge~1 .extended_lut = "off";
defparam \doing_precharge~1 .lut_mask = 64'h3370337033703370;
defparam \doing_precharge~1 .shared_arith = "off";

dffeas doing_precharge(
	.clk(ctl_clk),
	.d(\doing_precharge~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\doing_precharge~0_combout ),
	.q(\doing_precharge~q ),
	.prn(vcc));
defparam doing_precharge.is_wysiwyg = "true";
defparam doing_precharge.power_up = "low";

arriaii_lcell_comb \int_rdwr_to_valid_ready~0 (
	.dataa(!\doing_read~q ),
	.datab(!\general_counter[0]~q ),
	.datac(!\general_counter[1]~q ),
	.datad(!\doing_auto_precharge~q ),
	.datae(!\general_counter[3]~q ),
	.dataf(!\doing_precharge~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_rdwr_to_valid_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_rdwr_to_valid_ready~0 .extended_lut = "off";
defparam \int_rdwr_to_valid_ready~0 .lut_mask = 64'hA8EA000000000000;
defparam \int_rdwr_to_valid_ready~0 .shared_arith = "off";

arriaii_lcell_comb \int_rdwr_to_valid_ready~1 (
	.dataa(!\general_counter[0]~q ),
	.datab(!\general_counter[1]~q ),
	.datac(!\doing_precharge~q ),
	.datad(!\general_counter[5]~q ),
	.datae(!\general_counter[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_rdwr_to_valid_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_rdwr_to_valid_ready~1 .extended_lut = "off";
defparam \int_rdwr_to_valid_ready~1 .lut_mask = 64'hFE000000FE000000;
defparam \int_rdwr_to_valid_ready~1 .shared_arith = "off";

arriaii_lcell_comb \doing_read~0 (
	.dataa(!do_read_r),
	.datab(!to_chip_r_0),
	.datac(!do_write_r),
	.datad(!Equal0),
	.datae(!\doing_read~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_read~0 .extended_lut = "off";
defparam \doing_read~0 .lut_mask = 64'h0010FFFC0010FFFC;
defparam \doing_read~0 .shared_arith = "off";

dffeas doing_read(
	.clk(ctl_clk),
	.d(\doing_read~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_read~q ),
	.prn(vcc));
defparam doing_read.is_wysiwyg = "true";
defparam doing_read.power_up = "low";

arriaii_lcell_comb \int_rdwr_to_valid_ready~2 (
	.dataa(!act_to_rdwr_1),
	.datab(!\doing_read~q ),
	.datac(!\general_counter[1]~q ),
	.datad(!\doing_auto_precharge~q ),
	.datae(!\general_counter[3]~q ),
	.dataf(!\doing_precharge~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_rdwr_to_valid_ready~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_rdwr_to_valid_ready~2 .extended_lut = "off";
defparam \int_rdwr_to_valid_ready~2 .lut_mask = 64'h54550040FFFF0000;
defparam \int_rdwr_to_valid_ready~2 .shared_arith = "off";

arriaii_lcell_comb \int_rdwr_to_valid_ready~3 (
	.dataa(!close_4_0),
	.datab(!\general_counter[2]~q ),
	.datac(!\int_rdwr_to_valid_ready~0_combout ),
	.datad(!\int_rdwr_to_valid_ready~1_combout ),
	.datae(!\int_rdwr_to_valid_ready~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_rdwr_to_valid_ready~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_rdwr_to_valid_ready~3 .extended_lut = "off";
defparam \int_rdwr_to_valid_ready~3 .lut_mask = 64'h5555551055555510;
defparam \int_rdwr_to_valid_ready~3 .shared_arith = "off";

dffeas int_rdwr_to_valid_ready(
	.clk(ctl_clk),
	.d(\int_rdwr_to_valid_ready~3_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\int_rdwr_to_valid_ready~q ),
	.prn(vcc));
defparam int_rdwr_to_valid_ready.is_wysiwyg = "true";
defparam int_rdwr_to_valid_ready.power_up = "low";

arriaii_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~13 .shared_arith = "off";

arriaii_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \act_counter[4] (
	.clk(ctl_clk),
	.d(\Add0~17_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_4_0),
	.ena(vcc),
	.q(\act_counter[4]~q ),
	.prn(vcc));
defparam \act_counter[4] .is_wysiwyg = "true";
defparam \act_counter[4] .power_up = "low";

arriaii_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \act_counter[5] (
	.clk(ctl_clk),
	.d(\Add0~21_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_4_0),
	.ena(vcc),
	.q(\act_counter[5]~q ),
	.prn(vcc));
defparam \act_counter[5] .is_wysiwyg = "true";
defparam \act_counter[5] .power_up = "low";

arriaii_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Equal0~0_combout ),
	.datae(gnd),
	.dataf(!\act_counter[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF000000FF00;
defparam \Add0~1 .shared_arith = "off";

dffeas \act_counter[0] (
	.clk(ctl_clk),
	.d(\Add0~1_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_4_0),
	.ena(vcc),
	.q(\act_counter[0]~q ),
	.prn(vcc));
defparam \act_counter[0] .is_wysiwyg = "true";
defparam \act_counter[0] .power_up = "low";

arriaii_lcell_comb \Equal0~0 (
	.dataa(!\act_counter[3]~q ),
	.datab(!\act_counter[4]~q ),
	.datac(!\act_counter[5]~q ),
	.datad(!\act_counter[2]~q ),
	.datae(!\act_counter[1]~q ),
	.dataf(!\act_counter[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h0000000000000001;
defparam \Equal0~0 .shared_arith = "off";

arriaii_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \act_counter[1] (
	.clk(ctl_clk),
	.d(\Add0~5_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_4_0),
	.ena(vcc),
	.q(\act_counter[1]~q ),
	.prn(vcc));
defparam \act_counter[1] .is_wysiwyg = "true";
defparam \act_counter[1] .power_up = "low";

arriaii_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \act_counter[2] (
	.clk(ctl_clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_4_0),
	.ena(vcc),
	.q(\act_counter[2]~q ),
	.prn(vcc));
defparam \act_counter[2] .is_wysiwyg = "true";
defparam \act_counter[2] .power_up = "low";

dffeas \act_counter[3] (
	.clk(ctl_clk),
	.d(\Add0~13_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_4_0),
	.ena(vcc),
	.q(\act_counter[3]~q ),
	.prn(vcc));
defparam \act_counter[3] .is_wysiwyg = "true";
defparam \act_counter[3] .power_up = "low";

arriaii_lcell_comb \LessThan0~0 (
	.dataa(!act_to_rdwr_1),
	.datab(!\act_counter[3]~q ),
	.datac(!\act_counter[4]~q ),
	.datad(!\act_counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h4000400040004000;
defparam \LessThan0~0 .shared_arith = "off";

dffeas int_act_to_act_ready(
	.clk(ctl_clk),
	.d(\LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_4_0),
	.ena(vcc),
	.q(\int_act_to_act_ready~q ),
	.prn(vcc));
defparam int_act_to_act_ready.is_wysiwyg = "true";
defparam int_act_to_act_ready.power_up = "low";

arriaii_lcell_comb \rdwr_ready~0 (
	.dataa(!current_state1),
	.datab(!\LessThan0~0_combout ),
	.datac(!\act_counter[2]~q ),
	.datad(!\act_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdwr_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdwr_ready~0 .extended_lut = "off";
defparam \rdwr_ready~0 .lut_mask = 64'h4555455545554555;
defparam \rdwr_ready~0 .shared_arith = "off";

arriaii_lcell_comb \rdwr_ready~1 (
	.dataa(!act_to_rdwr_1),
	.datab(!close_4_0),
	.datac(!open_4_0),
	.datad(!\rdwr_ready~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdwr_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdwr_ready~1 .extended_lut = "off";
defparam \rdwr_ready~1 .lut_mask = 64'h0133013301330133;
defparam \rdwr_ready~1 .shared_arith = "off";

endmodule

module ddr3_int_alt_ddrx_bank_timer_info_5 (
	ctl_clk,
	do_read_r,
	do_write_r,
	current_state1,
	do_precharge_all_r,
	to_chip_r_0,
	always38,
	act_ready1,
	act_to_rdwr_1,
	always106,
	always145,
	ctl_reset_n,
	rdwr_ready1,
	always140,
	Equal0,
	close_5_0,
	open_5_0,
	general_counter,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	ctl_clk;
input 	do_read_r;
input 	do_write_r;
output 	current_state1;
input 	do_precharge_all_r;
input 	to_chip_r_0;
input 	always38;
output 	act_ready1;
input 	act_to_rdwr_1;
input 	always106;
input 	always145;
input 	ctl_reset_n;
output 	rdwr_ready1;
input 	always140;
input 	Equal0;
input 	close_5_0;
input 	open_5_0;
input 	general_counter;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \current_state~0_combout ;
wire \Add1~1_sumout ;
wire \general_counter~1_combout ;
wire \general_counter[0]~q ;
wire \Add1~10 ;
wire \Add1~13_sumout ;
wire \general_counter~3_combout ;
wire \general_counter[3]~q ;
wire \Add1~14 ;
wire \Add1~17_sumout ;
wire \general_counter~5_combout ;
wire \general_counter[4]~q ;
wire \Add1~18 ;
wire \Add1~21_sumout ;
wire \general_counter~4_combout ;
wire \general_counter[5]~q ;
wire \Equal1~0_combout ;
wire \Add1~2 ;
wire \Add1~5_sumout ;
wire \general_counter~2_combout ;
wire \general_counter[1]~q ;
wire \Add1~6 ;
wire \Add1~9_sumout ;
wire \general_counter~0_combout ;
wire \general_counter[2]~q ;
wire \doing_auto_precharge~0_combout ;
wire \doing_precharge~0_combout ;
wire \doing_auto_precharge~q ;
wire \doing_precharge~1_combout ;
wire \doing_precharge~q ;
wire \int_rdwr_to_valid_ready~0_combout ;
wire \int_rdwr_to_valid_ready~1_combout ;
wire \doing_read~0_combout ;
wire \doing_read~q ;
wire \int_rdwr_to_valid_ready~2_combout ;
wire \int_rdwr_to_valid_ready~3_combout ;
wire \int_rdwr_to_valid_ready~q ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \act_counter[4]~q ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \act_counter[5]~q ;
wire \Add0~1_sumout ;
wire \act_counter[0]~q ;
wire \Equal0~0_combout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \act_counter[1]~q ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \act_counter[2]~q ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \act_counter[3]~q ;
wire \LessThan0~0_combout ;
wire \int_act_to_act_ready~q ;
wire \rdwr_ready~0_combout ;
wire \rdwr_ready~1_combout ;


dffeas current_state(
	.clk(ctl_clk),
	.d(\current_state~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_5_0),
	.ena(vcc),
	.q(current_state1),
	.prn(vcc));
defparam current_state.is_wysiwyg = "true";
defparam current_state.power_up = "low";

arriaii_lcell_comb act_ready(
	.dataa(!\int_rdwr_to_valid_ready~q ),
	.datab(!\int_act_to_act_ready~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(act_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam act_ready.extended_lut = "off";
defparam act_ready.lut_mask = 64'h4444444444444444;
defparam act_ready.shared_arith = "off";

dffeas rdwr_ready(
	.clk(ctl_clk),
	.d(\rdwr_ready~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rdwr_ready1),
	.prn(vcc));
defparam rdwr_ready.is_wysiwyg = "true";
defparam rdwr_ready.power_up = "low";

arriaii_lcell_comb \current_state~0 (
	.dataa(!always38),
	.datab(!always106),
	.datac(!current_state1),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\current_state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \current_state~0 .extended_lut = "off";
defparam \current_state~0 .lut_mask = 64'h0C080C080C080C08;
defparam \current_state~0 .shared_arith = "off";

arriaii_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Equal1~0_combout ),
	.datae(gnd),
	.dataf(!\general_counter[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(\Add1~2 ),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h0000FF000000FF00;
defparam \Add1~1 .shared_arith = "off";

arriaii_lcell_comb \general_counter~1 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~1_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~1 .extended_lut = "off";
defparam \general_counter~1 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~1 .shared_arith = "off";

dffeas \general_counter[0] (
	.clk(ctl_clk),
	.d(\general_counter~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[0]~q ),
	.prn(vcc));
defparam \general_counter[0] .is_wysiwyg = "true";
defparam \general_counter[0] .power_up = "low";

arriaii_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~9 .shared_arith = "off";

arriaii_lcell_comb \Add1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~13 .shared_arith = "off";

arriaii_lcell_comb \general_counter~3 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~13_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~3 .extended_lut = "off";
defparam \general_counter~3 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~3 .shared_arith = "off";

dffeas \general_counter[3] (
	.clk(ctl_clk),
	.d(\general_counter~3_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[3]~q ),
	.prn(vcc));
defparam \general_counter[3] .is_wysiwyg = "true";
defparam \general_counter[3] .power_up = "low";

arriaii_lcell_comb \Add1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~17 .shared_arith = "off";

arriaii_lcell_comb \general_counter~5 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~17_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~5 .extended_lut = "off";
defparam \general_counter~5 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~5 .shared_arith = "off";

dffeas \general_counter[4] (
	.clk(ctl_clk),
	.d(\general_counter~5_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[4]~q ),
	.prn(vcc));
defparam \general_counter[4] .is_wysiwyg = "true";
defparam \general_counter[4] .power_up = "low";

arriaii_lcell_comb \Add1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~21_sumout ),
	.cout(),
	.shareout());
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~21 .shared_arith = "off";

arriaii_lcell_comb \general_counter~4 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~21_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~4 .extended_lut = "off";
defparam \general_counter~4 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~4 .shared_arith = "off";

dffeas \general_counter[5] (
	.clk(ctl_clk),
	.d(\general_counter~4_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[5]~q ),
	.prn(vcc));
defparam \general_counter[5] .is_wysiwyg = "true";
defparam \general_counter[5] .power_up = "low";

arriaii_lcell_comb \Equal1~0 (
	.dataa(!\general_counter[2]~q ),
	.datab(!\general_counter[0]~q ),
	.datac(!\general_counter[1]~q ),
	.datad(!\general_counter[3]~q ),
	.datae(!\general_counter[5]~q ),
	.dataf(!\general_counter[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'h0000000000000001;
defparam \Equal1~0 .shared_arith = "off";

arriaii_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~5 .shared_arith = "off";

arriaii_lcell_comb \general_counter~2 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~5_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~2 .extended_lut = "off";
defparam \general_counter~2 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~2 .shared_arith = "off";

dffeas \general_counter[1] (
	.clk(ctl_clk),
	.d(\general_counter~2_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[1]~q ),
	.prn(vcc));
defparam \general_counter[1] .is_wysiwyg = "true";
defparam \general_counter[1] .power_up = "low";

arriaii_lcell_comb \general_counter~0 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~9_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~0 .extended_lut = "off";
defparam \general_counter~0 .lut_mask = 64'h1311FFFF1311FFFF;
defparam \general_counter~0 .shared_arith = "off";

dffeas \general_counter[2] (
	.clk(ctl_clk),
	.d(\general_counter~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[2]~q ),
	.prn(vcc));
defparam \general_counter[2] .is_wysiwyg = "true";
defparam \general_counter[2] .power_up = "low";

arriaii_lcell_comb \doing_auto_precharge~0 (
	.dataa(!always38),
	.datab(!always106),
	.datac(!always140),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_auto_precharge~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_auto_precharge~0 .extended_lut = "off";
defparam \doing_auto_precharge~0 .lut_mask = 64'h0007000700070007;
defparam \doing_auto_precharge~0 .shared_arith = "off";

arriaii_lcell_comb \doing_precharge~0 (
	.dataa(!always38),
	.datab(!always145),
	.datac(!always106),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_precharge~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_precharge~0 .extended_lut = "off";
defparam \doing_precharge~0 .lut_mask = 64'h0F7F0F7F0F7F0F7F;
defparam \doing_precharge~0 .shared_arith = "off";

dffeas doing_auto_precharge(
	.clk(ctl_clk),
	.d(\doing_auto_precharge~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\doing_precharge~0_combout ),
	.q(\doing_auto_precharge~q ),
	.prn(vcc));
defparam doing_auto_precharge.is_wysiwyg = "true";
defparam doing_auto_precharge.power_up = "low";

arriaii_lcell_comb \doing_precharge~1 (
	.dataa(!always38),
	.datab(!always106),
	.datac(!always140),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_precharge~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_precharge~1 .extended_lut = "off";
defparam \doing_precharge~1 .lut_mask = 64'h3370337033703370;
defparam \doing_precharge~1 .shared_arith = "off";

dffeas doing_precharge(
	.clk(ctl_clk),
	.d(\doing_precharge~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\doing_precharge~0_combout ),
	.q(\doing_precharge~q ),
	.prn(vcc));
defparam doing_precharge.is_wysiwyg = "true";
defparam doing_precharge.power_up = "low";

arriaii_lcell_comb \int_rdwr_to_valid_ready~0 (
	.dataa(!\doing_read~q ),
	.datab(!\general_counter[0]~q ),
	.datac(!\general_counter[1]~q ),
	.datad(!\doing_auto_precharge~q ),
	.datae(!\general_counter[3]~q ),
	.dataf(!\doing_precharge~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_rdwr_to_valid_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_rdwr_to_valid_ready~0 .extended_lut = "off";
defparam \int_rdwr_to_valid_ready~0 .lut_mask = 64'hA8EA000000000000;
defparam \int_rdwr_to_valid_ready~0 .shared_arith = "off";

arriaii_lcell_comb \int_rdwr_to_valid_ready~1 (
	.dataa(!\general_counter[0]~q ),
	.datab(!\general_counter[1]~q ),
	.datac(!\doing_precharge~q ),
	.datad(!\general_counter[5]~q ),
	.datae(!\general_counter[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_rdwr_to_valid_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_rdwr_to_valid_ready~1 .extended_lut = "off";
defparam \int_rdwr_to_valid_ready~1 .lut_mask = 64'hFE000000FE000000;
defparam \int_rdwr_to_valid_ready~1 .shared_arith = "off";

arriaii_lcell_comb \doing_read~0 (
	.dataa(!do_read_r),
	.datab(!to_chip_r_0),
	.datac(!do_write_r),
	.datad(!Equal0),
	.datae(!\doing_read~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_read~0 .extended_lut = "off";
defparam \doing_read~0 .lut_mask = 64'h0010FFFC0010FFFC;
defparam \doing_read~0 .shared_arith = "off";

dffeas doing_read(
	.clk(ctl_clk),
	.d(\doing_read~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_read~q ),
	.prn(vcc));
defparam doing_read.is_wysiwyg = "true";
defparam doing_read.power_up = "low";

arriaii_lcell_comb \int_rdwr_to_valid_ready~2 (
	.dataa(!act_to_rdwr_1),
	.datab(!\doing_read~q ),
	.datac(!\general_counter[1]~q ),
	.datad(!\doing_auto_precharge~q ),
	.datae(!\general_counter[3]~q ),
	.dataf(!\doing_precharge~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_rdwr_to_valid_ready~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_rdwr_to_valid_ready~2 .extended_lut = "off";
defparam \int_rdwr_to_valid_ready~2 .lut_mask = 64'h54550040FFFF0000;
defparam \int_rdwr_to_valid_ready~2 .shared_arith = "off";

arriaii_lcell_comb \int_rdwr_to_valid_ready~3 (
	.dataa(!close_5_0),
	.datab(!\general_counter[2]~q ),
	.datac(!\int_rdwr_to_valid_ready~0_combout ),
	.datad(!\int_rdwr_to_valid_ready~1_combout ),
	.datae(!\int_rdwr_to_valid_ready~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_rdwr_to_valid_ready~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_rdwr_to_valid_ready~3 .extended_lut = "off";
defparam \int_rdwr_to_valid_ready~3 .lut_mask = 64'h5555551055555510;
defparam \int_rdwr_to_valid_ready~3 .shared_arith = "off";

dffeas int_rdwr_to_valid_ready(
	.clk(ctl_clk),
	.d(\int_rdwr_to_valid_ready~3_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\int_rdwr_to_valid_ready~q ),
	.prn(vcc));
defparam int_rdwr_to_valid_ready.is_wysiwyg = "true";
defparam int_rdwr_to_valid_ready.power_up = "low";

arriaii_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~13 .shared_arith = "off";

arriaii_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \act_counter[4] (
	.clk(ctl_clk),
	.d(\Add0~17_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_5_0),
	.ena(vcc),
	.q(\act_counter[4]~q ),
	.prn(vcc));
defparam \act_counter[4] .is_wysiwyg = "true";
defparam \act_counter[4] .power_up = "low";

arriaii_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \act_counter[5] (
	.clk(ctl_clk),
	.d(\Add0~21_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_5_0),
	.ena(vcc),
	.q(\act_counter[5]~q ),
	.prn(vcc));
defparam \act_counter[5] .is_wysiwyg = "true";
defparam \act_counter[5] .power_up = "low";

arriaii_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Equal0~0_combout ),
	.datae(gnd),
	.dataf(!\act_counter[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF000000FF00;
defparam \Add0~1 .shared_arith = "off";

dffeas \act_counter[0] (
	.clk(ctl_clk),
	.d(\Add0~1_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_5_0),
	.ena(vcc),
	.q(\act_counter[0]~q ),
	.prn(vcc));
defparam \act_counter[0] .is_wysiwyg = "true";
defparam \act_counter[0] .power_up = "low";

arriaii_lcell_comb \Equal0~0 (
	.dataa(!\act_counter[3]~q ),
	.datab(!\act_counter[4]~q ),
	.datac(!\act_counter[5]~q ),
	.datad(!\act_counter[2]~q ),
	.datae(!\act_counter[1]~q ),
	.dataf(!\act_counter[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h0000000000000001;
defparam \Equal0~0 .shared_arith = "off";

arriaii_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \act_counter[1] (
	.clk(ctl_clk),
	.d(\Add0~5_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_5_0),
	.ena(vcc),
	.q(\act_counter[1]~q ),
	.prn(vcc));
defparam \act_counter[1] .is_wysiwyg = "true";
defparam \act_counter[1] .power_up = "low";

arriaii_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \act_counter[2] (
	.clk(ctl_clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_5_0),
	.ena(vcc),
	.q(\act_counter[2]~q ),
	.prn(vcc));
defparam \act_counter[2] .is_wysiwyg = "true";
defparam \act_counter[2] .power_up = "low";

dffeas \act_counter[3] (
	.clk(ctl_clk),
	.d(\Add0~13_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_5_0),
	.ena(vcc),
	.q(\act_counter[3]~q ),
	.prn(vcc));
defparam \act_counter[3] .is_wysiwyg = "true";
defparam \act_counter[3] .power_up = "low";

arriaii_lcell_comb \LessThan0~0 (
	.dataa(!act_to_rdwr_1),
	.datab(!\act_counter[3]~q ),
	.datac(!\act_counter[4]~q ),
	.datad(!\act_counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h4000400040004000;
defparam \LessThan0~0 .shared_arith = "off";

dffeas int_act_to_act_ready(
	.clk(ctl_clk),
	.d(\LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_5_0),
	.ena(vcc),
	.q(\int_act_to_act_ready~q ),
	.prn(vcc));
defparam int_act_to_act_ready.is_wysiwyg = "true";
defparam int_act_to_act_ready.power_up = "low";

arriaii_lcell_comb \rdwr_ready~0 (
	.dataa(!current_state1),
	.datab(!\LessThan0~0_combout ),
	.datac(!\act_counter[2]~q ),
	.datad(!\act_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdwr_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdwr_ready~0 .extended_lut = "off";
defparam \rdwr_ready~0 .lut_mask = 64'h4555455545554555;
defparam \rdwr_ready~0 .shared_arith = "off";

arriaii_lcell_comb \rdwr_ready~1 (
	.dataa(!act_to_rdwr_1),
	.datab(!close_5_0),
	.datac(!open_5_0),
	.datad(!\rdwr_ready~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdwr_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdwr_ready~1 .extended_lut = "off";
defparam \rdwr_ready~1 .lut_mask = 64'h0133013301330133;
defparam \rdwr_ready~1 .shared_arith = "off";

endmodule

module ddr3_int_alt_ddrx_bank_timer_info_6 (
	ctl_clk,
	do_read_r,
	do_write_r,
	current_state1,
	do_precharge_all_r,
	to_chip_r_0,
	always38,
	act_ready1,
	act_to_rdwr_1,
	always106,
	always145,
	ctl_reset_n,
	rdwr_ready1,
	always140,
	Equal0,
	close_6_0,
	open_6_0,
	general_counter,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	ctl_clk;
input 	do_read_r;
input 	do_write_r;
output 	current_state1;
input 	do_precharge_all_r;
input 	to_chip_r_0;
input 	always38;
output 	act_ready1;
input 	act_to_rdwr_1;
input 	always106;
input 	always145;
input 	ctl_reset_n;
output 	rdwr_ready1;
input 	always140;
input 	Equal0;
input 	close_6_0;
input 	open_6_0;
input 	general_counter;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \current_state~0_combout ;
wire \Add1~1_sumout ;
wire \general_counter~1_combout ;
wire \general_counter[0]~q ;
wire \Add1~10 ;
wire \Add1~13_sumout ;
wire \general_counter~3_combout ;
wire \general_counter[3]~q ;
wire \Add1~14 ;
wire \Add1~17_sumout ;
wire \general_counter~5_combout ;
wire \general_counter[4]~q ;
wire \Add1~18 ;
wire \Add1~21_sumout ;
wire \general_counter~4_combout ;
wire \general_counter[5]~q ;
wire \Equal1~0_combout ;
wire \Add1~2 ;
wire \Add1~5_sumout ;
wire \general_counter~2_combout ;
wire \general_counter[1]~q ;
wire \Add1~6 ;
wire \Add1~9_sumout ;
wire \general_counter~0_combout ;
wire \general_counter[2]~q ;
wire \doing_auto_precharge~0_combout ;
wire \doing_precharge~0_combout ;
wire \doing_auto_precharge~q ;
wire \doing_precharge~1_combout ;
wire \doing_precharge~q ;
wire \int_rdwr_to_valid_ready~0_combout ;
wire \int_rdwr_to_valid_ready~1_combout ;
wire \doing_read~0_combout ;
wire \doing_read~q ;
wire \int_rdwr_to_valid_ready~2_combout ;
wire \int_rdwr_to_valid_ready~3_combout ;
wire \int_rdwr_to_valid_ready~q ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \act_counter[4]~q ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \act_counter[5]~q ;
wire \Add0~1_sumout ;
wire \act_counter[0]~q ;
wire \Equal0~0_combout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \act_counter[1]~q ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \act_counter[2]~q ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \act_counter[3]~q ;
wire \LessThan0~0_combout ;
wire \int_act_to_act_ready~q ;
wire \rdwr_ready~0_combout ;
wire \rdwr_ready~1_combout ;


dffeas current_state(
	.clk(ctl_clk),
	.d(\current_state~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_6_0),
	.ena(vcc),
	.q(current_state1),
	.prn(vcc));
defparam current_state.is_wysiwyg = "true";
defparam current_state.power_up = "low";

arriaii_lcell_comb act_ready(
	.dataa(!\int_rdwr_to_valid_ready~q ),
	.datab(!\int_act_to_act_ready~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(act_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam act_ready.extended_lut = "off";
defparam act_ready.lut_mask = 64'h4444444444444444;
defparam act_ready.shared_arith = "off";

dffeas rdwr_ready(
	.clk(ctl_clk),
	.d(\rdwr_ready~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rdwr_ready1),
	.prn(vcc));
defparam rdwr_ready.is_wysiwyg = "true";
defparam rdwr_ready.power_up = "low";

arriaii_lcell_comb \current_state~0 (
	.dataa(!always38),
	.datab(!always106),
	.datac(!current_state1),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\current_state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \current_state~0 .extended_lut = "off";
defparam \current_state~0 .lut_mask = 64'h0C080C080C080C08;
defparam \current_state~0 .shared_arith = "off";

arriaii_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Equal1~0_combout ),
	.datae(gnd),
	.dataf(!\general_counter[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(\Add1~2 ),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h0000FF000000FF00;
defparam \Add1~1 .shared_arith = "off";

arriaii_lcell_comb \general_counter~1 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~1_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~1 .extended_lut = "off";
defparam \general_counter~1 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~1 .shared_arith = "off";

dffeas \general_counter[0] (
	.clk(ctl_clk),
	.d(\general_counter~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[0]~q ),
	.prn(vcc));
defparam \general_counter[0] .is_wysiwyg = "true";
defparam \general_counter[0] .power_up = "low";

arriaii_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~9 .shared_arith = "off";

arriaii_lcell_comb \Add1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~13 .shared_arith = "off";

arriaii_lcell_comb \general_counter~3 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~13_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~3 .extended_lut = "off";
defparam \general_counter~3 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~3 .shared_arith = "off";

dffeas \general_counter[3] (
	.clk(ctl_clk),
	.d(\general_counter~3_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[3]~q ),
	.prn(vcc));
defparam \general_counter[3] .is_wysiwyg = "true";
defparam \general_counter[3] .power_up = "low";

arriaii_lcell_comb \Add1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~17 .shared_arith = "off";

arriaii_lcell_comb \general_counter~5 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~17_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~5 .extended_lut = "off";
defparam \general_counter~5 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~5 .shared_arith = "off";

dffeas \general_counter[4] (
	.clk(ctl_clk),
	.d(\general_counter~5_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[4]~q ),
	.prn(vcc));
defparam \general_counter[4] .is_wysiwyg = "true";
defparam \general_counter[4] .power_up = "low";

arriaii_lcell_comb \Add1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~21_sumout ),
	.cout(),
	.shareout());
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~21 .shared_arith = "off";

arriaii_lcell_comb \general_counter~4 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~21_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~4 .extended_lut = "off";
defparam \general_counter~4 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~4 .shared_arith = "off";

dffeas \general_counter[5] (
	.clk(ctl_clk),
	.d(\general_counter~4_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[5]~q ),
	.prn(vcc));
defparam \general_counter[5] .is_wysiwyg = "true";
defparam \general_counter[5] .power_up = "low";

arriaii_lcell_comb \Equal1~0 (
	.dataa(!\general_counter[2]~q ),
	.datab(!\general_counter[0]~q ),
	.datac(!\general_counter[1]~q ),
	.datad(!\general_counter[3]~q ),
	.datae(!\general_counter[5]~q ),
	.dataf(!\general_counter[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'h0000000000000001;
defparam \Equal1~0 .shared_arith = "off";

arriaii_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~5 .shared_arith = "off";

arriaii_lcell_comb \general_counter~2 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~5_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~2 .extended_lut = "off";
defparam \general_counter~2 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~2 .shared_arith = "off";

dffeas \general_counter[1] (
	.clk(ctl_clk),
	.d(\general_counter~2_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[1]~q ),
	.prn(vcc));
defparam \general_counter[1] .is_wysiwyg = "true";
defparam \general_counter[1] .power_up = "low";

arriaii_lcell_comb \general_counter~0 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~9_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~0 .extended_lut = "off";
defparam \general_counter~0 .lut_mask = 64'h1311FFFF1311FFFF;
defparam \general_counter~0 .shared_arith = "off";

dffeas \general_counter[2] (
	.clk(ctl_clk),
	.d(\general_counter~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[2]~q ),
	.prn(vcc));
defparam \general_counter[2] .is_wysiwyg = "true";
defparam \general_counter[2] .power_up = "low";

arriaii_lcell_comb \doing_auto_precharge~0 (
	.dataa(!always38),
	.datab(!always106),
	.datac(!always140),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_auto_precharge~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_auto_precharge~0 .extended_lut = "off";
defparam \doing_auto_precharge~0 .lut_mask = 64'h0007000700070007;
defparam \doing_auto_precharge~0 .shared_arith = "off";

arriaii_lcell_comb \doing_precharge~0 (
	.dataa(!always38),
	.datab(!always145),
	.datac(!always106),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_precharge~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_precharge~0 .extended_lut = "off";
defparam \doing_precharge~0 .lut_mask = 64'h0F7F0F7F0F7F0F7F;
defparam \doing_precharge~0 .shared_arith = "off";

dffeas doing_auto_precharge(
	.clk(ctl_clk),
	.d(\doing_auto_precharge~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\doing_precharge~0_combout ),
	.q(\doing_auto_precharge~q ),
	.prn(vcc));
defparam doing_auto_precharge.is_wysiwyg = "true";
defparam doing_auto_precharge.power_up = "low";

arriaii_lcell_comb \doing_precharge~1 (
	.dataa(!always38),
	.datab(!always106),
	.datac(!always140),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_precharge~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_precharge~1 .extended_lut = "off";
defparam \doing_precharge~1 .lut_mask = 64'h3370337033703370;
defparam \doing_precharge~1 .shared_arith = "off";

dffeas doing_precharge(
	.clk(ctl_clk),
	.d(\doing_precharge~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\doing_precharge~0_combout ),
	.q(\doing_precharge~q ),
	.prn(vcc));
defparam doing_precharge.is_wysiwyg = "true";
defparam doing_precharge.power_up = "low";

arriaii_lcell_comb \int_rdwr_to_valid_ready~0 (
	.dataa(!\doing_read~q ),
	.datab(!\general_counter[0]~q ),
	.datac(!\general_counter[1]~q ),
	.datad(!\doing_auto_precharge~q ),
	.datae(!\general_counter[3]~q ),
	.dataf(!\doing_precharge~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_rdwr_to_valid_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_rdwr_to_valid_ready~0 .extended_lut = "off";
defparam \int_rdwr_to_valid_ready~0 .lut_mask = 64'hA8EA000000000000;
defparam \int_rdwr_to_valid_ready~0 .shared_arith = "off";

arriaii_lcell_comb \int_rdwr_to_valid_ready~1 (
	.dataa(!\general_counter[0]~q ),
	.datab(!\general_counter[1]~q ),
	.datac(!\doing_precharge~q ),
	.datad(!\general_counter[5]~q ),
	.datae(!\general_counter[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_rdwr_to_valid_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_rdwr_to_valid_ready~1 .extended_lut = "off";
defparam \int_rdwr_to_valid_ready~1 .lut_mask = 64'hFE000000FE000000;
defparam \int_rdwr_to_valid_ready~1 .shared_arith = "off";

arriaii_lcell_comb \doing_read~0 (
	.dataa(!do_read_r),
	.datab(!to_chip_r_0),
	.datac(!do_write_r),
	.datad(!Equal0),
	.datae(!\doing_read~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_read~0 .extended_lut = "off";
defparam \doing_read~0 .lut_mask = 64'h0010FFFC0010FFFC;
defparam \doing_read~0 .shared_arith = "off";

dffeas doing_read(
	.clk(ctl_clk),
	.d(\doing_read~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_read~q ),
	.prn(vcc));
defparam doing_read.is_wysiwyg = "true";
defparam doing_read.power_up = "low";

arriaii_lcell_comb \int_rdwr_to_valid_ready~2 (
	.dataa(!act_to_rdwr_1),
	.datab(!\doing_read~q ),
	.datac(!\general_counter[1]~q ),
	.datad(!\doing_auto_precharge~q ),
	.datae(!\general_counter[3]~q ),
	.dataf(!\doing_precharge~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_rdwr_to_valid_ready~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_rdwr_to_valid_ready~2 .extended_lut = "off";
defparam \int_rdwr_to_valid_ready~2 .lut_mask = 64'h54550040FFFF0000;
defparam \int_rdwr_to_valid_ready~2 .shared_arith = "off";

arriaii_lcell_comb \int_rdwr_to_valid_ready~3 (
	.dataa(!close_6_0),
	.datab(!\general_counter[2]~q ),
	.datac(!\int_rdwr_to_valid_ready~0_combout ),
	.datad(!\int_rdwr_to_valid_ready~1_combout ),
	.datae(!\int_rdwr_to_valid_ready~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_rdwr_to_valid_ready~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_rdwr_to_valid_ready~3 .extended_lut = "off";
defparam \int_rdwr_to_valid_ready~3 .lut_mask = 64'h5555551055555510;
defparam \int_rdwr_to_valid_ready~3 .shared_arith = "off";

dffeas int_rdwr_to_valid_ready(
	.clk(ctl_clk),
	.d(\int_rdwr_to_valid_ready~3_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\int_rdwr_to_valid_ready~q ),
	.prn(vcc));
defparam int_rdwr_to_valid_ready.is_wysiwyg = "true";
defparam int_rdwr_to_valid_ready.power_up = "low";

arriaii_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~13 .shared_arith = "off";

arriaii_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \act_counter[4] (
	.clk(ctl_clk),
	.d(\Add0~17_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_6_0),
	.ena(vcc),
	.q(\act_counter[4]~q ),
	.prn(vcc));
defparam \act_counter[4] .is_wysiwyg = "true";
defparam \act_counter[4] .power_up = "low";

arriaii_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \act_counter[5] (
	.clk(ctl_clk),
	.d(\Add0~21_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_6_0),
	.ena(vcc),
	.q(\act_counter[5]~q ),
	.prn(vcc));
defparam \act_counter[5] .is_wysiwyg = "true";
defparam \act_counter[5] .power_up = "low";

arriaii_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Equal0~0_combout ),
	.datae(gnd),
	.dataf(!\act_counter[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF000000FF00;
defparam \Add0~1 .shared_arith = "off";

dffeas \act_counter[0] (
	.clk(ctl_clk),
	.d(\Add0~1_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_6_0),
	.ena(vcc),
	.q(\act_counter[0]~q ),
	.prn(vcc));
defparam \act_counter[0] .is_wysiwyg = "true";
defparam \act_counter[0] .power_up = "low";

arriaii_lcell_comb \Equal0~0 (
	.dataa(!\act_counter[3]~q ),
	.datab(!\act_counter[4]~q ),
	.datac(!\act_counter[5]~q ),
	.datad(!\act_counter[2]~q ),
	.datae(!\act_counter[1]~q ),
	.dataf(!\act_counter[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h0000000000000001;
defparam \Equal0~0 .shared_arith = "off";

arriaii_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \act_counter[1] (
	.clk(ctl_clk),
	.d(\Add0~5_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_6_0),
	.ena(vcc),
	.q(\act_counter[1]~q ),
	.prn(vcc));
defparam \act_counter[1] .is_wysiwyg = "true";
defparam \act_counter[1] .power_up = "low";

arriaii_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \act_counter[2] (
	.clk(ctl_clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_6_0),
	.ena(vcc),
	.q(\act_counter[2]~q ),
	.prn(vcc));
defparam \act_counter[2] .is_wysiwyg = "true";
defparam \act_counter[2] .power_up = "low";

dffeas \act_counter[3] (
	.clk(ctl_clk),
	.d(\Add0~13_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_6_0),
	.ena(vcc),
	.q(\act_counter[3]~q ),
	.prn(vcc));
defparam \act_counter[3] .is_wysiwyg = "true";
defparam \act_counter[3] .power_up = "low";

arriaii_lcell_comb \LessThan0~0 (
	.dataa(!act_to_rdwr_1),
	.datab(!\act_counter[3]~q ),
	.datac(!\act_counter[4]~q ),
	.datad(!\act_counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h4000400040004000;
defparam \LessThan0~0 .shared_arith = "off";

dffeas int_act_to_act_ready(
	.clk(ctl_clk),
	.d(\LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_6_0),
	.ena(vcc),
	.q(\int_act_to_act_ready~q ),
	.prn(vcc));
defparam int_act_to_act_ready.is_wysiwyg = "true";
defparam int_act_to_act_ready.power_up = "low";

arriaii_lcell_comb \rdwr_ready~0 (
	.dataa(!current_state1),
	.datab(!\LessThan0~0_combout ),
	.datac(!\act_counter[2]~q ),
	.datad(!\act_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdwr_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdwr_ready~0 .extended_lut = "off";
defparam \rdwr_ready~0 .lut_mask = 64'h4555455545554555;
defparam \rdwr_ready~0 .shared_arith = "off";

arriaii_lcell_comb \rdwr_ready~1 (
	.dataa(!act_to_rdwr_1),
	.datab(!close_6_0),
	.datac(!open_6_0),
	.datad(!\rdwr_ready~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdwr_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdwr_ready~1 .extended_lut = "off";
defparam \rdwr_ready~1 .lut_mask = 64'h0133013301330133;
defparam \rdwr_ready~1 .shared_arith = "off";

endmodule

module ddr3_int_alt_ddrx_bank_timer_info_7 (
	ctl_clk,
	do_read_r,
	do_write_r,
	current_state1,
	do_precharge_all_r,
	to_chip_r_0,
	always38,
	act_ready1,
	act_to_rdwr_1,
	always106,
	always145,
	ctl_reset_n,
	rdwr_ready1,
	always140,
	Equal0,
	close_7_0,
	open_7_0,
	general_counter,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	ctl_clk;
input 	do_read_r;
input 	do_write_r;
output 	current_state1;
input 	do_precharge_all_r;
input 	to_chip_r_0;
input 	always38;
output 	act_ready1;
input 	act_to_rdwr_1;
input 	always106;
input 	always145;
input 	ctl_reset_n;
output 	rdwr_ready1;
input 	always140;
input 	Equal0;
input 	close_7_0;
input 	open_7_0;
input 	general_counter;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \current_state~0_combout ;
wire \Add1~1_sumout ;
wire \general_counter~1_combout ;
wire \general_counter[0]~q ;
wire \Add1~10 ;
wire \Add1~13_sumout ;
wire \general_counter~3_combout ;
wire \general_counter[3]~q ;
wire \Add1~14 ;
wire \Add1~17_sumout ;
wire \general_counter~5_combout ;
wire \general_counter[4]~q ;
wire \Add1~18 ;
wire \Add1~21_sumout ;
wire \general_counter~4_combout ;
wire \general_counter[5]~q ;
wire \Equal1~0_combout ;
wire \Add1~2 ;
wire \Add1~5_sumout ;
wire \general_counter~2_combout ;
wire \general_counter[1]~q ;
wire \Add1~6 ;
wire \Add1~9_sumout ;
wire \general_counter~0_combout ;
wire \general_counter[2]~q ;
wire \doing_auto_precharge~0_combout ;
wire \doing_auto_precharge~1_combout ;
wire \doing_auto_precharge~q ;
wire \doing_precharge~0_combout ;
wire \doing_precharge~q ;
wire \int_rdwr_to_valid_ready~0_combout ;
wire \int_rdwr_to_valid_ready~1_combout ;
wire \doing_read~0_combout ;
wire \doing_read~q ;
wire \int_rdwr_to_valid_ready~2_combout ;
wire \int_rdwr_to_valid_ready~3_combout ;
wire \int_rdwr_to_valid_ready~q ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \act_counter[4]~q ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \act_counter[5]~q ;
wire \Add0~1_sumout ;
wire \act_counter[0]~q ;
wire \Equal0~0_combout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \act_counter[1]~q ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \act_counter[2]~q ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \act_counter[3]~q ;
wire \LessThan0~0_combout ;
wire \int_act_to_act_ready~q ;
wire \rdwr_ready~0_combout ;
wire \rdwr_ready~1_combout ;


dffeas current_state(
	.clk(ctl_clk),
	.d(\current_state~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_7_0),
	.ena(vcc),
	.q(current_state1),
	.prn(vcc));
defparam current_state.is_wysiwyg = "true";
defparam current_state.power_up = "low";

arriaii_lcell_comb act_ready(
	.dataa(!\int_rdwr_to_valid_ready~q ),
	.datab(!\int_act_to_act_ready~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(act_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam act_ready.extended_lut = "off";
defparam act_ready.lut_mask = 64'h4444444444444444;
defparam act_ready.shared_arith = "off";

dffeas rdwr_ready(
	.clk(ctl_clk),
	.d(\rdwr_ready~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rdwr_ready1),
	.prn(vcc));
defparam rdwr_ready.is_wysiwyg = "true";
defparam rdwr_ready.power_up = "low";

arriaii_lcell_comb \current_state~0 (
	.dataa(!always38),
	.datab(!always106),
	.datac(!current_state1),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\current_state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \current_state~0 .extended_lut = "off";
defparam \current_state~0 .lut_mask = 64'h0C080C080C080C08;
defparam \current_state~0 .shared_arith = "off";

arriaii_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Equal1~0_combout ),
	.datae(gnd),
	.dataf(!\general_counter[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(\Add1~2 ),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h0000FF000000FF00;
defparam \Add1~1 .shared_arith = "off";

arriaii_lcell_comb \general_counter~1 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!\Add1~1_sumout ),
	.datae(!general_counter),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~1 .extended_lut = "off";
defparam \general_counter~1 .lut_mask = 64'h00EC00EE00EC00EE;
defparam \general_counter~1 .shared_arith = "off";

dffeas \general_counter[0] (
	.clk(ctl_clk),
	.d(\general_counter~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[0]~q ),
	.prn(vcc));
defparam \general_counter[0] .is_wysiwyg = "true";
defparam \general_counter[0] .power_up = "low";

arriaii_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~9 .shared_arith = "off";

arriaii_lcell_comb \Add1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~13 .shared_arith = "off";

arriaii_lcell_comb \general_counter~3 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~13_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~3 .extended_lut = "off";
defparam \general_counter~3 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~3 .shared_arith = "off";

dffeas \general_counter[3] (
	.clk(ctl_clk),
	.d(\general_counter~3_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[3]~q ),
	.prn(vcc));
defparam \general_counter[3] .is_wysiwyg = "true";
defparam \general_counter[3] .power_up = "low";

arriaii_lcell_comb \Add1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~17 .shared_arith = "off";

arriaii_lcell_comb \general_counter~5 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~17_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~5 .extended_lut = "off";
defparam \general_counter~5 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~5 .shared_arith = "off";

dffeas \general_counter[4] (
	.clk(ctl_clk),
	.d(\general_counter~5_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[4]~q ),
	.prn(vcc));
defparam \general_counter[4] .is_wysiwyg = "true";
defparam \general_counter[4] .power_up = "low";

arriaii_lcell_comb \Add1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~21_sumout ),
	.cout(),
	.shareout());
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~21 .shared_arith = "off";

arriaii_lcell_comb \general_counter~4 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!general_counter),
	.datae(!\Add1~21_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~4 .extended_lut = "off";
defparam \general_counter~4 .lut_mask = 64'h0000ECEE0000ECEE;
defparam \general_counter~4 .shared_arith = "off";

dffeas \general_counter[5] (
	.clk(ctl_clk),
	.d(\general_counter~4_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[5]~q ),
	.prn(vcc));
defparam \general_counter[5] .is_wysiwyg = "true";
defparam \general_counter[5] .power_up = "low";

arriaii_lcell_comb \Equal1~0 (
	.dataa(!\general_counter[2]~q ),
	.datab(!\general_counter[0]~q ),
	.datac(!\general_counter[1]~q ),
	.datad(!\general_counter[3]~q ),
	.datae(!\general_counter[5]~q ),
	.dataf(!\general_counter[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'h0000000000000001;
defparam \Equal1~0 .shared_arith = "off";

arriaii_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\general_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~5 .shared_arith = "off";

arriaii_lcell_comb \general_counter~2 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!\Add1~5_sumout ),
	.datae(!general_counter),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~2 .extended_lut = "off";
defparam \general_counter~2 .lut_mask = 64'h00EC00EE00EC00EE;
defparam \general_counter~2 .shared_arith = "off";

dffeas \general_counter[1] (
	.clk(ctl_clk),
	.d(\general_counter~2_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[1]~q ),
	.prn(vcc));
defparam \general_counter[1] .is_wysiwyg = "true";
defparam \general_counter[1] .power_up = "low";

arriaii_lcell_comb \general_counter~0 (
	.dataa(!do_precharge_all_r),
	.datab(!to_chip_r_0),
	.datac(!Equal0),
	.datad(!\Add1~9_sumout ),
	.datae(!general_counter),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\general_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \general_counter~0 .extended_lut = "off";
defparam \general_counter~0 .lut_mask = 64'h13FF11FF13FF11FF;
defparam \general_counter~0 .shared_arith = "off";

dffeas \general_counter[2] (
	.clk(ctl_clk),
	.d(\general_counter~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\general_counter[2]~q ),
	.prn(vcc));
defparam \general_counter[2] .is_wysiwyg = "true";
defparam \general_counter[2] .power_up = "low";

arriaii_lcell_comb \doing_auto_precharge~0 (
	.dataa(!always38),
	.datab(!always106),
	.datac(!always140),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_auto_precharge~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_auto_precharge~0 .extended_lut = "off";
defparam \doing_auto_precharge~0 .lut_mask = 64'h0007000700070007;
defparam \doing_auto_precharge~0 .shared_arith = "off";

arriaii_lcell_comb \doing_auto_precharge~1 (
	.dataa(!always38),
	.datab(!always145),
	.datac(!always106),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_auto_precharge~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_auto_precharge~1 .extended_lut = "off";
defparam \doing_auto_precharge~1 .lut_mask = 64'h0F7F0F7F0F7F0F7F;
defparam \doing_auto_precharge~1 .shared_arith = "off";

dffeas doing_auto_precharge(
	.clk(ctl_clk),
	.d(\doing_auto_precharge~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\doing_auto_precharge~1_combout ),
	.q(\doing_auto_precharge~q ),
	.prn(vcc));
defparam doing_auto_precharge.is_wysiwyg = "true";
defparam doing_auto_precharge.power_up = "low";

arriaii_lcell_comb \doing_precharge~0 (
	.dataa(!always38),
	.datab(!always106),
	.datac(!always140),
	.datad(!Equal0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_precharge~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_precharge~0 .extended_lut = "off";
defparam \doing_precharge~0 .lut_mask = 64'h3370337033703370;
defparam \doing_precharge~0 .shared_arith = "off";

dffeas doing_precharge(
	.clk(ctl_clk),
	.d(\doing_precharge~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\doing_auto_precharge~1_combout ),
	.q(\doing_precharge~q ),
	.prn(vcc));
defparam doing_precharge.is_wysiwyg = "true";
defparam doing_precharge.power_up = "low";

arriaii_lcell_comb \int_rdwr_to_valid_ready~0 (
	.dataa(!\doing_read~q ),
	.datab(!\general_counter[0]~q ),
	.datac(!\general_counter[1]~q ),
	.datad(!\doing_auto_precharge~q ),
	.datae(!\general_counter[3]~q ),
	.dataf(!\doing_precharge~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_rdwr_to_valid_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_rdwr_to_valid_ready~0 .extended_lut = "off";
defparam \int_rdwr_to_valid_ready~0 .lut_mask = 64'hA8EA000000000000;
defparam \int_rdwr_to_valid_ready~0 .shared_arith = "off";

arriaii_lcell_comb \int_rdwr_to_valid_ready~1 (
	.dataa(!\general_counter[0]~q ),
	.datab(!\general_counter[1]~q ),
	.datac(!\doing_precharge~q ),
	.datad(!\general_counter[5]~q ),
	.datae(!\general_counter[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_rdwr_to_valid_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_rdwr_to_valid_ready~1 .extended_lut = "off";
defparam \int_rdwr_to_valid_ready~1 .lut_mask = 64'hFE000000FE000000;
defparam \int_rdwr_to_valid_ready~1 .shared_arith = "off";

arriaii_lcell_comb \doing_read~0 (
	.dataa(!do_read_r),
	.datab(!to_chip_r_0),
	.datac(!do_write_r),
	.datad(!Equal0),
	.datae(!\doing_read~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_read~0 .extended_lut = "off";
defparam \doing_read~0 .lut_mask = 64'h0010FFFC0010FFFC;
defparam \doing_read~0 .shared_arith = "off";

dffeas doing_read(
	.clk(ctl_clk),
	.d(\doing_read~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_read~q ),
	.prn(vcc));
defparam doing_read.is_wysiwyg = "true";
defparam doing_read.power_up = "low";

arriaii_lcell_comb \int_rdwr_to_valid_ready~2 (
	.dataa(!act_to_rdwr_1),
	.datab(!\doing_read~q ),
	.datac(!\general_counter[1]~q ),
	.datad(!\doing_auto_precharge~q ),
	.datae(!\general_counter[3]~q ),
	.dataf(!\doing_precharge~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_rdwr_to_valid_ready~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_rdwr_to_valid_ready~2 .extended_lut = "off";
defparam \int_rdwr_to_valid_ready~2 .lut_mask = 64'h54550040FFFF0000;
defparam \int_rdwr_to_valid_ready~2 .shared_arith = "off";

arriaii_lcell_comb \int_rdwr_to_valid_ready~3 (
	.dataa(!close_7_0),
	.datab(!\general_counter[2]~q ),
	.datac(!\int_rdwr_to_valid_ready~0_combout ),
	.datad(!\int_rdwr_to_valid_ready~1_combout ),
	.datae(!\int_rdwr_to_valid_ready~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_rdwr_to_valid_ready~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_rdwr_to_valid_ready~3 .extended_lut = "off";
defparam \int_rdwr_to_valid_ready~3 .lut_mask = 64'h5555551055555510;
defparam \int_rdwr_to_valid_ready~3 .shared_arith = "off";

dffeas int_rdwr_to_valid_ready(
	.clk(ctl_clk),
	.d(\int_rdwr_to_valid_ready~3_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\int_rdwr_to_valid_ready~q ),
	.prn(vcc));
defparam int_rdwr_to_valid_ready.is_wysiwyg = "true";
defparam int_rdwr_to_valid_ready.power_up = "low";

arriaii_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~13 .shared_arith = "off";

arriaii_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \act_counter[4] (
	.clk(ctl_clk),
	.d(\Add0~17_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_7_0),
	.ena(vcc),
	.q(\act_counter[4]~q ),
	.prn(vcc));
defparam \act_counter[4] .is_wysiwyg = "true";
defparam \act_counter[4] .power_up = "low";

arriaii_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \act_counter[5] (
	.clk(ctl_clk),
	.d(\Add0~21_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_7_0),
	.ena(vcc),
	.q(\act_counter[5]~q ),
	.prn(vcc));
defparam \act_counter[5] .is_wysiwyg = "true";
defparam \act_counter[5] .power_up = "low";

arriaii_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Equal0~0_combout ),
	.datae(gnd),
	.dataf(!\act_counter[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF000000FF00;
defparam \Add0~1 .shared_arith = "off";

dffeas \act_counter[0] (
	.clk(ctl_clk),
	.d(\Add0~1_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_7_0),
	.ena(vcc),
	.q(\act_counter[0]~q ),
	.prn(vcc));
defparam \act_counter[0] .is_wysiwyg = "true";
defparam \act_counter[0] .power_up = "low";

arriaii_lcell_comb \Equal0~0 (
	.dataa(!\act_counter[3]~q ),
	.datab(!\act_counter[4]~q ),
	.datac(!\act_counter[5]~q ),
	.datad(!\act_counter[2]~q ),
	.datae(!\act_counter[1]~q ),
	.dataf(!\act_counter[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h0000000000000001;
defparam \Equal0~0 .shared_arith = "off";

arriaii_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \act_counter[1] (
	.clk(ctl_clk),
	.d(\Add0~5_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_7_0),
	.ena(vcc),
	.q(\act_counter[1]~q ),
	.prn(vcc));
defparam \act_counter[1] .is_wysiwyg = "true";
defparam \act_counter[1] .power_up = "low";

arriaii_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \act_counter[2] (
	.clk(ctl_clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_7_0),
	.ena(vcc),
	.q(\act_counter[2]~q ),
	.prn(vcc));
defparam \act_counter[2] .is_wysiwyg = "true";
defparam \act_counter[2] .power_up = "low";

dffeas \act_counter[3] (
	.clk(ctl_clk),
	.d(\Add0~13_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_7_0),
	.ena(vcc),
	.q(\act_counter[3]~q ),
	.prn(vcc));
defparam \act_counter[3] .is_wysiwyg = "true";
defparam \act_counter[3] .power_up = "low";

arriaii_lcell_comb \LessThan0~0 (
	.dataa(!act_to_rdwr_1),
	.datab(!\act_counter[3]~q ),
	.datac(!\act_counter[4]~q ),
	.datad(!\act_counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h4000400040004000;
defparam \LessThan0~0 .shared_arith = "off";

dffeas int_act_to_act_ready(
	.clk(ctl_clk),
	.d(\LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(open_7_0),
	.ena(vcc),
	.q(\int_act_to_act_ready~q ),
	.prn(vcc));
defparam int_act_to_act_ready.is_wysiwyg = "true";
defparam int_act_to_act_ready.power_up = "low";

arriaii_lcell_comb \rdwr_ready~0 (
	.dataa(!current_state1),
	.datab(!\LessThan0~0_combout ),
	.datac(!\act_counter[2]~q ),
	.datad(!\act_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdwr_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdwr_ready~0 .extended_lut = "off";
defparam \rdwr_ready~0 .lut_mask = 64'h4555455545554555;
defparam \rdwr_ready~0 .shared_arith = "off";

arriaii_lcell_comb \rdwr_ready~1 (
	.dataa(!act_to_rdwr_1),
	.datab(!close_7_0),
	.datac(!open_7_0),
	.datad(!\rdwr_ready~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdwr_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdwr_ready~1 .extended_lut = "off";
defparam \rdwr_ready~1 .lut_mask = 64'h0133013301330133;
defparam \rdwr_ready~1 .shared_arith = "off";

endmodule

module ddr3_int_alt_ddrx_bypass (
	ctl_clk,
	out_cmd_info_valid_0,
	do_read,
	do_auto_precharge,
	do_write,
	out_cmd_info_valid_2,
	out_cmd_info_valid_3,
	out_cmd_info_valid_4,
	out_cmd_info_valid_1,
	pipe_10_0,
	pipe_12_0,
	pipe_11_0,
	act_cmd_monitor_per_chip0act_cmd_cnt0,
	act_trrd_ready_0,
	Mux0,
	pipe_12_2,
	pipe_12_3,
	pipe_12_1,
	pipe_10_2,
	pipe_10_3,
	pipe_10_1,
	pipe_11_2,
	pipe_11_3,
	pipe_11_1,
	pipe_12_4,
	pipe_11_4,
	pipe_10_4,
	Mux25,
	Mux5,
	fetch,
	do_precharge_all,
	out_cs_can_refresh_0,
	pipefull_0,
	out_cmd_can_activate_0,
	out_cmd_bank_is_open_0,
	to_chip,
	always38,
	to_bank_addr_r_2,
	current_bank_2,
	to_bank_addr_r_0,
	current_bank_0,
	to_bank_addr_r_1,
	current_bank_1,
	always381,
	out_cmd_can_write_0,
	out_cmd_can_read_0,
	out_cs_all_banks_closed_0,
	out_cs_can_precharge_all_0,
	do_activate,
	act_ready,
	act_ready1,
	act_ready2,
	act_ready3,
	act_ready4,
	power_saving_logic_per_chip0int_enter_power_saving_ready,
	act_ready5,
	act_ready6,
	act_ready7,
	Selector20,
	ctl_reset_n,
	pipefull_1,
	act_to_rdwr_1,
	int_cmd_info_valid,
	out_cmd_can_activate_2,
	out_cmd_bank_is_open_2,
	out_cmd_can_activate_3,
	out_cmd_bank_is_open_3,
	out_cmd_can_activate_4,
	out_cmd_bank_is_open_4,
	out_cmd_can_activate_1,
	out_cmd_bank_is_open_1,
	Mux10,
	Mux13,
	always106,
	always145,
	act_cmd_monitor_per_chip0act_cmd_cnt1,
	act_cmd_monitor_per_chip0act_cmd_cnt2,
	Mux1,
	can_al_activate_write,
	Mux12,
	rdwr_ready,
	rdwr_ready1,
	rdwr_ready2,
	rdwr_ready3,
	Mux9,
	can_al_activate_read,
	pipefull_4,
	cs_all_banks_closed_0,
	always140,
	pipefull_2,
	Mux16,
	Mux19,
	Mux3,
	Mux2,
	pipefull_3,
	Mux22,
	Mux4,
	always71,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	ctl_clk;
output 	out_cmd_info_valid_0;
input 	do_read;
input 	do_auto_precharge;
input 	do_write;
output 	out_cmd_info_valid_2;
output 	out_cmd_info_valid_3;
output 	out_cmd_info_valid_4;
output 	out_cmd_info_valid_1;
input 	pipe_10_0;
input 	pipe_12_0;
input 	pipe_11_0;
input 	act_cmd_monitor_per_chip0act_cmd_cnt0;
input 	act_trrd_ready_0;
input 	Mux0;
input 	pipe_12_2;
input 	pipe_12_3;
input 	pipe_12_1;
input 	pipe_10_2;
input 	pipe_10_3;
input 	pipe_10_1;
input 	pipe_11_2;
input 	pipe_11_3;
input 	pipe_11_1;
input 	pipe_12_4;
input 	pipe_11_4;
input 	pipe_10_4;
input 	Mux25;
input 	Mux5;
input 	fetch;
input 	do_precharge_all;
output 	out_cs_can_refresh_0;
input 	pipefull_0;
output 	out_cmd_can_activate_0;
output 	out_cmd_bank_is_open_0;
input 	[0:0] to_chip;
input 	always38;
input 	to_bank_addr_r_2;
input 	current_bank_2;
input 	to_bank_addr_r_0;
input 	current_bank_0;
input 	to_bank_addr_r_1;
input 	current_bank_1;
input 	always381;
output 	out_cmd_can_write_0;
output 	out_cmd_can_read_0;
output 	out_cs_all_banks_closed_0;
output 	out_cs_can_precharge_all_0;
input 	do_activate;
input 	act_ready;
input 	act_ready1;
input 	act_ready2;
input 	act_ready3;
input 	act_ready4;
input 	power_saving_logic_per_chip0int_enter_power_saving_ready;
input 	act_ready5;
input 	act_ready6;
input 	act_ready7;
input 	Selector20;
input 	ctl_reset_n;
input 	pipefull_1;
input 	act_to_rdwr_1;
input 	int_cmd_info_valid;
output 	out_cmd_can_activate_2;
output 	out_cmd_bank_is_open_2;
output 	out_cmd_can_activate_3;
output 	out_cmd_bank_is_open_3;
output 	out_cmd_can_activate_4;
output 	out_cmd_bank_is_open_4;
output 	out_cmd_can_activate_1;
output 	out_cmd_bank_is_open_1;
input 	Mux10;
input 	Mux13;
input 	always106;
output 	always145;
input 	act_cmd_monitor_per_chip0act_cmd_cnt1;
input 	act_cmd_monitor_per_chip0act_cmd_cnt2;
input 	Mux1;
input 	can_al_activate_write;
input 	Mux12;
input 	rdwr_ready;
input 	rdwr_ready1;
input 	rdwr_ready2;
input 	rdwr_ready3;
input 	Mux9;
input 	can_al_activate_read;
input 	pipefull_4;
input 	cs_all_banks_closed_0;
output 	always140;
input 	pipefull_2;
input 	Mux16;
input 	Mux19;
input 	Mux3;
input 	Mux2;
input 	pipefull_3;
input 	Mux22;
input 	Mux4;
output 	always71;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \out_cs_can_refresh~0_combout ;
wire \out_cs_can_refresh~1_combout ;
wire \do_auto_precharge_r1~q ;
wire \do_precharge_all_r1~q ;
wire \out_cs_can_refresh~2_combout ;
wire \out_cs_can_refresh~3_combout ;
wire \Equal1~0_combout ;
wire \cmd_close[0]~0_combout ;
wire \out_cmd_can_activate~0_combout ;
wire \always13~0_combout ;
wire \int_cmd_close_r1[1]~q ;
wire \cache_r1~q ;
wire \always5~0_combout ;
wire \int_cmd_close_r1[0]~q ;
wire \out_cmd_can_activate~1_combout ;
wire \out_cmd_can_activate~2_combout ;
wire \cmd_open[0]~0_combout ;
wire \out_cmd_bank_is_open~0_combout ;
wire \out_cmd_can_write~0_combout ;
wire \out_cmd_can_write~1_combout ;
wire \int_cmd_open_r1[1]~q ;
wire \int_cmd_open_r1[0]~q ;
wire \out_cmd_can_read~0_combout ;
wire \out_cmd_can_write~2_combout ;
wire \out_cmd_can_write~3_combout ;
wire \out_cmd_can_write~4_combout ;
wire \out_cmd_can_write~5_combout ;
wire \out_cmd_can_read~1_combout ;
wire \to_chip_r1[0]~q ;
wire \do_activate_r1~q ;
wire \out_cs_all_banks_closed~0_combout ;
wire \out_cs_all_banks_closed~1_combout ;
wire \do_write_r1~q ;
wire \do_read_r1~q ;
wire \out_cs_can_precharge_all~0_combout ;
wire \Equal2~0_combout ;
wire \Equal3~0_combout ;
wire \cmd_close[2]~1_combout ;
wire \always29~0_combout ;
wire \int_cmd_close_r1[3]~q ;
wire \always21~0_combout ;
wire \int_cmd_close_r1[2]~q ;
wire \out_cmd_can_activate~3_combout ;
wire \out_cmd_can_activate~4_combout ;
wire \out_cmd_bank_is_open~13_combout ;
wire \Equal4~0_combout ;
wire \cmd_close[3]~2_combout ;
wire \always37~0_combout ;
wire \int_cmd_close_r1[4]~q ;
wire \out_cmd_can_activate~5_combout ;
wire \out_cmd_can_activate~6_combout ;
wire \out_cmd_bank_is_open~9_combout ;
wire \always45~0_combout ;
wire \cmd_close[4]~3_combout ;
wire \always45~1_combout ;
wire \int_cmd_close_r1[5]~q ;
wire \out_cmd_can_activate~7_combout ;
wire \out_cmd_can_activate~8_combout ;
wire \out_cmd_bank_is_open~5_combout ;
wire \cmd_close[1]~4_combout ;
wire \out_cmd_can_activate~9_combout ;
wire \out_cmd_can_activate~10_combout ;
wire \out_cmd_bank_is_open~1_combout ;


dffeas \out_cmd_info_valid[0] (
	.clk(ctl_clk),
	.d(int_cmd_info_valid),
	.asdata(pipefull_0),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(fetch),
	.ena(vcc),
	.q(out_cmd_info_valid_0),
	.prn(vcc));
defparam \out_cmd_info_valid[0] .is_wysiwyg = "true";
defparam \out_cmd_info_valid[0] .power_up = "low";

dffeas \out_cmd_info_valid[2] (
	.clk(ctl_clk),
	.d(pipefull_1),
	.asdata(pipefull_2),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(fetch),
	.ena(vcc),
	.q(out_cmd_info_valid_2),
	.prn(vcc));
defparam \out_cmd_info_valid[2] .is_wysiwyg = "true";
defparam \out_cmd_info_valid[2] .power_up = "low";

dffeas \out_cmd_info_valid[3] (
	.clk(ctl_clk),
	.d(pipefull_2),
	.asdata(pipefull_3),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(fetch),
	.ena(vcc),
	.q(out_cmd_info_valid_3),
	.prn(vcc));
defparam \out_cmd_info_valid[3] .is_wysiwyg = "true";
defparam \out_cmd_info_valid[3] .power_up = "low";

dffeas \out_cmd_info_valid[4] (
	.clk(ctl_clk),
	.d(pipefull_3),
	.asdata(pipefull_4),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(fetch),
	.ena(vcc),
	.q(out_cmd_info_valid_4),
	.prn(vcc));
defparam \out_cmd_info_valid[4] .is_wysiwyg = "true";
defparam \out_cmd_info_valid[4] .power_up = "low";

dffeas \out_cmd_info_valid[1] (
	.clk(ctl_clk),
	.d(pipefull_0),
	.asdata(pipefull_1),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(fetch),
	.ena(vcc),
	.q(out_cmd_info_valid_1),
	.prn(vcc));
defparam \out_cmd_info_valid[1] .is_wysiwyg = "true";
defparam \out_cmd_info_valid[1] .power_up = "low";

dffeas \out_cs_can_refresh[0] (
	.clk(ctl_clk),
	.d(\out_cs_can_refresh~3_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_cs_can_refresh_0),
	.prn(vcc));
defparam \out_cs_can_refresh[0] .is_wysiwyg = "true";
defparam \out_cs_can_refresh[0] .power_up = "low";

dffeas \out_cmd_can_activate[0] (
	.clk(ctl_clk),
	.d(\out_cmd_can_activate~2_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_cmd_can_activate_0),
	.prn(vcc));
defparam \out_cmd_can_activate[0] .is_wysiwyg = "true";
defparam \out_cmd_can_activate[0] .power_up = "low";

dffeas \out_cmd_bank_is_open[0] (
	.clk(ctl_clk),
	.d(\out_cmd_bank_is_open~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_cmd_bank_is_open_0),
	.prn(vcc));
defparam \out_cmd_bank_is_open[0] .is_wysiwyg = "true";
defparam \out_cmd_bank_is_open[0] .power_up = "low";

dffeas \out_cmd_can_write[0] (
	.clk(ctl_clk),
	.d(\out_cmd_can_write~5_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_cmd_can_write_0),
	.prn(vcc));
defparam \out_cmd_can_write[0] .is_wysiwyg = "true";
defparam \out_cmd_can_write[0] .power_up = "low";

dffeas \out_cmd_can_read[0] (
	.clk(ctl_clk),
	.d(\out_cmd_can_read~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_cmd_can_read_0),
	.prn(vcc));
defparam \out_cmd_can_read[0] .is_wysiwyg = "true";
defparam \out_cmd_can_read[0] .power_up = "low";

dffeas \out_cs_all_banks_closed[0] (
	.clk(ctl_clk),
	.d(\out_cs_all_banks_closed~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_cs_all_banks_closed_0),
	.prn(vcc));
defparam \out_cs_all_banks_closed[0] .is_wysiwyg = "true";
defparam \out_cs_all_banks_closed[0] .power_up = "low";

dffeas \out_cs_can_precharge_all[0] (
	.clk(ctl_clk),
	.d(\out_cs_can_precharge_all~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_cs_can_precharge_all_0),
	.prn(vcc));
defparam \out_cs_can_precharge_all[0] .is_wysiwyg = "true";
defparam \out_cs_can_precharge_all[0] .power_up = "low";

dffeas \out_cmd_can_activate[2] (
	.clk(ctl_clk),
	.d(\out_cmd_can_activate~4_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_cmd_can_activate_2),
	.prn(vcc));
defparam \out_cmd_can_activate[2] .is_wysiwyg = "true";
defparam \out_cmd_can_activate[2] .power_up = "low";

dffeas \out_cmd_bank_is_open[2] (
	.clk(ctl_clk),
	.d(\out_cmd_bank_is_open~13_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_cmd_bank_is_open_2),
	.prn(vcc));
defparam \out_cmd_bank_is_open[2] .is_wysiwyg = "true";
defparam \out_cmd_bank_is_open[2] .power_up = "low";

dffeas \out_cmd_can_activate[3] (
	.clk(ctl_clk),
	.d(\out_cmd_can_activate~6_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_cmd_can_activate_3),
	.prn(vcc));
defparam \out_cmd_can_activate[3] .is_wysiwyg = "true";
defparam \out_cmd_can_activate[3] .power_up = "low";

dffeas \out_cmd_bank_is_open[3] (
	.clk(ctl_clk),
	.d(\out_cmd_bank_is_open~9_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_cmd_bank_is_open_3),
	.prn(vcc));
defparam \out_cmd_bank_is_open[3] .is_wysiwyg = "true";
defparam \out_cmd_bank_is_open[3] .power_up = "low";

dffeas \out_cmd_can_activate[4] (
	.clk(ctl_clk),
	.d(\out_cmd_can_activate~8_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_cmd_can_activate_4),
	.prn(vcc));
defparam \out_cmd_can_activate[4] .is_wysiwyg = "true";
defparam \out_cmd_can_activate[4] .power_up = "low";

dffeas \out_cmd_bank_is_open[4] (
	.clk(ctl_clk),
	.d(\out_cmd_bank_is_open~5_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_cmd_bank_is_open_4),
	.prn(vcc));
defparam \out_cmd_bank_is_open[4] .is_wysiwyg = "true";
defparam \out_cmd_bank_is_open[4] .power_up = "low";

dffeas \out_cmd_can_activate[1] (
	.clk(ctl_clk),
	.d(\out_cmd_can_activate~10_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_cmd_can_activate_1),
	.prn(vcc));
defparam \out_cmd_can_activate[1] .is_wysiwyg = "true";
defparam \out_cmd_can_activate[1] .power_up = "low";

dffeas \out_cmd_bank_is_open[1] (
	.clk(ctl_clk),
	.d(\out_cmd_bank_is_open~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_cmd_bank_is_open_1),
	.prn(vcc));
defparam \out_cmd_bank_is_open[1] .is_wysiwyg = "true";
defparam \out_cmd_bank_is_open[1] .power_up = "low";

arriaii_lcell_comb \always145~0 (
	.dataa(!to_chip[0]),
	.datab(!do_activate),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always145),
	.sumout(),
	.cout(),
	.shareout());
defparam \always145~0 .extended_lut = "off";
defparam \always145~0 .lut_mask = 64'h1111111111111111;
defparam \always145~0 .shared_arith = "off";

arriaii_lcell_comb \always140~0 (
	.dataa(!do_read),
	.datab(!to_chip[0]),
	.datac(!do_write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always140),
	.sumout(),
	.cout(),
	.shareout());
defparam \always140~0 .extended_lut = "off";
defparam \always140~0 .lut_mask = 64'h1313131313131313;
defparam \always140~0 .shared_arith = "off";

arriaii_lcell_comb \always71~0 (
	.dataa(!to_chip[0]),
	.datab(!do_write),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always71),
	.sumout(),
	.cout(),
	.shareout());
defparam \always71~0 .extended_lut = "off";
defparam \always71~0 .lut_mask = 64'h1111111111111111;
defparam \always71~0 .shared_arith = "off";

arriaii_lcell_comb \out_cs_can_refresh~0 (
	.dataa(!act_ready3),
	.datab(!act_ready4),
	.datac(!power_saving_logic_per_chip0int_enter_power_saving_ready),
	.datad(!act_ready5),
	.datae(!act_ready6),
	.dataf(!act_ready7),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cs_can_refresh~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cs_can_refresh~0 .extended_lut = "off";
defparam \out_cs_can_refresh~0 .lut_mask = 64'h0000000000000001;
defparam \out_cs_can_refresh~0 .shared_arith = "off";

arriaii_lcell_comb \out_cs_can_refresh~1 (
	.dataa(!\out_cs_all_banks_closed~0_combout ),
	.datab(!act_ready),
	.datac(!act_ready1),
	.datad(!act_ready2),
	.datae(!\out_cs_can_refresh~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cs_can_refresh~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cs_can_refresh~1 .extended_lut = "off";
defparam \out_cs_can_refresh~1 .lut_mask = 64'h0000000200000002;
defparam \out_cs_can_refresh~1 .shared_arith = "off";

dffeas do_auto_precharge_r1(
	.clk(ctl_clk),
	.d(do_auto_precharge),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\do_auto_precharge_r1~q ),
	.prn(vcc));
defparam do_auto_precharge_r1.is_wysiwyg = "true";
defparam do_auto_precharge_r1.power_up = "low";

dffeas do_precharge_all_r1(
	.clk(ctl_clk),
	.d(do_precharge_all),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\do_precharge_all_r1~q ),
	.prn(vcc));
defparam do_precharge_all_r1.is_wysiwyg = "true";
defparam do_precharge_all_r1.power_up = "low";

arriaii_lcell_comb \out_cs_can_refresh~2 (
	.dataa(!\to_chip_r1[0]~q ),
	.datab(!\do_auto_precharge_r1~q ),
	.datac(!\do_precharge_all_r1~q ),
	.datad(!Selector20),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cs_can_refresh~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cs_can_refresh~2 .extended_lut = "off";
defparam \out_cs_can_refresh~2 .lut_mask = 64'hEA00EA00EA00EA00;
defparam \out_cs_can_refresh~2 .shared_arith = "off";

arriaii_lcell_comb \out_cs_can_refresh~3 (
	.dataa(!do_precharge_all),
	.datab(!to_chip[0]),
	.datac(!do_auto_precharge),
	.datad(!\out_cs_can_refresh~1_combout ),
	.datae(!\out_cs_can_refresh~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cs_can_refresh~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cs_can_refresh~3 .extended_lut = "off";
defparam \out_cs_can_refresh~3 .lut_mask = 64'h000000EC000000EC;
defparam \out_cs_can_refresh~3 .shared_arith = "off";

arriaii_lcell_comb \Equal1~0 (
	.dataa(!to_bank_addr_r_2),
	.datab(!to_bank_addr_r_0),
	.datac(!to_bank_addr_r_1),
	.datad(!pipe_10_0),
	.datae(!pipe_12_0),
	.dataf(!pipe_11_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'h8020401008020401;
defparam \Equal1~0 .shared_arith = "off";

arriaii_lcell_comb \cmd_close[0]~0 (
	.dataa(!fetch),
	.datab(!always38),
	.datac(!always381),
	.datad(!always106),
	.datae(!\Equal1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cmd_close[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cmd_close[0]~0 .extended_lut = "off";
defparam \cmd_close[0]~0 .lut_mask = 64'hFD00EC00FD00EC00;
defparam \cmd_close[0]~0 .shared_arith = "off";

arriaii_lcell_comb \out_cmd_can_activate~0 (
	.dataa(!always145),
	.datab(!power_saving_logic_per_chip0int_enter_power_saving_ready),
	.datac(!act_cmd_monitor_per_chip0act_cmd_cnt1),
	.datad(!act_cmd_monitor_per_chip0act_cmd_cnt0),
	.datae(!act_trrd_ready_0),
	.dataf(!act_cmd_monitor_per_chip0act_cmd_cnt2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cmd_can_activate~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cmd_can_activate~0 .extended_lut = "off";
defparam \out_cmd_can_activate~0 .lut_mask = 64'h0000333200000000;
defparam \out_cmd_can_activate~0 .shared_arith = "off";

arriaii_lcell_comb \always13~0 (
	.dataa(!always38),
	.datab(!always106),
	.datac(!\Equal1~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always13~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always13~0 .extended_lut = "off";
defparam \always13~0 .lut_mask = 64'h3737373737373737;
defparam \always13~0 .shared_arith = "off";

dffeas \int_cmd_close_r1[1] (
	.clk(ctl_clk),
	.d(\always13~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\int_cmd_close_r1[1]~q ),
	.prn(vcc));
defparam \int_cmd_close_r1[1] .is_wysiwyg = "true";
defparam \int_cmd_close_r1[1] .power_up = "low";

dffeas cache_r1(
	.clk(ctl_clk),
	.d(fetch),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\cache_r1~q ),
	.prn(vcc));
defparam cache_r1.is_wysiwyg = "true";
defparam cache_r1.power_up = "low";

arriaii_lcell_comb \always5~0 (
	.dataa(!always38),
	.datab(!always381),
	.datac(!always106),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always5~0 .extended_lut = "off";
defparam \always5~0 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \always5~0 .shared_arith = "off";

dffeas \int_cmd_close_r1[0] (
	.clk(ctl_clk),
	.d(\always5~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\int_cmd_close_r1[0]~q ),
	.prn(vcc));
defparam \int_cmd_close_r1[0] .is_wysiwyg = "true";
defparam \int_cmd_close_r1[0] .power_up = "low";

arriaii_lcell_comb \out_cmd_can_activate~1 (
	.dataa(!fetch),
	.datab(!\out_cmd_can_activate~0_combout ),
	.datac(!\int_cmd_close_r1[1]~q ),
	.datad(!\cache_r1~q ),
	.datae(!\int_cmd_close_r1[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cmd_can_activate~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cmd_can_activate~1 .extended_lut = "off";
defparam \out_cmd_can_activate~1 .lut_mask = 64'h3230103032301030;
defparam \out_cmd_can_activate~1 .shared_arith = "off";

arriaii_lcell_comb \out_cmd_can_activate~2 (
	.dataa(!fetch),
	.datab(!Mux10),
	.datac(!Mux13),
	.datad(!\cmd_close[0]~0_combout ),
	.datae(!\out_cmd_can_activate~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cmd_can_activate~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cmd_can_activate~2 .extended_lut = "off";
defparam \out_cmd_can_activate~2 .lut_mask = 64'h0000002700000027;
defparam \out_cmd_can_activate~2 .shared_arith = "off";

arriaii_lcell_comb \cmd_open[0]~0 (
	.dataa(!fetch),
	.datab(!always381),
	.datac(!always145),
	.datad(!\Equal1~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cmd_open[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cmd_open[0]~0 .extended_lut = "off";
defparam \cmd_open[0]~0 .lut_mask = 64'h0207020702070207;
defparam \cmd_open[0]~0 .shared_arith = "off";

arriaii_lcell_comb \out_cmd_bank_is_open~0 (
	.dataa(!fetch),
	.datab(!\cmd_close[0]~0_combout ),
	.datac(!Mux0),
	.datad(!\cmd_open[0]~0_combout ),
	.datae(!Mux1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cmd_bank_is_open~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cmd_bank_is_open~0 .extended_lut = "off";
defparam \out_cmd_bank_is_open~0 .lut_mask = 64'h02FF13FF02FF13FF;
defparam \out_cmd_bank_is_open~0 .shared_arith = "off";

arriaii_lcell_comb \out_cmd_can_write~0 (
	.dataa(!pipe_12_0),
	.datab(!pipe_11_0),
	.datac(!rdwr_ready),
	.datad(!rdwr_ready1),
	.datae(!rdwr_ready2),
	.dataf(!rdwr_ready3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cmd_can_write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cmd_can_write~0 .extended_lut = "off";
defparam \out_cmd_can_write~0 .lut_mask = 64'h084C2A6E195D3B7F;
defparam \out_cmd_can_write~0 .shared_arith = "off";

arriaii_lcell_comb \out_cmd_can_write~1 (
	.dataa(!fetch),
	.datab(!pipe_10_0),
	.datac(!Mux12),
	.datad(!\out_cmd_can_write~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cmd_can_write~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cmd_can_write~1 .extended_lut = "off";
defparam \out_cmd_can_write~1 .lut_mask = 64'h0145014501450145;
defparam \out_cmd_can_write~1 .shared_arith = "off";

dffeas \int_cmd_open_r1[1] (
	.clk(ctl_clk),
	.d(GND_port),
	.asdata(\Equal1~0_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(always145),
	.ena(vcc),
	.q(\int_cmd_open_r1[1]~q ),
	.prn(vcc));
defparam \int_cmd_open_r1[1] .is_wysiwyg = "true";
defparam \int_cmd_open_r1[1] .power_up = "low";

dffeas \int_cmd_open_r1[0] (
	.clk(ctl_clk),
	.d(GND_port),
	.asdata(always381),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(always145),
	.ena(vcc),
	.q(\int_cmd_open_r1[0]~q ),
	.prn(vcc));
defparam \int_cmd_open_r1[0] .is_wysiwyg = "true";
defparam \int_cmd_open_r1[0] .power_up = "low";

arriaii_lcell_comb \out_cmd_can_read~0 (
	.dataa(!fetch),
	.datab(!\cache_r1~q ),
	.datac(!\int_cmd_open_r1[1]~q ),
	.datad(!\int_cmd_open_r1[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cmd_can_read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cmd_can_read~0 .extended_lut = "off";
defparam \out_cmd_can_read~0 .lut_mask = 64'h078F078F078F078F;
defparam \out_cmd_can_read~0 .shared_arith = "off";

arriaii_lcell_comb \out_cmd_can_write~2 (
	.dataa(!current_bank_2),
	.datab(!current_bank_1),
	.datac(!rdwr_ready),
	.datad(!rdwr_ready1),
	.datae(!rdwr_ready2),
	.dataf(!rdwr_ready3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cmd_can_write~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cmd_can_write~2 .extended_lut = "off";
defparam \out_cmd_can_write~2 .lut_mask = 64'h084C2A6E195D3B7F;
defparam \out_cmd_can_write~2 .shared_arith = "off";

arriaii_lcell_comb \out_cmd_can_write~3 (
	.dataa(!fetch),
	.datab(!current_bank_0),
	.datac(!Mux9),
	.datad(!\out_cmd_can_write~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cmd_can_write~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cmd_can_write~3 .extended_lut = "off";
defparam \out_cmd_can_write~3 .lut_mask = 64'h028A028A028A028A;
defparam \out_cmd_can_write~3 .shared_arith = "off";

arriaii_lcell_comb \out_cmd_can_write~4 (
	.dataa(!act_to_rdwr_1),
	.datab(!\cmd_open[0]~0_combout ),
	.datac(!\out_cmd_can_write~1_combout ),
	.datad(!\out_cmd_can_read~0_combout ),
	.datae(!\out_cmd_can_write~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cmd_can_write~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cmd_can_write~4 .extended_lut = "off";
defparam \out_cmd_can_write~4 .lut_mask = 64'hE0A00000E0A00000;
defparam \out_cmd_can_write~4 .shared_arith = "off";

arriaii_lcell_comb \out_cmd_can_write~5 (
	.dataa(!can_al_activate_write),
	.datab(!\out_cmd_can_write~4_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cmd_can_write~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cmd_can_write~5 .extended_lut = "off";
defparam \out_cmd_can_write~5 .lut_mask = 64'h4444444444444444;
defparam \out_cmd_can_write~5 .shared_arith = "off";

arriaii_lcell_comb \out_cmd_can_read~1 (
	.dataa(!\out_cmd_can_write~4_combout ),
	.datab(!can_al_activate_read),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cmd_can_read~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cmd_can_read~1 .extended_lut = "off";
defparam \out_cmd_can_read~1 .lut_mask = 64'h2222222222222222;
defparam \out_cmd_can_read~1 .shared_arith = "off";

dffeas \to_chip_r1[0] (
	.clk(ctl_clk),
	.d(to_chip[0]),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\to_chip_r1[0]~q ),
	.prn(vcc));
defparam \to_chip_r1[0] .is_wysiwyg = "true";
defparam \to_chip_r1[0] .power_up = "low";

dffeas do_activate_r1(
	.clk(ctl_clk),
	.d(do_activate),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\do_activate_r1~q ),
	.prn(vcc));
defparam do_activate_r1.is_wysiwyg = "true";
defparam do_activate_r1.power_up = "low";

arriaii_lcell_comb \out_cs_all_banks_closed~0 (
	.dataa(!to_chip[0]),
	.datab(!\do_activate_r1~q ),
	.datac(!\to_chip_r1[0]~q ),
	.datad(!do_activate),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cs_all_banks_closed~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cs_all_banks_closed~0 .extended_lut = "off";
defparam \out_cs_all_banks_closed~0 .lut_mask = 64'h0357035703570357;
defparam \out_cs_all_banks_closed~0 .shared_arith = "off";

arriaii_lcell_comb \out_cs_all_banks_closed~1 (
	.dataa(!\to_chip_r1[0]~q ),
	.datab(!\out_cs_all_banks_closed~0_combout ),
	.datac(!\do_precharge_all_r1~q ),
	.datad(!always106),
	.datae(!cs_all_banks_closed_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cs_all_banks_closed~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cs_all_banks_closed~1 .extended_lut = "off";
defparam \out_cs_all_banks_closed~1 .lut_mask = 64'h04CCCCCC04CCCCCC;
defparam \out_cs_all_banks_closed~1 .shared_arith = "off";

dffeas do_write_r1(
	.clk(ctl_clk),
	.d(do_write),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\do_write_r1~q ),
	.prn(vcc));
defparam do_write_r1.is_wysiwyg = "true";
defparam do_write_r1.power_up = "low";

dffeas do_read_r1(
	.clk(ctl_clk),
	.d(do_read),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\do_read_r1~q ),
	.prn(vcc));
defparam do_read_r1.is_wysiwyg = "true";
defparam do_read_r1.power_up = "low";

arriaii_lcell_comb \out_cs_can_precharge_all~0 (
	.dataa(!\to_chip_r1[0]~q ),
	.datab(!\out_cs_can_refresh~1_combout ),
	.datac(!always140),
	.datad(!\do_write_r1~q ),
	.datae(!\do_read_r1~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cs_can_precharge_all~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cs_can_precharge_all~0 .extended_lut = "off";
defparam \out_cs_can_precharge_all~0 .lut_mask = 64'h3020202030202020;
defparam \out_cs_can_precharge_all~0 .shared_arith = "off";

arriaii_lcell_comb \Equal2~0 (
	.dataa(!to_bank_addr_r_2),
	.datab(!to_bank_addr_r_0),
	.datac(!to_bank_addr_r_1),
	.datad(!pipe_12_1),
	.datae(!pipe_10_1),
	.dataf(!pipe_11_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~0 .extended_lut = "off";
defparam \Equal2~0 .lut_mask = 64'h8040201008040201;
defparam \Equal2~0 .shared_arith = "off";

arriaii_lcell_comb \Equal3~0 (
	.dataa(!to_bank_addr_r_2),
	.datab(!to_bank_addr_r_0),
	.datac(!to_bank_addr_r_1),
	.datad(!pipe_12_2),
	.datae(!pipe_10_2),
	.dataf(!pipe_11_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~0 .extended_lut = "off";
defparam \Equal3~0 .lut_mask = 64'h8040201008040201;
defparam \Equal3~0 .shared_arith = "off";

arriaii_lcell_comb \cmd_close[2]~1 (
	.dataa(!fetch),
	.datab(!always38),
	.datac(!always106),
	.datad(!\Equal2~0_combout ),
	.datae(!\Equal3~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cmd_close[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cmd_close[2]~1 .extended_lut = "off";
defparam \cmd_close[2]~1 .lut_mask = 64'h0F2F1F3F0F2F1F3F;
defparam \cmd_close[2]~1 .shared_arith = "off";

arriaii_lcell_comb \always29~0 (
	.dataa(!always38),
	.datab(!always106),
	.datac(!\Equal3~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always29~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always29~0 .extended_lut = "off";
defparam \always29~0 .lut_mask = 64'h3737373737373737;
defparam \always29~0 .shared_arith = "off";

dffeas \int_cmd_close_r1[3] (
	.clk(ctl_clk),
	.d(\always29~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\int_cmd_close_r1[3]~q ),
	.prn(vcc));
defparam \int_cmd_close_r1[3] .is_wysiwyg = "true";
defparam \int_cmd_close_r1[3] .power_up = "low";

arriaii_lcell_comb \always21~0 (
	.dataa(!always38),
	.datab(!always106),
	.datac(!\Equal2~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always21~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always21~0 .extended_lut = "off";
defparam \always21~0 .lut_mask = 64'h3737373737373737;
defparam \always21~0 .shared_arith = "off";

dffeas \int_cmd_close_r1[2] (
	.clk(ctl_clk),
	.d(\always21~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\int_cmd_close_r1[2]~q ),
	.prn(vcc));
defparam \int_cmd_close_r1[2] .is_wysiwyg = "true";
defparam \int_cmd_close_r1[2] .power_up = "low";

arriaii_lcell_comb \out_cmd_can_activate~3 (
	.dataa(!fetch),
	.datab(!\out_cmd_can_activate~0_combout ),
	.datac(!\cache_r1~q ),
	.datad(!\int_cmd_close_r1[3]~q ),
	.datae(!\int_cmd_close_r1[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cmd_can_activate~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cmd_can_activate~3 .extended_lut = "off";
defparam \out_cmd_can_activate~3 .lut_mask = 64'h3320130033201300;
defparam \out_cmd_can_activate~3 .shared_arith = "off";

arriaii_lcell_comb \out_cmd_can_activate~4 (
	.dataa(!fetch),
	.datab(!Mux16),
	.datac(!Mux19),
	.datad(!\cmd_close[2]~1_combout ),
	.datae(!\out_cmd_can_activate~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cmd_can_activate~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cmd_can_activate~4 .extended_lut = "off";
defparam \out_cmd_can_activate~4 .lut_mask = 64'h0000270000002700;
defparam \out_cmd_can_activate~4 .shared_arith = "off";

arriaii_lcell_comb \out_cmd_bank_is_open~13 (
	.dataa(!always145),
	.datab(!\Equal3~0_combout ),
	.datac(!Mux3),
	.datad(!\Equal2~0_combout ),
	.datae(!fetch),
	.dataf(!\cmd_close[2]~1_combout ),
	.datag(!Mux2),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cmd_bank_is_open~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cmd_bank_is_open~13 .extended_lut = "on";
defparam \out_cmd_bank_is_open~13 .lut_mask = 64'h0F5F1F1F00551111;
defparam \out_cmd_bank_is_open~13 .shared_arith = "off";

arriaii_lcell_comb \Equal4~0 (
	.dataa(!to_bank_addr_r_2),
	.datab(!to_bank_addr_r_0),
	.datac(!to_bank_addr_r_1),
	.datad(!pipe_12_3),
	.datae(!pipe_10_3),
	.dataf(!pipe_11_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~0 .extended_lut = "off";
defparam \Equal4~0 .lut_mask = 64'h8040201008040201;
defparam \Equal4~0 .shared_arith = "off";

arriaii_lcell_comb \cmd_close[3]~2 (
	.dataa(!fetch),
	.datab(!always38),
	.datac(!always106),
	.datad(!\Equal3~0_combout ),
	.datae(!\Equal4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cmd_close[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cmd_close[3]~2 .extended_lut = "off";
defparam \cmd_close[3]~2 .lut_mask = 64'h0F2F1F3F0F2F1F3F;
defparam \cmd_close[3]~2 .shared_arith = "off";

arriaii_lcell_comb \always37~0 (
	.dataa(!always38),
	.datab(!always106),
	.datac(!\Equal4~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always37~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always37~0 .extended_lut = "off";
defparam \always37~0 .lut_mask = 64'h3737373737373737;
defparam \always37~0 .shared_arith = "off";

dffeas \int_cmd_close_r1[4] (
	.clk(ctl_clk),
	.d(\always37~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\int_cmd_close_r1[4]~q ),
	.prn(vcc));
defparam \int_cmd_close_r1[4] .is_wysiwyg = "true";
defparam \int_cmd_close_r1[4] .power_up = "low";

arriaii_lcell_comb \out_cmd_can_activate~5 (
	.dataa(!fetch),
	.datab(!\out_cmd_can_activate~0_combout ),
	.datac(!\cache_r1~q ),
	.datad(!\int_cmd_close_r1[3]~q ),
	.datae(!\int_cmd_close_r1[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cmd_can_activate~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cmd_can_activate~5 .extended_lut = "off";
defparam \out_cmd_can_activate~5 .lut_mask = 64'h3313200033132000;
defparam \out_cmd_can_activate~5 .shared_arith = "off";

arriaii_lcell_comb \out_cmd_can_activate~6 (
	.dataa(!fetch),
	.datab(!Mux19),
	.datac(!Mux22),
	.datad(!\cmd_close[3]~2_combout ),
	.datae(!\out_cmd_can_activate~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cmd_can_activate~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cmd_can_activate~6 .extended_lut = "off";
defparam \out_cmd_can_activate~6 .lut_mask = 64'h0000270000002700;
defparam \out_cmd_can_activate~6 .shared_arith = "off";

arriaii_lcell_comb \out_cmd_bank_is_open~9 (
	.dataa(!always145),
	.datab(!\Equal4~0_combout ),
	.datac(!Mux4),
	.datad(!\Equal3~0_combout ),
	.datae(!fetch),
	.dataf(!\cmd_close[3]~2_combout ),
	.datag(!Mux3),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cmd_bank_is_open~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cmd_bank_is_open~9 .extended_lut = "on";
defparam \out_cmd_bank_is_open~9 .lut_mask = 64'h0F5F1F1F00551111;
defparam \out_cmd_bank_is_open~9 .shared_arith = "off";

arriaii_lcell_comb \always45~0 (
	.dataa(!to_bank_addr_r_2),
	.datab(!to_bank_addr_r_0),
	.datac(!to_bank_addr_r_1),
	.datad(!pipe_12_4),
	.datae(!pipe_11_4),
	.dataf(!pipe_10_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always45~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always45~0 .extended_lut = "off";
defparam \always45~0 .lut_mask = 64'h8040080420100201;
defparam \always45~0 .shared_arith = "off";

arriaii_lcell_comb \cmd_close[4]~3 (
	.dataa(!fetch),
	.datab(!always38),
	.datac(!always106),
	.datad(!\Equal4~0_combout ),
	.datae(!\always45~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cmd_close[4]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cmd_close[4]~3 .extended_lut = "off";
defparam \cmd_close[4]~3 .lut_mask = 64'h0F2F1F3F0F2F1F3F;
defparam \cmd_close[4]~3 .shared_arith = "off";

arriaii_lcell_comb \always45~1 (
	.dataa(!always38),
	.datab(!always106),
	.datac(!\always45~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always45~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always45~1 .extended_lut = "off";
defparam \always45~1 .lut_mask = 64'h3737373737373737;
defparam \always45~1 .shared_arith = "off";

dffeas \int_cmd_close_r1[5] (
	.clk(ctl_clk),
	.d(\always45~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\int_cmd_close_r1[5]~q ),
	.prn(vcc));
defparam \int_cmd_close_r1[5] .is_wysiwyg = "true";
defparam \int_cmd_close_r1[5] .power_up = "low";

arriaii_lcell_comb \out_cmd_can_activate~7 (
	.dataa(!fetch),
	.datab(!\out_cmd_can_activate~0_combout ),
	.datac(!\cache_r1~q ),
	.datad(!\cmd_close[4]~3_combout ),
	.datae(!\int_cmd_close_r1[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cmd_can_activate~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cmd_can_activate~7 .extended_lut = "off";
defparam \out_cmd_can_activate~7 .lut_mask = 64'h3300200033002000;
defparam \out_cmd_can_activate~7 .shared_arith = "off";

arriaii_lcell_comb \out_cmd_can_activate~8 (
	.dataa(!fetch),
	.datab(!\cache_r1~q ),
	.datac(!Mux22),
	.datad(!\int_cmd_close_r1[4]~q ),
	.datae(!Mux25),
	.dataf(!\out_cmd_can_activate~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cmd_can_activate~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cmd_can_activate~8 .extended_lut = "off";
defparam \out_cmd_can_activate~8 .lut_mask = 64'h000000000A025F57;
defparam \out_cmd_can_activate~8 .shared_arith = "off";

arriaii_lcell_comb \out_cmd_bank_is_open~5 (
	.dataa(!always145),
	.datab(!\always45~0_combout ),
	.datac(!Mux5),
	.datad(!\Equal4~0_combout ),
	.datae(!fetch),
	.dataf(!\cmd_close[4]~3_combout ),
	.datag(!Mux4),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cmd_bank_is_open~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cmd_bank_is_open~5 .extended_lut = "on";
defparam \out_cmd_bank_is_open~5 .lut_mask = 64'h0F5F1F1F00551111;
defparam \out_cmd_bank_is_open~5 .shared_arith = "off";

arriaii_lcell_comb \cmd_close[1]~4 (
	.dataa(!fetch),
	.datab(!always38),
	.datac(!always106),
	.datad(!\Equal1~0_combout ),
	.datae(!\Equal2~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cmd_close[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cmd_close[1]~4 .extended_lut = "off";
defparam \cmd_close[1]~4 .lut_mask = 64'h0F2F1F3F0F2F1F3F;
defparam \cmd_close[1]~4 .shared_arith = "off";

arriaii_lcell_comb \out_cmd_can_activate~9 (
	.dataa(!fetch),
	.datab(!\out_cmd_can_activate~0_combout ),
	.datac(!\int_cmd_close_r1[1]~q ),
	.datad(!\cache_r1~q ),
	.datae(!\int_cmd_close_r1[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cmd_can_activate~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cmd_can_activate~9 .extended_lut = "off";
defparam \out_cmd_can_activate~9 .lut_mask = 64'h3133200031332000;
defparam \out_cmd_can_activate~9 .shared_arith = "off";

arriaii_lcell_comb \out_cmd_can_activate~10 (
	.dataa(!fetch),
	.datab(!Mux13),
	.datac(!Mux16),
	.datad(!\cmd_close[1]~4_combout ),
	.datae(!\out_cmd_can_activate~9_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cmd_can_activate~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cmd_can_activate~10 .extended_lut = "off";
defparam \out_cmd_can_activate~10 .lut_mask = 64'h0000270000002700;
defparam \out_cmd_can_activate~10 .shared_arith = "off";

arriaii_lcell_comb \out_cmd_bank_is_open~1 (
	.dataa(!always145),
	.datab(!\Equal2~0_combout ),
	.datac(!Mux2),
	.datad(!\Equal1~0_combout ),
	.datae(!fetch),
	.dataf(!\cmd_close[1]~4_combout ),
	.datag(!Mux1),
	.cin(gnd),
	.sharein(gnd),
	.combout(\out_cmd_bank_is_open~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \out_cmd_bank_is_open~1 .extended_lut = "on";
defparam \out_cmd_bank_is_open~1 .lut_mask = 64'h0F5F1F1F00551111;
defparam \out_cmd_bank_is_open~1 .shared_arith = "off";

endmodule

module ddr3_int_alt_ddrx_cache (
	ctl_clk,
	fetch,
	int_cmd_info_valid,
	ctl_reset_n)/* synthesis synthesis_greybox=0 */;
input 	ctl_clk;
input 	fetch;
output 	int_cmd_info_valid;
input 	ctl_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fetch_r1~q ;
wire \int_cmd_info_valid[0]~1_combout ;
wire \int_current_info_valid_r1~q ;


arriaii_lcell_comb \int_cmd_info_valid~0 (
	.dataa(!\int_current_info_valid_r1~q ),
	.datab(!\fetch_r1~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(int_cmd_info_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_cmd_info_valid~0 .extended_lut = "off";
defparam \int_cmd_info_valid~0 .lut_mask = 64'h7777777777777777;
defparam \int_cmd_info_valid~0 .shared_arith = "off";

dffeas fetch_r1(
	.clk(ctl_clk),
	.d(fetch),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fetch_r1~q ),
	.prn(vcc));
defparam fetch_r1.is_wysiwyg = "true";
defparam fetch_r1.power_up = "low";

arriaii_lcell_comb \int_cmd_info_valid[0]~1 (
	.dataa(!fetch),
	.datab(!\int_current_info_valid_r1~q ),
	.datac(!\fetch_r1~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_cmd_info_valid[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_cmd_info_valid[0]~1 .extended_lut = "off";
defparam \int_cmd_info_valid[0]~1 .lut_mask = 64'h2A2A2A2A2A2A2A2A;
defparam \int_cmd_info_valid[0]~1 .shared_arith = "off";

dffeas int_current_info_valid_r1(
	.clk(ctl_clk),
	.d(\int_cmd_info_valid[0]~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\int_current_info_valid_r1~q ),
	.prn(vcc));
defparam int_current_info_valid_r1.is_wysiwyg = "true";
defparam int_current_info_valid_r1.power_up = "low";

endmodule

module ddr3_int_alt_ddrx_rank_monitor (
	ctl_clk,
	auto_refresh_logic_per_chip0int_refresh_req,
	do_read_r,
	do_write_r,
	act_cmd_monitor_per_chip0act_cmd_cnt0,
	act_trrd_ready_0,
	write_dqs_ready1,
	read_dqs_ready1,
	do_burst_chop_r,
	do_precharge_all_r,
	do_refresh_r,
	add_lat_on,
	to_chip_r_0,
	power_saving_logic_per_chip0int_enter_power_saving_ready,
	Selector20,
	act_to_rdwr_1,
	ctl_reset_n,
	always145,
	act_cmd_monitor_per_chip0act_cmd_cnt1,
	act_cmd_monitor_per_chip0act_cmd_cnt2,
	write_to_read_finish_twtr_0,
	always1,
	always71,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	ctl_clk;
output 	auto_refresh_logic_per_chip0int_refresh_req;
input 	do_read_r;
input 	do_write_r;
output 	act_cmd_monitor_per_chip0act_cmd_cnt0;
output 	act_trrd_ready_0;
output 	write_dqs_ready1;
output 	read_dqs_ready1;
input 	do_burst_chop_r;
input 	do_precharge_all_r;
input 	do_refresh_r;
input 	add_lat_on;
input 	to_chip_r_0;
output 	power_saving_logic_per_chip0int_enter_power_saving_ready;
output 	Selector20;
input 	act_to_rdwr_1;
input 	ctl_reset_n;
input 	always145;
output 	act_cmd_monitor_per_chip0act_cmd_cnt1;
output 	act_cmd_monitor_per_chip0act_cmd_cnt2;
output 	write_to_read_finish_twtr_0;
input 	always1;
input 	always71;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add6~1_sumout ;
wire \refresh_cnt~1_combout ;
wire \auto_refresh_logic_per_chip[0].refresh_cnt[0]~q ;
wire \Equal10~0_combout ;
wire \Add6~42 ;
wire \Add6~45_sumout ;
wire \auto_refresh_logic_per_chip[0].refresh_cnt[11]~q ;
wire \Add6~46 ;
wire \Add6~49_sumout ;
wire \auto_refresh_logic_per_chip[0].refresh_cnt[12]~q ;
wire \Equal10~1_combout ;
wire \Equal10~2_combout ;
wire \Add6~2 ;
wire \Add6~5_sumout ;
wire \refresh_cnt~0_combout ;
wire \auto_refresh_logic_per_chip[0].refresh_cnt[1]~q ;
wire \Add6~6 ;
wire \Add6~9_sumout ;
wire \auto_refresh_logic_per_chip[0].refresh_cnt[2]~q ;
wire \Add6~10 ;
wire \Add6~13_sumout ;
wire \auto_refresh_logic_per_chip[0].refresh_cnt[3]~q ;
wire \Add6~14 ;
wire \Add6~17_sumout ;
wire \auto_refresh_logic_per_chip[0].refresh_cnt[4]~q ;
wire \Add6~18 ;
wire \Add6~21_sumout ;
wire \auto_refresh_logic_per_chip[0].refresh_cnt[5]~q ;
wire \Add6~22 ;
wire \Add6~25_sumout ;
wire \auto_refresh_logic_per_chip[0].refresh_cnt[6]~q ;
wire \Add6~26 ;
wire \Add6~29_sumout ;
wire \auto_refresh_logic_per_chip[0].refresh_cnt[7]~q ;
wire \Add6~30 ;
wire \Add6~33_sumout ;
wire \auto_refresh_logic_per_chip[0].refresh_cnt[8]~q ;
wire \Add6~34 ;
wire \Add6~37_sumout ;
wire \auto_refresh_logic_per_chip[0].refresh_cnt[9]~q ;
wire \Add6~38 ;
wire \Add6~41_sumout ;
wire \auto_refresh_logic_per_chip[0].refresh_cnt[10]~q ;
wire \LessThan12~0_combout ;
wire \LessThan12~1_combout ;
wire \LessThan12~2_combout ;
wire \act_cmd_monitor_per_chip[0].act_cmd_cnt[0]~_wirecell_combout ;
wire \act_cmd_monitor_per_chip[0].act_tfaw_shift_reg[0]~q ;
wire \act_cmd_monitor_per_chip[0].act_tfaw_shift_reg[1]~q ;
wire \act_cmd_monitor_per_chip[0].act_tfaw_shift_reg[2]~q ;
wire \act_cmd_monitor_per_chip[0].act_tfaw_shift_reg[3]~q ;
wire \Add0~0_combout ;
wire \Mux0~0_combout ;
wire \act_cmd_monitor_per_chip[0].act_cmd_cnt[1]~1_combout ;
wire \Add2~6 ;
wire \Add2~9_sumout ;
wire \act_cmd_monitor_per_chip[0].act_trrd_cnt[2]~q ;
wire \Add2~10 ;
wire \Add2~13_sumout ;
wire \act_cmd_monitor_per_chip[0].act_trrd_cnt[3]~q ;
wire \Add2~14 ;
wire \Add2~17_sumout ;
wire \act_cmd_monitor_per_chip[0].act_trrd_cnt[4]~q ;
wire \Add2~18 ;
wire \Add2~21_sumout ;
wire \act_cmd_monitor_per_chip[0].act_trrd_cnt[5]~q ;
wire \Add2~1_sumout ;
wire \act_cmd_monitor_per_chip[0].act_trrd_cnt[0]~q ;
wire \Equal1~0_combout ;
wire \Add2~2 ;
wire \Add2~5_sumout ;
wire \act_cmd_monitor_per_chip[0].act_trrd_cnt[1]~q ;
wire \LessThan1~0_combout ;
wire \Selector4~0_combout ;
wire \rdwr_state.IDLE~q ;
wire \Selector1~0_combout ;
wire \rdwr_state.WR~q ;
wire \Add3~1_sumout ;
wire \rdwr_cnt[0]~q ;
wire \Add3~14 ;
wire \Add3~17_sumout ;
wire \rdwr_cnt[4]~q ;
wire \Add3~18 ;
wire \Add3~21_sumout ;
wire \rdwr_cnt[5]~q ;
wire \Add3~22 ;
wire \Add3~25_sumout ;
wire \rdwr_cnt[6]~q ;
wire \Equal2~0_combout ;
wire \Equal2~1_combout ;
wire \Add3~2 ;
wire \Add3~5_sumout ;
wire \rdwr_cnt[1]~q ;
wire \Add3~6 ;
wire \Add3~9_sumout ;
wire \rdwr_cnt[2]~q ;
wire \Add3~10 ;
wire \Add3~13_sumout ;
wire \rdwr_cnt[3]~q ;
wire \LessThan5~0_combout ;
wire \LessThan5~1_combout ;
wire \rdwr_state.RD~0_combout ;
wire \rdwr_state.RD~q ;
wire \doing_burst_chop~0_combout ;
wire \doing_burst_chop~q ;
wire \Selector4~1_combout ;
wire \Selector4~2_combout ;
wire \Selector3~0_combout ;
wire \Selector3~1_combout ;
wire \Add5~10 ;
wire \Add5~13_sumout ;
wire \int_enter_power_saving_ready~0_combout ;
wire \power_saving_logic_per_chip[0].power_saving_cnt[3]~q ;
wire \Add5~14 ;
wire \Add5~17_sumout ;
wire \power_saving_logic_per_chip[0].power_saving_cnt[4]~q ;
wire \Add5~18 ;
wire \Add5~21_sumout ;
wire \power_saving_logic_per_chip[0].power_saving_cnt[5]~q ;
wire \Add5~22 ;
wire \Add5~25_sumout ;
wire \power_saving_logic_per_chip[0].power_saving_cnt[6]~q ;
wire \Add5~26 ;
wire \Add5~29_sumout ;
wire \power_saving_logic_per_chip[0].power_saving_cnt[7]~q ;
wire \Add5~30 ;
wire \Add5~33_sumout ;
wire \power_saving_logic_per_chip[0].power_saving_cnt[8]~q ;
wire \Add5~34 ;
wire \Add5~37_sumout ;
wire \power_saving_logic_per_chip[0].power_saving_cnt[9]~q ;
wire \Equal4~0_combout ;
wire \Equal4~1_combout ;
wire \Add5~1_sumout ;
wire \power_saving_logic_per_chip[0].power_saving_cnt[0]~q ;
wire \Add5~2 ;
wire \Add5~5_sumout ;
wire \power_saving_logic_per_chip[0].power_saving_cnt[1]~q ;
wire \Add5~6 ;
wire \Add5~9_sumout ;
wire \power_saving_cnt~0_combout ;
wire \power_saving_logic_per_chip[0].power_saving_cnt[2]~q ;
wire \LessThan10~0_combout ;
wire \LessThan9~0_combout ;
wire \Selector20~1_combout ;
wire \power_saving_logic_per_chip[0].power_saving_state[30]~q ;
wire \LessThan9~1_combout ;
wire \Selector6~0_combout ;
wire \act_cmd_monitor_per_chip[0].act_cmd_cnt[1]~0_combout ;
wire \act_cmd_monitor_per_chip[0].act_cmd_cnt[2]~0_combout ;
wire \Add4~2 ;
wire \Add4~5_sumout ;
wire \twtr_cnt[0][1]~q ;
wire \Add4~6 ;
wire \Add4~9_sumout ;
wire \twtr_cnt[0][2]~q ;
wire \Add4~10 ;
wire \Add4~13_sumout ;
wire \twtr_cnt[0][3]~q ;
wire \Add4~14 ;
wire \Add4~17_sumout ;
wire \twtr_cnt[0][4]~q ;
wire \Equal3~0_combout ;
wire \Add4~1_sumout ;
wire \twtr_cnt[0][0]~q ;
wire \LessThan8~0_combout ;


dffeas \auto_refresh_logic_per_chip[0].int_refresh_req (
	.clk(ctl_clk),
	.d(\LessThan12~2_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(Selector20),
	.sload(gnd),
	.ena(vcc),
	.q(auto_refresh_logic_per_chip0int_refresh_req),
	.prn(vcc));
defparam \auto_refresh_logic_per_chip[0].int_refresh_req .is_wysiwyg = "true";
defparam \auto_refresh_logic_per_chip[0].int_refresh_req .power_up = "low";

dffeas \act_cmd_monitor_per_chip[0].act_cmd_cnt[0] (
	.clk(ctl_clk),
	.d(\act_cmd_monitor_per_chip[0].act_cmd_cnt[0]~_wirecell_combout ),
	.asdata(\Add0~0_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(always145),
	.ena(\act_cmd_monitor_per_chip[0].act_cmd_cnt[1]~1_combout ),
	.q(act_cmd_monitor_per_chip0act_cmd_cnt0),
	.prn(vcc));
defparam \act_cmd_monitor_per_chip[0].act_cmd_cnt[0] .is_wysiwyg = "true";
defparam \act_cmd_monitor_per_chip[0].act_cmd_cnt[0] .power_up = "low";

dffeas \act_trrd_ready[0] (
	.clk(ctl_clk),
	.d(\LessThan1~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(always145),
	.ena(vcc),
	.q(act_trrd_ready_0),
	.prn(vcc));
defparam \act_trrd_ready[0] .is_wysiwyg = "true";
defparam \act_trrd_ready[0] .power_up = "low";

dffeas write_dqs_ready(
	.clk(ctl_clk),
	.d(\Selector4~2_combout ),
	.asdata(act_to_rdwr_1),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(do_write_r),
	.ena(vcc),
	.q(write_dqs_ready1),
	.prn(vcc));
defparam write_dqs_ready.is_wysiwyg = "true";
defparam write_dqs_ready.power_up = "low";

dffeas read_dqs_ready(
	.clk(ctl_clk),
	.d(\Selector3~1_combout ),
	.asdata(add_lat_on),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(do_write_r),
	.ena(vcc),
	.q(read_dqs_ready1),
	.prn(vcc));
defparam read_dqs_ready.is_wysiwyg = "true";
defparam read_dqs_ready.power_up = "low";

dffeas \power_saving_logic_per_chip[0].int_enter_power_saving_ready (
	.clk(ctl_clk),
	.d(\Selector6~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(power_saving_logic_per_chip0int_enter_power_saving_ready),
	.prn(vcc));
defparam \power_saving_logic_per_chip[0].int_enter_power_saving_ready .is_wysiwyg = "true";
defparam \power_saving_logic_per_chip[0].int_enter_power_saving_ready .power_up = "low";

arriaii_lcell_comb \Selector20~0 (
	.dataa(!do_refresh_r),
	.datab(!to_chip_r_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector20),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector20~0 .extended_lut = "off";
defparam \Selector20~0 .lut_mask = 64'h1111111111111111;
defparam \Selector20~0 .shared_arith = "off";

dffeas \act_cmd_monitor_per_chip[0].act_cmd_cnt[1] (
	.clk(ctl_clk),
	.d(\act_cmd_monitor_per_chip[0].act_cmd_cnt[1]~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(act_cmd_monitor_per_chip0act_cmd_cnt1),
	.prn(vcc));
defparam \act_cmd_monitor_per_chip[0].act_cmd_cnt[1] .is_wysiwyg = "true";
defparam \act_cmd_monitor_per_chip[0].act_cmd_cnt[1] .power_up = "low";

dffeas \act_cmd_monitor_per_chip[0].act_cmd_cnt[2] (
	.clk(ctl_clk),
	.d(\act_cmd_monitor_per_chip[0].act_cmd_cnt[2]~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(act_cmd_monitor_per_chip0act_cmd_cnt2),
	.prn(vcc));
defparam \act_cmd_monitor_per_chip[0].act_cmd_cnt[2] .is_wysiwyg = "true";
defparam \act_cmd_monitor_per_chip[0].act_cmd_cnt[2] .power_up = "low";

dffeas \write_to_read_finish_twtr[0] (
	.clk(ctl_clk),
	.d(\LessThan8~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(write_to_read_finish_twtr_0),
	.prn(vcc));
defparam \write_to_read_finish_twtr[0] .is_wysiwyg = "true";
defparam \write_to_read_finish_twtr[0] .power_up = "low";

arriaii_lcell_comb \Add6~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Equal10~2_combout ),
	.datae(gnd),
	.dataf(!\auto_refresh_logic_per_chip[0].refresh_cnt[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~1_sumout ),
	.cout(\Add6~2 ),
	.shareout());
defparam \Add6~1 .extended_lut = "off";
defparam \Add6~1 .lut_mask = 64'h0000FF000000FF00;
defparam \Add6~1 .shared_arith = "off";

arriaii_lcell_comb \refresh_cnt~1 (
	.dataa(!Selector20),
	.datab(!\Add6~1_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\refresh_cnt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \refresh_cnt~1 .extended_lut = "off";
defparam \refresh_cnt~1 .lut_mask = 64'h7777777777777777;
defparam \refresh_cnt~1 .shared_arith = "off";

dffeas \auto_refresh_logic_per_chip[0].refresh_cnt[0] (
	.clk(ctl_clk),
	.d(\refresh_cnt~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_refresh_logic_per_chip[0].refresh_cnt[0]~q ),
	.prn(vcc));
defparam \auto_refresh_logic_per_chip[0].refresh_cnt[0] .is_wysiwyg = "true";
defparam \auto_refresh_logic_per_chip[0].refresh_cnt[0] .power_up = "low";

arriaii_lcell_comb \Equal10~0 (
	.dataa(!\auto_refresh_logic_per_chip[0].refresh_cnt[7]~q ),
	.datab(!\auto_refresh_logic_per_chip[0].refresh_cnt[4]~q ),
	.datac(!\auto_refresh_logic_per_chip[0].refresh_cnt[3]~q ),
	.datad(!\auto_refresh_logic_per_chip[0].refresh_cnt[6]~q ),
	.datae(!\auto_refresh_logic_per_chip[0].refresh_cnt[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal10~0 .extended_lut = "off";
defparam \Equal10~0 .lut_mask = 64'h0000000100000001;
defparam \Equal10~0 .shared_arith = "off";

arriaii_lcell_comb \Add6~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\auto_refresh_logic_per_chip[0].refresh_cnt[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~41_sumout ),
	.cout(\Add6~42 ),
	.shareout());
defparam \Add6~41 .extended_lut = "off";
defparam \Add6~41 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add6~41 .shared_arith = "off";

arriaii_lcell_comb \Add6~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\auto_refresh_logic_per_chip[0].refresh_cnt[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~45_sumout ),
	.cout(\Add6~46 ),
	.shareout());
defparam \Add6~45 .extended_lut = "off";
defparam \Add6~45 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add6~45 .shared_arith = "off";

dffeas \auto_refresh_logic_per_chip[0].refresh_cnt[11] (
	.clk(ctl_clk),
	.d(\Add6~45_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(Selector20),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_refresh_logic_per_chip[0].refresh_cnt[11]~q ),
	.prn(vcc));
defparam \auto_refresh_logic_per_chip[0].refresh_cnt[11] .is_wysiwyg = "true";
defparam \auto_refresh_logic_per_chip[0].refresh_cnt[11] .power_up = "low";

arriaii_lcell_comb \Add6~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\auto_refresh_logic_per_chip[0].refresh_cnt[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~49_sumout ),
	.cout(),
	.shareout());
defparam \Add6~49 .extended_lut = "off";
defparam \Add6~49 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add6~49 .shared_arith = "off";

dffeas \auto_refresh_logic_per_chip[0].refresh_cnt[12] (
	.clk(ctl_clk),
	.d(\Add6~49_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(Selector20),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_refresh_logic_per_chip[0].refresh_cnt[12]~q ),
	.prn(vcc));
defparam \auto_refresh_logic_per_chip[0].refresh_cnt[12] .is_wysiwyg = "true";
defparam \auto_refresh_logic_per_chip[0].refresh_cnt[12] .power_up = "low";

arriaii_lcell_comb \Equal10~1 (
	.dataa(!\auto_refresh_logic_per_chip[0].refresh_cnt[10]~q ),
	.datab(!\auto_refresh_logic_per_chip[0].refresh_cnt[8]~q ),
	.datac(!\auto_refresh_logic_per_chip[0].refresh_cnt[9]~q ),
	.datad(!\auto_refresh_logic_per_chip[0].refresh_cnt[11]~q ),
	.datae(!\auto_refresh_logic_per_chip[0].refresh_cnt[12]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal10~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal10~1 .extended_lut = "off";
defparam \Equal10~1 .lut_mask = 64'h0000000100000001;
defparam \Equal10~1 .shared_arith = "off";

arriaii_lcell_comb \Equal10~2 (
	.dataa(!\auto_refresh_logic_per_chip[0].refresh_cnt[1]~q ),
	.datab(!\auto_refresh_logic_per_chip[0].refresh_cnt[0]~q ),
	.datac(!\auto_refresh_logic_per_chip[0].refresh_cnt[2]~q ),
	.datad(!\Equal10~0_combout ),
	.datae(!\Equal10~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal10~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal10~2 .extended_lut = "off";
defparam \Equal10~2 .lut_mask = 64'h0000000100000001;
defparam \Equal10~2 .shared_arith = "off";

arriaii_lcell_comb \Add6~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\auto_refresh_logic_per_chip[0].refresh_cnt[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~5_sumout ),
	.cout(\Add6~6 ),
	.shareout());
defparam \Add6~5 .extended_lut = "off";
defparam \Add6~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add6~5 .shared_arith = "off";

arriaii_lcell_comb \refresh_cnt~0 (
	.dataa(!Selector20),
	.datab(!\Add6~5_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\refresh_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \refresh_cnt~0 .extended_lut = "off";
defparam \refresh_cnt~0 .lut_mask = 64'h7777777777777777;
defparam \refresh_cnt~0 .shared_arith = "off";

dffeas \auto_refresh_logic_per_chip[0].refresh_cnt[1] (
	.clk(ctl_clk),
	.d(\refresh_cnt~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_refresh_logic_per_chip[0].refresh_cnt[1]~q ),
	.prn(vcc));
defparam \auto_refresh_logic_per_chip[0].refresh_cnt[1] .is_wysiwyg = "true";
defparam \auto_refresh_logic_per_chip[0].refresh_cnt[1] .power_up = "low";

arriaii_lcell_comb \Add6~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\auto_refresh_logic_per_chip[0].refresh_cnt[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~9_sumout ),
	.cout(\Add6~10 ),
	.shareout());
defparam \Add6~9 .extended_lut = "off";
defparam \Add6~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add6~9 .shared_arith = "off";

dffeas \auto_refresh_logic_per_chip[0].refresh_cnt[2] (
	.clk(ctl_clk),
	.d(\Add6~9_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(Selector20),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_refresh_logic_per_chip[0].refresh_cnt[2]~q ),
	.prn(vcc));
defparam \auto_refresh_logic_per_chip[0].refresh_cnt[2] .is_wysiwyg = "true";
defparam \auto_refresh_logic_per_chip[0].refresh_cnt[2] .power_up = "low";

arriaii_lcell_comb \Add6~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\auto_refresh_logic_per_chip[0].refresh_cnt[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~13_sumout ),
	.cout(\Add6~14 ),
	.shareout());
defparam \Add6~13 .extended_lut = "off";
defparam \Add6~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add6~13 .shared_arith = "off";

dffeas \auto_refresh_logic_per_chip[0].refresh_cnt[3] (
	.clk(ctl_clk),
	.d(\Add6~13_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(Selector20),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_refresh_logic_per_chip[0].refresh_cnt[3]~q ),
	.prn(vcc));
defparam \auto_refresh_logic_per_chip[0].refresh_cnt[3] .is_wysiwyg = "true";
defparam \auto_refresh_logic_per_chip[0].refresh_cnt[3] .power_up = "low";

arriaii_lcell_comb \Add6~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\auto_refresh_logic_per_chip[0].refresh_cnt[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~17_sumout ),
	.cout(\Add6~18 ),
	.shareout());
defparam \Add6~17 .extended_lut = "off";
defparam \Add6~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add6~17 .shared_arith = "off";

dffeas \auto_refresh_logic_per_chip[0].refresh_cnt[4] (
	.clk(ctl_clk),
	.d(\Add6~17_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(Selector20),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_refresh_logic_per_chip[0].refresh_cnt[4]~q ),
	.prn(vcc));
defparam \auto_refresh_logic_per_chip[0].refresh_cnt[4] .is_wysiwyg = "true";
defparam \auto_refresh_logic_per_chip[0].refresh_cnt[4] .power_up = "low";

arriaii_lcell_comb \Add6~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\auto_refresh_logic_per_chip[0].refresh_cnt[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~21_sumout ),
	.cout(\Add6~22 ),
	.shareout());
defparam \Add6~21 .extended_lut = "off";
defparam \Add6~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add6~21 .shared_arith = "off";

dffeas \auto_refresh_logic_per_chip[0].refresh_cnt[5] (
	.clk(ctl_clk),
	.d(\Add6~21_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(Selector20),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_refresh_logic_per_chip[0].refresh_cnt[5]~q ),
	.prn(vcc));
defparam \auto_refresh_logic_per_chip[0].refresh_cnt[5] .is_wysiwyg = "true";
defparam \auto_refresh_logic_per_chip[0].refresh_cnt[5] .power_up = "low";

arriaii_lcell_comb \Add6~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\auto_refresh_logic_per_chip[0].refresh_cnt[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~25_sumout ),
	.cout(\Add6~26 ),
	.shareout());
defparam \Add6~25 .extended_lut = "off";
defparam \Add6~25 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add6~25 .shared_arith = "off";

dffeas \auto_refresh_logic_per_chip[0].refresh_cnt[6] (
	.clk(ctl_clk),
	.d(\Add6~25_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(Selector20),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_refresh_logic_per_chip[0].refresh_cnt[6]~q ),
	.prn(vcc));
defparam \auto_refresh_logic_per_chip[0].refresh_cnt[6] .is_wysiwyg = "true";
defparam \auto_refresh_logic_per_chip[0].refresh_cnt[6] .power_up = "low";

arriaii_lcell_comb \Add6~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\auto_refresh_logic_per_chip[0].refresh_cnt[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~29_sumout ),
	.cout(\Add6~30 ),
	.shareout());
defparam \Add6~29 .extended_lut = "off";
defparam \Add6~29 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add6~29 .shared_arith = "off";

dffeas \auto_refresh_logic_per_chip[0].refresh_cnt[7] (
	.clk(ctl_clk),
	.d(\Add6~29_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(Selector20),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_refresh_logic_per_chip[0].refresh_cnt[7]~q ),
	.prn(vcc));
defparam \auto_refresh_logic_per_chip[0].refresh_cnt[7] .is_wysiwyg = "true";
defparam \auto_refresh_logic_per_chip[0].refresh_cnt[7] .power_up = "low";

arriaii_lcell_comb \Add6~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\auto_refresh_logic_per_chip[0].refresh_cnt[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~33_sumout ),
	.cout(\Add6~34 ),
	.shareout());
defparam \Add6~33 .extended_lut = "off";
defparam \Add6~33 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add6~33 .shared_arith = "off";

dffeas \auto_refresh_logic_per_chip[0].refresh_cnt[8] (
	.clk(ctl_clk),
	.d(\Add6~33_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(Selector20),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_refresh_logic_per_chip[0].refresh_cnt[8]~q ),
	.prn(vcc));
defparam \auto_refresh_logic_per_chip[0].refresh_cnt[8] .is_wysiwyg = "true";
defparam \auto_refresh_logic_per_chip[0].refresh_cnt[8] .power_up = "low";

arriaii_lcell_comb \Add6~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\auto_refresh_logic_per_chip[0].refresh_cnt[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~37_sumout ),
	.cout(\Add6~38 ),
	.shareout());
defparam \Add6~37 .extended_lut = "off";
defparam \Add6~37 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add6~37 .shared_arith = "off";

dffeas \auto_refresh_logic_per_chip[0].refresh_cnt[9] (
	.clk(ctl_clk),
	.d(\Add6~37_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(Selector20),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_refresh_logic_per_chip[0].refresh_cnt[9]~q ),
	.prn(vcc));
defparam \auto_refresh_logic_per_chip[0].refresh_cnt[9] .is_wysiwyg = "true";
defparam \auto_refresh_logic_per_chip[0].refresh_cnt[9] .power_up = "low";

dffeas \auto_refresh_logic_per_chip[0].refresh_cnt[10] (
	.clk(ctl_clk),
	.d(\Add6~41_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(Selector20),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_refresh_logic_per_chip[0].refresh_cnt[10]~q ),
	.prn(vcc));
defparam \auto_refresh_logic_per_chip[0].refresh_cnt[10] .is_wysiwyg = "true";
defparam \auto_refresh_logic_per_chip[0].refresh_cnt[10] .power_up = "low";

arriaii_lcell_comb \LessThan12~0 (
	.dataa(!\auto_refresh_logic_per_chip[0].refresh_cnt[4]~q ),
	.datab(!\auto_refresh_logic_per_chip[0].refresh_cnt[1]~q ),
	.datac(!\auto_refresh_logic_per_chip[0].refresh_cnt[0]~q ),
	.datad(!\auto_refresh_logic_per_chip[0].refresh_cnt[3]~q ),
	.datae(!\auto_refresh_logic_per_chip[0].refresh_cnt[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan12~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan12~0 .extended_lut = "off";
defparam \LessThan12~0 .lut_mask = 64'h0155555501555555;
defparam \LessThan12~0 .shared_arith = "off";

arriaii_lcell_comb \LessThan12~1 (
	.dataa(!\auto_refresh_logic_per_chip[0].refresh_cnt[7]~q ),
	.datab(!\LessThan12~0_combout ),
	.datac(!\auto_refresh_logic_per_chip[0].refresh_cnt[6]~q ),
	.datad(!\auto_refresh_logic_per_chip[0].refresh_cnt[5]~q ),
	.datae(!\auto_refresh_logic_per_chip[0].refresh_cnt[8]~q ),
	.dataf(!\auto_refresh_logic_per_chip[0].refresh_cnt[9]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan12~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan12~1 .extended_lut = "off";
defparam \LessThan12~1 .lut_mask = 64'hEAAA000000000000;
defparam \LessThan12~1 .shared_arith = "off";

arriaii_lcell_comb \LessThan12~2 (
	.dataa(!\auto_refresh_logic_per_chip[0].refresh_cnt[10]~q ),
	.datab(!\LessThan12~1_combout ),
	.datac(!\auto_refresh_logic_per_chip[0].refresh_cnt[11]~q ),
	.datad(!act_to_rdwr_1),
	.datae(!\auto_refresh_logic_per_chip[0].refresh_cnt[12]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan12~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan12~2 .extended_lut = "off";
defparam \LessThan12~2 .lut_mask = 64'hFF4FFFFFFF4FFFFF;
defparam \LessThan12~2 .shared_arith = "off";

arriaii_lcell_comb \act_cmd_monitor_per_chip[0].act_cmd_cnt[0]~_wirecell (
	.dataa(!act_cmd_monitor_per_chip0act_cmd_cnt0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\act_cmd_monitor_per_chip[0].act_cmd_cnt[0]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \act_cmd_monitor_per_chip[0].act_cmd_cnt[0]~_wirecell .extended_lut = "off";
defparam \act_cmd_monitor_per_chip[0].act_cmd_cnt[0]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \act_cmd_monitor_per_chip[0].act_cmd_cnt[0]~_wirecell .shared_arith = "off";

dffeas \act_cmd_monitor_per_chip[0].act_tfaw_shift_reg[0] (
	.clk(ctl_clk),
	.d(always145),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\act_cmd_monitor_per_chip[0].act_tfaw_shift_reg[0]~q ),
	.prn(vcc));
defparam \act_cmd_monitor_per_chip[0].act_tfaw_shift_reg[0] .is_wysiwyg = "true";
defparam \act_cmd_monitor_per_chip[0].act_tfaw_shift_reg[0] .power_up = "low";

dffeas \act_cmd_monitor_per_chip[0].act_tfaw_shift_reg[1] (
	.clk(ctl_clk),
	.d(\act_cmd_monitor_per_chip[0].act_tfaw_shift_reg[0]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\act_cmd_monitor_per_chip[0].act_tfaw_shift_reg[1]~q ),
	.prn(vcc));
defparam \act_cmd_monitor_per_chip[0].act_tfaw_shift_reg[1] .is_wysiwyg = "true";
defparam \act_cmd_monitor_per_chip[0].act_tfaw_shift_reg[1] .power_up = "low";

dffeas \act_cmd_monitor_per_chip[0].act_tfaw_shift_reg[2] (
	.clk(ctl_clk),
	.d(\act_cmd_monitor_per_chip[0].act_tfaw_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\act_cmd_monitor_per_chip[0].act_tfaw_shift_reg[2]~q ),
	.prn(vcc));
defparam \act_cmd_monitor_per_chip[0].act_tfaw_shift_reg[2] .is_wysiwyg = "true";
defparam \act_cmd_monitor_per_chip[0].act_tfaw_shift_reg[2] .power_up = "low";

dffeas \act_cmd_monitor_per_chip[0].act_tfaw_shift_reg[3] (
	.clk(ctl_clk),
	.d(\act_cmd_monitor_per_chip[0].act_tfaw_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\act_cmd_monitor_per_chip[0].act_tfaw_shift_reg[3]~q ),
	.prn(vcc));
defparam \act_cmd_monitor_per_chip[0].act_tfaw_shift_reg[3] .is_wysiwyg = "true";
defparam \act_cmd_monitor_per_chip[0].act_tfaw_shift_reg[3] .power_up = "low";

arriaii_lcell_comb \Add0~0 (
	.dataa(!act_to_rdwr_1),
	.datab(!act_cmd_monitor_per_chip0act_cmd_cnt0),
	.datac(!\act_cmd_monitor_per_chip[0].act_tfaw_shift_reg[3]~q ),
	.datad(!\act_cmd_monitor_per_chip[0].act_tfaw_shift_reg[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'hC963C963C963C963;
defparam \Add0~0 .shared_arith = "off";

arriaii_lcell_comb \Mux0~0 (
	.dataa(!act_to_rdwr_1),
	.datab(!\act_cmd_monitor_per_chip[0].act_tfaw_shift_reg[3]~q ),
	.datac(!\act_cmd_monitor_per_chip[0].act_tfaw_shift_reg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~0 .extended_lut = "off";
defparam \Mux0~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \Mux0~0 .shared_arith = "off";

arriaii_lcell_comb \act_cmd_monitor_per_chip[0].act_cmd_cnt[1]~1 (
	.dataa(!always145),
	.datab(!\Mux0~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\act_cmd_monitor_per_chip[0].act_cmd_cnt[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \act_cmd_monitor_per_chip[0].act_cmd_cnt[1]~1 .extended_lut = "off";
defparam \act_cmd_monitor_per_chip[0].act_cmd_cnt[1]~1 .lut_mask = 64'h7777777777777777;
defparam \act_cmd_monitor_per_chip[0].act_cmd_cnt[1]~1 .shared_arith = "off";

arriaii_lcell_comb \Add2~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_cmd_monitor_per_chip[0].act_trrd_cnt[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~5_sumout ),
	.cout(\Add2~6 ),
	.shareout());
defparam \Add2~5 .extended_lut = "off";
defparam \Add2~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add2~5 .shared_arith = "off";

arriaii_lcell_comb \Add2~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_cmd_monitor_per_chip[0].act_trrd_cnt[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~9_sumout ),
	.cout(\Add2~10 ),
	.shareout());
defparam \Add2~9 .extended_lut = "off";
defparam \Add2~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add2~9 .shared_arith = "off";

dffeas \act_cmd_monitor_per_chip[0].act_trrd_cnt[2] (
	.clk(ctl_clk),
	.d(\Add2~9_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(always145),
	.ena(vcc),
	.q(\act_cmd_monitor_per_chip[0].act_trrd_cnt[2]~q ),
	.prn(vcc));
defparam \act_cmd_monitor_per_chip[0].act_trrd_cnt[2] .is_wysiwyg = "true";
defparam \act_cmd_monitor_per_chip[0].act_trrd_cnt[2] .power_up = "low";

arriaii_lcell_comb \Add2~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_cmd_monitor_per_chip[0].act_trrd_cnt[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~13_sumout ),
	.cout(\Add2~14 ),
	.shareout());
defparam \Add2~13 .extended_lut = "off";
defparam \Add2~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add2~13 .shared_arith = "off";

dffeas \act_cmd_monitor_per_chip[0].act_trrd_cnt[3] (
	.clk(ctl_clk),
	.d(\Add2~13_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(always145),
	.ena(vcc),
	.q(\act_cmd_monitor_per_chip[0].act_trrd_cnt[3]~q ),
	.prn(vcc));
defparam \act_cmd_monitor_per_chip[0].act_trrd_cnt[3] .is_wysiwyg = "true";
defparam \act_cmd_monitor_per_chip[0].act_trrd_cnt[3] .power_up = "low";

arriaii_lcell_comb \Add2~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_cmd_monitor_per_chip[0].act_trrd_cnt[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~17_sumout ),
	.cout(\Add2~18 ),
	.shareout());
defparam \Add2~17 .extended_lut = "off";
defparam \Add2~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add2~17 .shared_arith = "off";

dffeas \act_cmd_monitor_per_chip[0].act_trrd_cnt[4] (
	.clk(ctl_clk),
	.d(\Add2~17_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(always145),
	.ena(vcc),
	.q(\act_cmd_monitor_per_chip[0].act_trrd_cnt[4]~q ),
	.prn(vcc));
defparam \act_cmd_monitor_per_chip[0].act_trrd_cnt[4] .is_wysiwyg = "true";
defparam \act_cmd_monitor_per_chip[0].act_trrd_cnt[4] .power_up = "low";

arriaii_lcell_comb \Add2~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\act_cmd_monitor_per_chip[0].act_trrd_cnt[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~21_sumout ),
	.cout(),
	.shareout());
defparam \Add2~21 .extended_lut = "off";
defparam \Add2~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add2~21 .shared_arith = "off";

dffeas \act_cmd_monitor_per_chip[0].act_trrd_cnt[5] (
	.clk(ctl_clk),
	.d(\Add2~21_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(always145),
	.ena(vcc),
	.q(\act_cmd_monitor_per_chip[0].act_trrd_cnt[5]~q ),
	.prn(vcc));
defparam \act_cmd_monitor_per_chip[0].act_trrd_cnt[5] .is_wysiwyg = "true";
defparam \act_cmd_monitor_per_chip[0].act_trrd_cnt[5] .power_up = "low";

arriaii_lcell_comb \Add2~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Equal1~0_combout ),
	.datae(gnd),
	.dataf(!\act_cmd_monitor_per_chip[0].act_trrd_cnt[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~1_sumout ),
	.cout(\Add2~2 ),
	.shareout());
defparam \Add2~1 .extended_lut = "off";
defparam \Add2~1 .lut_mask = 64'h0000FF000000FF00;
defparam \Add2~1 .shared_arith = "off";

dffeas \act_cmd_monitor_per_chip[0].act_trrd_cnt[0] (
	.clk(ctl_clk),
	.d(\Add2~1_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(always145),
	.ena(vcc),
	.q(\act_cmd_monitor_per_chip[0].act_trrd_cnt[0]~q ),
	.prn(vcc));
defparam \act_cmd_monitor_per_chip[0].act_trrd_cnt[0] .is_wysiwyg = "true";
defparam \act_cmd_monitor_per_chip[0].act_trrd_cnt[0] .power_up = "low";

arriaii_lcell_comb \Equal1~0 (
	.dataa(!\act_cmd_monitor_per_chip[0].act_trrd_cnt[1]~q ),
	.datab(!\act_cmd_monitor_per_chip[0].act_trrd_cnt[2]~q ),
	.datac(!\act_cmd_monitor_per_chip[0].act_trrd_cnt[3]~q ),
	.datad(!\act_cmd_monitor_per_chip[0].act_trrd_cnt[4]~q ),
	.datae(!\act_cmd_monitor_per_chip[0].act_trrd_cnt[5]~q ),
	.dataf(!\act_cmd_monitor_per_chip[0].act_trrd_cnt[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'h0000000000000001;
defparam \Equal1~0 .shared_arith = "off";

dffeas \act_cmd_monitor_per_chip[0].act_trrd_cnt[1] (
	.clk(ctl_clk),
	.d(\Add2~5_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(always145),
	.ena(vcc),
	.q(\act_cmd_monitor_per_chip[0].act_trrd_cnt[1]~q ),
	.prn(vcc));
defparam \act_cmd_monitor_per_chip[0].act_trrd_cnt[1] .is_wysiwyg = "true";
defparam \act_cmd_monitor_per_chip[0].act_trrd_cnt[1] .power_up = "low";

arriaii_lcell_comb \LessThan1~0 (
	.dataa(!act_to_rdwr_1),
	.datab(!\act_cmd_monitor_per_chip[0].act_trrd_cnt[1]~q ),
	.datac(!\act_cmd_monitor_per_chip[0].act_trrd_cnt[2]~q ),
	.datad(!\act_cmd_monitor_per_chip[0].act_trrd_cnt[3]~q ),
	.datae(!\act_cmd_monitor_per_chip[0].act_trrd_cnt[4]~q ),
	.dataf(!\act_cmd_monitor_per_chip[0].act_trrd_cnt[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan1~0 .extended_lut = "off";
defparam \LessThan1~0 .lut_mask = 64'hBFFFFFFFFFFFFFFF;
defparam \LessThan1~0 .shared_arith = "off";

arriaii_lcell_comb \Selector4~0 (
	.dataa(!add_lat_on),
	.datab(!act_to_rdwr_1),
	.datac(!do_burst_chop_r),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~0 .extended_lut = "off";
defparam \Selector4~0 .lut_mask = 64'h5353535353535353;
defparam \Selector4~0 .shared_arith = "off";

dffeas \rdwr_state.IDLE (
	.clk(ctl_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.q(\rdwr_state.IDLE~q ),
	.prn(vcc));
defparam \rdwr_state.IDLE .is_wysiwyg = "true";
defparam \rdwr_state.IDLE .power_up = "low";

arriaii_lcell_comb \Selector1~0 (
	.dataa(!do_read_r),
	.datab(!do_write_r),
	.datac(!\rdwr_state.WR~q ),
	.datad(!\rdwr_state.IDLE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h333B333B333B333B;
defparam \Selector1~0 .shared_arith = "off";

dffeas \rdwr_state.WR (
	.clk(ctl_clk),
	.d(\Selector1~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdwr_state.WR~q ),
	.prn(vcc));
defparam \rdwr_state.WR .is_wysiwyg = "true";
defparam \rdwr_state.WR .power_up = "low";

arriaii_lcell_comb \Add3~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Equal2~1_combout ),
	.datae(gnd),
	.dataf(!\rdwr_cnt[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~1_sumout ),
	.cout(\Add3~2 ),
	.shareout());
defparam \Add3~1 .extended_lut = "off";
defparam \Add3~1 .lut_mask = 64'h0000FF000000FF00;
defparam \Add3~1 .shared_arith = "off";

dffeas \rdwr_cnt[0] (
	.clk(ctl_clk),
	.d(\Add3~1_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(always1),
	.ena(vcc),
	.q(\rdwr_cnt[0]~q ),
	.prn(vcc));
defparam \rdwr_cnt[0] .is_wysiwyg = "true";
defparam \rdwr_cnt[0] .power_up = "low";

arriaii_lcell_comb \Add3~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\rdwr_cnt[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~13_sumout ),
	.cout(\Add3~14 ),
	.shareout());
defparam \Add3~13 .extended_lut = "off";
defparam \Add3~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add3~13 .shared_arith = "off";

arriaii_lcell_comb \Add3~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\rdwr_cnt[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~17_sumout ),
	.cout(\Add3~18 ),
	.shareout());
defparam \Add3~17 .extended_lut = "off";
defparam \Add3~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add3~17 .shared_arith = "off";

dffeas \rdwr_cnt[4] (
	.clk(ctl_clk),
	.d(\Add3~17_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(always1),
	.ena(vcc),
	.q(\rdwr_cnt[4]~q ),
	.prn(vcc));
defparam \rdwr_cnt[4] .is_wysiwyg = "true";
defparam \rdwr_cnt[4] .power_up = "low";

arriaii_lcell_comb \Add3~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\rdwr_cnt[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~21_sumout ),
	.cout(\Add3~22 ),
	.shareout());
defparam \Add3~21 .extended_lut = "off";
defparam \Add3~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add3~21 .shared_arith = "off";

dffeas \rdwr_cnt[5] (
	.clk(ctl_clk),
	.d(\Add3~21_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(always1),
	.ena(vcc),
	.q(\rdwr_cnt[5]~q ),
	.prn(vcc));
defparam \rdwr_cnt[5] .is_wysiwyg = "true";
defparam \rdwr_cnt[5] .power_up = "low";

arriaii_lcell_comb \Add3~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\rdwr_cnt[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~25_sumout ),
	.cout(),
	.shareout());
defparam \Add3~25 .extended_lut = "off";
defparam \Add3~25 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add3~25 .shared_arith = "off";

dffeas \rdwr_cnt[6] (
	.clk(ctl_clk),
	.d(\Add3~25_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(always1),
	.ena(vcc),
	.q(\rdwr_cnt[6]~q ),
	.prn(vcc));
defparam \rdwr_cnt[6] .is_wysiwyg = "true";
defparam \rdwr_cnt[6] .power_up = "low";

arriaii_lcell_comb \Equal2~0 (
	.dataa(!\rdwr_cnt[3]~q ),
	.datab(!\rdwr_cnt[4]~q ),
	.datac(!\rdwr_cnt[5]~q ),
	.datad(!\rdwr_cnt[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~0 .extended_lut = "off";
defparam \Equal2~0 .lut_mask = 64'h0001000100010001;
defparam \Equal2~0 .shared_arith = "off";

arriaii_lcell_comb \Equal2~1 (
	.dataa(!\rdwr_cnt[2]~q ),
	.datab(!\rdwr_cnt[1]~q ),
	.datac(!\rdwr_cnt[0]~q ),
	.datad(!\Equal2~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~1 .extended_lut = "off";
defparam \Equal2~1 .lut_mask = 64'h0001000100010001;
defparam \Equal2~1 .shared_arith = "off";

arriaii_lcell_comb \Add3~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\rdwr_cnt[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~5_sumout ),
	.cout(\Add3~6 ),
	.shareout());
defparam \Add3~5 .extended_lut = "off";
defparam \Add3~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add3~5 .shared_arith = "off";

dffeas \rdwr_cnt[1] (
	.clk(ctl_clk),
	.d(\Add3~5_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(always1),
	.ena(vcc),
	.q(\rdwr_cnt[1]~q ),
	.prn(vcc));
defparam \rdwr_cnt[1] .is_wysiwyg = "true";
defparam \rdwr_cnt[1] .power_up = "low";

arriaii_lcell_comb \Add3~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\rdwr_cnt[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~9_sumout ),
	.cout(\Add3~10 ),
	.shareout());
defparam \Add3~9 .extended_lut = "off";
defparam \Add3~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add3~9 .shared_arith = "off";

dffeas \rdwr_cnt[2] (
	.clk(ctl_clk),
	.d(\Add3~9_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(always1),
	.ena(vcc),
	.q(\rdwr_cnt[2]~q ),
	.prn(vcc));
defparam \rdwr_cnt[2] .is_wysiwyg = "true";
defparam \rdwr_cnt[2] .power_up = "low";

dffeas \rdwr_cnt[3] (
	.clk(ctl_clk),
	.d(\Add3~13_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(always1),
	.ena(vcc),
	.q(\rdwr_cnt[3]~q ),
	.prn(vcc));
defparam \rdwr_cnt[3] .is_wysiwyg = "true";
defparam \rdwr_cnt[3] .power_up = "low";

arriaii_lcell_comb \LessThan5~0 (
	.dataa(!act_to_rdwr_1),
	.datab(!\rdwr_cnt[3]~q ),
	.datac(!\rdwr_cnt[4]~q ),
	.datad(!\rdwr_cnt[5]~q ),
	.datae(!\rdwr_cnt[6]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan5~0 .extended_lut = "off";
defparam \LessThan5~0 .lut_mask = 64'h4000000040000000;
defparam \LessThan5~0 .shared_arith = "off";

arriaii_lcell_comb \LessThan5~1 (
	.dataa(!\LessThan5~0_combout ),
	.datab(!\rdwr_cnt[2]~q ),
	.datac(!\rdwr_cnt[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan5~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan5~1 .extended_lut = "off";
defparam \LessThan5~1 .lut_mask = 64'h4040404040404040;
defparam \LessThan5~1 .shared_arith = "off";

arriaii_lcell_comb \rdwr_state.RD~0 (
	.dataa(!do_write_r),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdwr_state.RD~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdwr_state.RD~0 .extended_lut = "off";
defparam \rdwr_state.RD~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdwr_state.RD~0 .shared_arith = "off";

dffeas \rdwr_state.RD (
	.clk(ctl_clk),
	.d(\rdwr_state.RD~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.q(\rdwr_state.RD~q ),
	.prn(vcc));
defparam \rdwr_state.RD .is_wysiwyg = "true";
defparam \rdwr_state.RD .power_up = "low";

arriaii_lcell_comb \doing_burst_chop~0 (
	.dataa(!do_read_r),
	.datab(!do_write_r),
	.datac(!do_burst_chop_r),
	.datad(!\doing_burst_chop~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\doing_burst_chop~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \doing_burst_chop~0 .extended_lut = "off";
defparam \doing_burst_chop~0 .lut_mask = 64'h078F078F078F078F;
defparam \doing_burst_chop~0 .shared_arith = "off";

dffeas doing_burst_chop(
	.clk(ctl_clk),
	.d(\doing_burst_chop~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\doing_burst_chop~q ),
	.prn(vcc));
defparam doing_burst_chop.is_wysiwyg = "true";
defparam doing_burst_chop.power_up = "low";

arriaii_lcell_comb \Selector4~1 (
	.dataa(!\rdwr_cnt[2]~q ),
	.datab(!\rdwr_cnt[1]~q ),
	.datac(!\rdwr_state.RD~q ),
	.datad(!\rdwr_cnt[0]~q ),
	.datae(!\doing_burst_chop~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector4~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~1 .extended_lut = "off";
defparam \Selector4~1 .lut_mask = 64'h0E0A0A0A0E0A0A0A;
defparam \Selector4~1 .shared_arith = "off";

arriaii_lcell_comb \Selector4~2 (
	.dataa(!do_read_r),
	.datab(!\Selector4~0_combout ),
	.datac(!\rdwr_state.WR~q ),
	.datad(!\LessThan5~0_combout ),
	.datae(!\LessThan5~1_combout ),
	.dataf(!\Selector4~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector4~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~2 .extended_lut = "off";
defparam \Selector4~2 .lut_mask = 64'hBBBBB1B1BB11B111;
defparam \Selector4~2 .shared_arith = "off";

arriaii_lcell_comb \Selector3~0 (
	.dataa(!\rdwr_state.WR~q ),
	.datab(!\LessThan5~0_combout ),
	.datac(!\rdwr_cnt[2]~q ),
	.datad(!\rdwr_cnt[1]~q ),
	.datae(!\rdwr_cnt[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'h1111111011111110;
defparam \Selector3~0 .shared_arith = "off";

arriaii_lcell_comb \Selector3~1 (
	.dataa(!do_read_r),
	.datab(!act_to_rdwr_1),
	.datac(!\LessThan5~1_combout ),
	.datad(!\rdwr_state.RD~q ),
	.datae(!\Selector3~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~1 .extended_lut = "off";
defparam \Selector3~1 .lut_mask = 64'hBBB11111BBB11111;
defparam \Selector3~1 .shared_arith = "off";

arriaii_lcell_comb \Add5~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\power_saving_logic_per_chip[0].power_saving_cnt[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~9_sumout ),
	.cout(\Add5~10 ),
	.shareout());
defparam \Add5~9 .extended_lut = "off";
defparam \Add5~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add5~9 .shared_arith = "off";

arriaii_lcell_comb \Add5~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\power_saving_logic_per_chip[0].power_saving_cnt[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~13_sumout ),
	.cout(\Add5~14 ),
	.shareout());
defparam \Add5~13 .extended_lut = "off";
defparam \Add5~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add5~13 .shared_arith = "off";

arriaii_lcell_comb \int_enter_power_saving_ready~0 (
	.dataa(!do_precharge_all_r),
	.datab(!do_refresh_r),
	.datac(!to_chip_r_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\int_enter_power_saving_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \int_enter_power_saving_ready~0 .extended_lut = "off";
defparam \int_enter_power_saving_ready~0 .lut_mask = 64'h0707070707070707;
defparam \int_enter_power_saving_ready~0 .shared_arith = "off";

dffeas \power_saving_logic_per_chip[0].power_saving_cnt[3] (
	.clk(ctl_clk),
	.d(\Add5~13_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\int_enter_power_saving_ready~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\power_saving_logic_per_chip[0].power_saving_cnt[3]~q ),
	.prn(vcc));
defparam \power_saving_logic_per_chip[0].power_saving_cnt[3] .is_wysiwyg = "true";
defparam \power_saving_logic_per_chip[0].power_saving_cnt[3] .power_up = "low";

arriaii_lcell_comb \Add5~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\power_saving_logic_per_chip[0].power_saving_cnt[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~17_sumout ),
	.cout(\Add5~18 ),
	.shareout());
defparam \Add5~17 .extended_lut = "off";
defparam \Add5~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add5~17 .shared_arith = "off";

dffeas \power_saving_logic_per_chip[0].power_saving_cnt[4] (
	.clk(ctl_clk),
	.d(\Add5~17_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\int_enter_power_saving_ready~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\power_saving_logic_per_chip[0].power_saving_cnt[4]~q ),
	.prn(vcc));
defparam \power_saving_logic_per_chip[0].power_saving_cnt[4] .is_wysiwyg = "true";
defparam \power_saving_logic_per_chip[0].power_saving_cnt[4] .power_up = "low";

arriaii_lcell_comb \Add5~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\power_saving_logic_per_chip[0].power_saving_cnt[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~21_sumout ),
	.cout(\Add5~22 ),
	.shareout());
defparam \Add5~21 .extended_lut = "off";
defparam \Add5~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add5~21 .shared_arith = "off";

dffeas \power_saving_logic_per_chip[0].power_saving_cnt[5] (
	.clk(ctl_clk),
	.d(\Add5~21_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\int_enter_power_saving_ready~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\power_saving_logic_per_chip[0].power_saving_cnt[5]~q ),
	.prn(vcc));
defparam \power_saving_logic_per_chip[0].power_saving_cnt[5] .is_wysiwyg = "true";
defparam \power_saving_logic_per_chip[0].power_saving_cnt[5] .power_up = "low";

arriaii_lcell_comb \Add5~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\power_saving_logic_per_chip[0].power_saving_cnt[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~25_sumout ),
	.cout(\Add5~26 ),
	.shareout());
defparam \Add5~25 .extended_lut = "off";
defparam \Add5~25 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add5~25 .shared_arith = "off";

dffeas \power_saving_logic_per_chip[0].power_saving_cnt[6] (
	.clk(ctl_clk),
	.d(\Add5~25_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\int_enter_power_saving_ready~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\power_saving_logic_per_chip[0].power_saving_cnt[6]~q ),
	.prn(vcc));
defparam \power_saving_logic_per_chip[0].power_saving_cnt[6] .is_wysiwyg = "true";
defparam \power_saving_logic_per_chip[0].power_saving_cnt[6] .power_up = "low";

arriaii_lcell_comb \Add5~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\power_saving_logic_per_chip[0].power_saving_cnt[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~29_sumout ),
	.cout(\Add5~30 ),
	.shareout());
defparam \Add5~29 .extended_lut = "off";
defparam \Add5~29 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add5~29 .shared_arith = "off";

dffeas \power_saving_logic_per_chip[0].power_saving_cnt[7] (
	.clk(ctl_clk),
	.d(\Add5~29_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\int_enter_power_saving_ready~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\power_saving_logic_per_chip[0].power_saving_cnt[7]~q ),
	.prn(vcc));
defparam \power_saving_logic_per_chip[0].power_saving_cnt[7] .is_wysiwyg = "true";
defparam \power_saving_logic_per_chip[0].power_saving_cnt[7] .power_up = "low";

arriaii_lcell_comb \Add5~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\power_saving_logic_per_chip[0].power_saving_cnt[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~33_sumout ),
	.cout(\Add5~34 ),
	.shareout());
defparam \Add5~33 .extended_lut = "off";
defparam \Add5~33 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add5~33 .shared_arith = "off";

dffeas \power_saving_logic_per_chip[0].power_saving_cnt[8] (
	.clk(ctl_clk),
	.d(\Add5~33_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\int_enter_power_saving_ready~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\power_saving_logic_per_chip[0].power_saving_cnt[8]~q ),
	.prn(vcc));
defparam \power_saving_logic_per_chip[0].power_saving_cnt[8] .is_wysiwyg = "true";
defparam \power_saving_logic_per_chip[0].power_saving_cnt[8] .power_up = "low";

arriaii_lcell_comb \Add5~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\power_saving_logic_per_chip[0].power_saving_cnt[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~37_sumout ),
	.cout(),
	.shareout());
defparam \Add5~37 .extended_lut = "off";
defparam \Add5~37 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add5~37 .shared_arith = "off";

dffeas \power_saving_logic_per_chip[0].power_saving_cnt[9] (
	.clk(ctl_clk),
	.d(\Add5~37_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\int_enter_power_saving_ready~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\power_saving_logic_per_chip[0].power_saving_cnt[9]~q ),
	.prn(vcc));
defparam \power_saving_logic_per_chip[0].power_saving_cnt[9] .is_wysiwyg = "true";
defparam \power_saving_logic_per_chip[0].power_saving_cnt[9] .power_up = "low";

arriaii_lcell_comb \Equal4~0 (
	.dataa(!\power_saving_logic_per_chip[0].power_saving_cnt[4]~q ),
	.datab(!\power_saving_logic_per_chip[0].power_saving_cnt[2]~q ),
	.datac(!\power_saving_logic_per_chip[0].power_saving_cnt[3]~q ),
	.datad(!\power_saving_logic_per_chip[0].power_saving_cnt[5]~q ),
	.datae(!\power_saving_logic_per_chip[0].power_saving_cnt[9]~q ),
	.dataf(!\power_saving_logic_per_chip[0].power_saving_cnt[7]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~0 .extended_lut = "off";
defparam \Equal4~0 .lut_mask = 64'h0000000000000001;
defparam \Equal4~0 .shared_arith = "off";

arriaii_lcell_comb \Equal4~1 (
	.dataa(!\power_saving_logic_per_chip[0].power_saving_cnt[1]~q ),
	.datab(!\power_saving_logic_per_chip[0].power_saving_cnt[0]~q ),
	.datac(!\power_saving_logic_per_chip[0].power_saving_cnt[8]~q ),
	.datad(!\power_saving_logic_per_chip[0].power_saving_cnt[6]~q ),
	.datae(!\Equal4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~1 .extended_lut = "off";
defparam \Equal4~1 .lut_mask = 64'h0000000100000001;
defparam \Equal4~1 .shared_arith = "off";

arriaii_lcell_comb \Add5~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\power_saving_logic_per_chip[0].power_saving_cnt[0]~q ),
	.datae(gnd),
	.dataf(!\Equal4~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~1_sumout ),
	.cout(\Add5~2 ),
	.shareout());
defparam \Add5~1 .extended_lut = "off";
defparam \Add5~1 .lut_mask = 64'h000000FF000000FF;
defparam \Add5~1 .shared_arith = "off";

dffeas \power_saving_logic_per_chip[0].power_saving_cnt[0] (
	.clk(ctl_clk),
	.d(\Add5~1_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\int_enter_power_saving_ready~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\power_saving_logic_per_chip[0].power_saving_cnt[0]~q ),
	.prn(vcc));
defparam \power_saving_logic_per_chip[0].power_saving_cnt[0] .is_wysiwyg = "true";
defparam \power_saving_logic_per_chip[0].power_saving_cnt[0] .power_up = "low";

arriaii_lcell_comb \Add5~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\power_saving_logic_per_chip[0].power_saving_cnt[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add5~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~5_sumout ),
	.cout(\Add5~6 ),
	.shareout());
defparam \Add5~5 .extended_lut = "off";
defparam \Add5~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add5~5 .shared_arith = "off";

dffeas \power_saving_logic_per_chip[0].power_saving_cnt[1] (
	.clk(ctl_clk),
	.d(\Add5~5_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\int_enter_power_saving_ready~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\power_saving_logic_per_chip[0].power_saving_cnt[1]~q ),
	.prn(vcc));
defparam \power_saving_logic_per_chip[0].power_saving_cnt[1] .is_wysiwyg = "true";
defparam \power_saving_logic_per_chip[0].power_saving_cnt[1] .power_up = "low";

arriaii_lcell_comb \power_saving_cnt~0 (
	.dataa(!\int_enter_power_saving_ready~0_combout ),
	.datab(!\Add5~9_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\power_saving_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \power_saving_cnt~0 .extended_lut = "off";
defparam \power_saving_cnt~0 .lut_mask = 64'h7777777777777777;
defparam \power_saving_cnt~0 .shared_arith = "off";

dffeas \power_saving_logic_per_chip[0].power_saving_cnt[2] (
	.clk(ctl_clk),
	.d(\power_saving_cnt~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\power_saving_logic_per_chip[0].power_saving_cnt[2]~q ),
	.prn(vcc));
defparam \power_saving_logic_per_chip[0].power_saving_cnt[2] .is_wysiwyg = "true";
defparam \power_saving_logic_per_chip[0].power_saving_cnt[2] .power_up = "low";

arriaii_lcell_comb \LessThan10~0 (
	.dataa(!\power_saving_logic_per_chip[0].power_saving_cnt[4]~q ),
	.datab(!\power_saving_logic_per_chip[0].power_saving_cnt[2]~q ),
	.datac(!\power_saving_logic_per_chip[0].power_saving_cnt[3]~q ),
	.datad(!\power_saving_logic_per_chip[0].power_saving_cnt[1]~q ),
	.datae(!\power_saving_logic_per_chip[0].power_saving_cnt[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan10~0 .extended_lut = "off";
defparam \LessThan10~0 .lut_mask = 64'h1555555515555555;
defparam \LessThan10~0 .shared_arith = "off";

arriaii_lcell_comb \LessThan9~0 (
	.dataa(!act_to_rdwr_1),
	.datab(!\power_saving_logic_per_chip[0].power_saving_cnt[8]~q ),
	.datac(!\power_saving_logic_per_chip[0].power_saving_cnt[6]~q ),
	.datad(!\power_saving_logic_per_chip[0].power_saving_cnt[5]~q ),
	.datae(!\power_saving_logic_per_chip[0].power_saving_cnt[9]~q ),
	.dataf(!\power_saving_logic_per_chip[0].power_saving_cnt[7]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan9~0 .extended_lut = "off";
defparam \LessThan9~0 .lut_mask = 64'h4000000000000000;
defparam \LessThan9~0 .shared_arith = "off";

arriaii_lcell_comb \Selector20~1 (
	.dataa(!Selector20),
	.datab(!\power_saving_logic_per_chip[0].power_saving_state[30]~q ),
	.datac(!\LessThan10~0_combout ),
	.datad(!\LessThan9~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector20~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector20~1 .extended_lut = "off";
defparam \Selector20~1 .lut_mask = 64'h4474447444744474;
defparam \Selector20~1 .shared_arith = "off";

dffeas \power_saving_logic_per_chip[0].power_saving_state[30] (
	.clk(ctl_clk),
	.d(\Selector20~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\power_saving_logic_per_chip[0].power_saving_state[30]~q ),
	.prn(vcc));
defparam \power_saving_logic_per_chip[0].power_saving_state[30] .is_wysiwyg = "true";
defparam \power_saving_logic_per_chip[0].power_saving_state[30] .power_up = "low";

arriaii_lcell_comb \LessThan9~1 (
	.dataa(!\power_saving_logic_per_chip[0].power_saving_cnt[4]~q ),
	.datab(!\power_saving_logic_per_chip[0].power_saving_cnt[2]~q ),
	.datac(!\power_saving_logic_per_chip[0].power_saving_cnt[3]~q ),
	.datad(!\power_saving_logic_per_chip[0].power_saving_cnt[1]~q ),
	.datae(!\power_saving_logic_per_chip[0].power_saving_cnt[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan9~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan9~1 .extended_lut = "off";
defparam \LessThan9~1 .lut_mask = 64'h8080800080808000;
defparam \LessThan9~1 .shared_arith = "off";

arriaii_lcell_comb \Selector6~0 (
	.dataa(!\power_saving_logic_per_chip[0].power_saving_state[30]~q ),
	.datab(!\LessThan10~0_combout ),
	.datac(!\LessThan9~0_combout ),
	.datad(!\LessThan9~1_combout ),
	.datae(!\int_enter_power_saving_ready~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~0 .extended_lut = "off";
defparam \Selector6~0 .lut_mask = 64'hFBF15151FBF15151;
defparam \Selector6~0 .shared_arith = "off";

arriaii_lcell_comb \act_cmd_monitor_per_chip[0].act_cmd_cnt[1]~0 (
	.dataa(!always145),
	.datab(!act_cmd_monitor_per_chip0act_cmd_cnt1),
	.datac(!act_cmd_monitor_per_chip0act_cmd_cnt0),
	.datad(!\Mux0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\act_cmd_monitor_per_chip[0].act_cmd_cnt[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \act_cmd_monitor_per_chip[0].act_cmd_cnt[1]~0 .extended_lut = "off";
defparam \act_cmd_monitor_per_chip[0].act_cmd_cnt[1]~0 .lut_mask = 64'h3693369336933693;
defparam \act_cmd_monitor_per_chip[0].act_cmd_cnt[1]~0 .shared_arith = "off";

arriaii_lcell_comb \act_cmd_monitor_per_chip[0].act_cmd_cnt[2]~0 (
	.dataa(!always145),
	.datab(!act_cmd_monitor_per_chip0act_cmd_cnt1),
	.datac(!act_cmd_monitor_per_chip0act_cmd_cnt0),
	.datad(!act_cmd_monitor_per_chip0act_cmd_cnt2),
	.datae(!\Mux0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\act_cmd_monitor_per_chip[0].act_cmd_cnt[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \act_cmd_monitor_per_chip[0].act_cmd_cnt[2]~0 .extended_lut = "off";
defparam \act_cmd_monitor_per_chip[0].act_cmd_cnt[2]~0 .lut_mask = 64'h01FE807F01FE807F;
defparam \act_cmd_monitor_per_chip[0].act_cmd_cnt[2]~0 .shared_arith = "off";

arriaii_lcell_comb \Add4~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\Equal3~0_combout ),
	.datae(gnd),
	.dataf(!\twtr_cnt[0][0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~1_sumout ),
	.cout(\Add4~2 ),
	.shareout());
defparam \Add4~1 .extended_lut = "off";
defparam \Add4~1 .lut_mask = 64'h0000FF000000FF00;
defparam \Add4~1 .shared_arith = "off";

arriaii_lcell_comb \Add4~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\twtr_cnt[0][1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~5_sumout ),
	.cout(\Add4~6 ),
	.shareout());
defparam \Add4~5 .extended_lut = "off";
defparam \Add4~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add4~5 .shared_arith = "off";

dffeas \twtr_cnt[0][1] (
	.clk(ctl_clk),
	.d(\Add4~5_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(always71),
	.ena(vcc),
	.q(\twtr_cnt[0][1]~q ),
	.prn(vcc));
defparam \twtr_cnt[0][1] .is_wysiwyg = "true";
defparam \twtr_cnt[0][1] .power_up = "low";

arriaii_lcell_comb \Add4~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\twtr_cnt[0][2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~9_sumout ),
	.cout(\Add4~10 ),
	.shareout());
defparam \Add4~9 .extended_lut = "off";
defparam \Add4~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add4~9 .shared_arith = "off";

dffeas \twtr_cnt[0][2] (
	.clk(ctl_clk),
	.d(\Add4~9_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(always71),
	.ena(vcc),
	.q(\twtr_cnt[0][2]~q ),
	.prn(vcc));
defparam \twtr_cnt[0][2] .is_wysiwyg = "true";
defparam \twtr_cnt[0][2] .power_up = "low";

arriaii_lcell_comb \Add4~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\twtr_cnt[0][3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~13_sumout ),
	.cout(\Add4~14 ),
	.shareout());
defparam \Add4~13 .extended_lut = "off";
defparam \Add4~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add4~13 .shared_arith = "off";

dffeas \twtr_cnt[0][3] (
	.clk(ctl_clk),
	.d(\Add4~13_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(always71),
	.ena(vcc),
	.q(\twtr_cnt[0][3]~q ),
	.prn(vcc));
defparam \twtr_cnt[0][3] .is_wysiwyg = "true";
defparam \twtr_cnt[0][3] .power_up = "low";

arriaii_lcell_comb \Add4~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\twtr_cnt[0][4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~17_sumout ),
	.cout(),
	.shareout());
defparam \Add4~17 .extended_lut = "off";
defparam \Add4~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add4~17 .shared_arith = "off";

dffeas \twtr_cnt[0][4] (
	.clk(ctl_clk),
	.d(\Add4~17_sumout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(always71),
	.ena(vcc),
	.q(\twtr_cnt[0][4]~q ),
	.prn(vcc));
defparam \twtr_cnt[0][4] .is_wysiwyg = "true";
defparam \twtr_cnt[0][4] .power_up = "low";

arriaii_lcell_comb \Equal3~0 (
	.dataa(!\twtr_cnt[0][0]~q ),
	.datab(!\twtr_cnt[0][2]~q ),
	.datac(!\twtr_cnt[0][1]~q ),
	.datad(!\twtr_cnt[0][3]~q ),
	.datae(!\twtr_cnt[0][4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~0 .extended_lut = "off";
defparam \Equal3~0 .lut_mask = 64'h0000000100000001;
defparam \Equal3~0 .shared_arith = "off";

dffeas \twtr_cnt[0][0] (
	.clk(ctl_clk),
	.d(\Add4~1_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(always71),
	.ena(vcc),
	.q(\twtr_cnt[0][0]~q ),
	.prn(vcc));
defparam \twtr_cnt[0][0] .is_wysiwyg = "true";
defparam \twtr_cnt[0][0] .power_up = "low";

arriaii_lcell_comb \LessThan8~0 (
	.dataa(!act_to_rdwr_1),
	.datab(!\twtr_cnt[0][0]~q ),
	.datac(!\twtr_cnt[0][2]~q ),
	.datad(!\twtr_cnt[0][1]~q ),
	.datae(!\twtr_cnt[0][3]~q ),
	.dataf(!\twtr_cnt[0][4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan8~0 .extended_lut = "off";
defparam \LessThan8~0 .lut_mask = 64'hAAABFFFFFFFFFFFF;
defparam \LessThan8~0 .shared_arith = "off";

endmodule

module ddr3_int_alt_ddrx_timing_param (
	clk_0,
	add_lat_on1,
	act_to_rdwr_1,
	reset_reg_12,
	more_than_3_wr_to_pch1)/* synthesis synthesis_greybox=0 */;
input 	clk_0;
output 	add_lat_on1;
output 	act_to_rdwr_1;
input 	reset_reg_12;
output 	more_than_3_wr_to_pch1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_lat_on~0_combout ;


dffeas add_lat_on(
	.clk(clk_0),
	.d(\add_lat_on~0_combout ),
	.asdata(vcc),
	.clrn(reset_reg_12),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(add_lat_on1),
	.prn(vcc));
defparam add_lat_on.is_wysiwyg = "true";
defparam add_lat_on.power_up = "low";

dffeas \act_to_rdwr[1] (
	.clk(clk_0),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset_reg_12),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(act_to_rdwr_1),
	.prn(vcc));
defparam \act_to_rdwr[1] .is_wysiwyg = "true";
defparam \act_to_rdwr[1] .power_up = "low";

dffeas more_than_3_wr_to_pch(
	.clk(clk_0),
	.d(act_to_rdwr_1),
	.asdata(vcc),
	.clrn(reset_reg_12),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(more_than_3_wr_to_pch1),
	.prn(vcc));
defparam more_than_3_wr_to_pch.is_wysiwyg = "true";
defparam more_than_3_wr_to_pch.power_up = "low";

arriaii_lcell_comb \add_lat_on~0 (
	.dataa(!act_to_rdwr_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\add_lat_on~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \add_lat_on~0 .extended_lut = "off";
defparam \add_lat_on~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \add_lat_on~0 .shared_arith = "off";

endmodule

module ddr3_int_alt_ddrx_clock_and_reset (
	clk_0,
	reset_phy_clk_1x_n,
	reset_reg_4,
	reset_reg_5,
	reset_reg_7,
	reset_reg_3,
	reset_reg_14,
	reset_reg_16,
	reset_reg_11,
	reset_reg_9,
	reset_reg_12,
	reset_reg_8,
	reset_reg_10,
	reset_reg_15)/* synthesis synthesis_greybox=0 */;
input 	clk_0;
input 	reset_phy_clk_1x_n;
output 	reset_reg_4;
output 	reset_reg_5;
output 	reset_reg_7;
output 	reset_reg_3;
output 	reset_reg_14;
output 	reset_reg_16;
output 	reset_reg_11;
output 	reset_reg_9;
output 	reset_reg_12;
output 	reset_reg_8;
output 	reset_reg_10;
output 	reset_reg_15;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_alt_ddrx_reset_sync_1 reset_sync_inst(
	.clk(clk_0),
	.reset_n(reset_phy_clk_1x_n),
	.reset_reg_4(reset_reg_4),
	.reset_reg_5(reset_reg_5),
	.reset_reg_7(reset_reg_7),
	.reset_reg_3(reset_reg_3),
	.reset_reg_14(reset_reg_14),
	.reset_reg_16(reset_reg_16),
	.reset_reg_11(reset_reg_11),
	.reset_reg_9(reset_reg_9),
	.reset_reg_12(reset_reg_12),
	.reset_reg_8(reset_reg_8),
	.reset_reg_10(reset_reg_10),
	.reset_reg_15(reset_reg_15));

endmodule

module ddr3_int_alt_ddrx_reset_sync_1 (
	clk,
	reset_n,
	reset_reg_4,
	reset_reg_5,
	reset_reg_7,
	reset_reg_3,
	reset_reg_14,
	reset_reg_16,
	reset_reg_11,
	reset_reg_9,
	reset_reg_12,
	reset_reg_8,
	reset_reg_10,
	reset_reg_15)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	reset_n;
output 	reset_reg_4;
output 	reset_reg_5;
output 	reset_reg_7;
output 	reset_reg_3;
output 	reset_reg_14;
output 	reset_reg_16;
output 	reset_reg_11;
output 	reset_reg_9;
output 	reset_reg_12;
output 	reset_reg_8;
output 	reset_reg_10;
output 	reset_reg_15;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \reset_reg[0]~q ;
wire \reset_reg[1]~q ;
wire \reset_reg[2]~q ;


dffeas \reset_reg[4] (
	.clk(clk),
	.d(\reset_reg[2]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(reset_reg_4),
	.prn(vcc));
defparam \reset_reg[4] .is_wysiwyg = "true";
defparam \reset_reg[4] .power_up = "low";

dffeas \reset_reg[5] (
	.clk(clk),
	.d(\reset_reg[2]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(reset_reg_5),
	.prn(vcc));
defparam \reset_reg[5] .is_wysiwyg = "true";
defparam \reset_reg[5] .power_up = "low";

dffeas \reset_reg[7] (
	.clk(clk),
	.d(\reset_reg[2]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(reset_reg_7),
	.prn(vcc));
defparam \reset_reg[7] .is_wysiwyg = "true";
defparam \reset_reg[7] .power_up = "low";

dffeas \reset_reg[3] (
	.clk(clk),
	.d(\reset_reg[2]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(reset_reg_3),
	.prn(vcc));
defparam \reset_reg[3] .is_wysiwyg = "true";
defparam \reset_reg[3] .power_up = "low";

dffeas \reset_reg[14] (
	.clk(clk),
	.d(\reset_reg[2]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(reset_reg_14),
	.prn(vcc));
defparam \reset_reg[14] .is_wysiwyg = "true";
defparam \reset_reg[14] .power_up = "low";

dffeas \reset_reg[16] (
	.clk(clk),
	.d(\reset_reg[2]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(reset_reg_16),
	.prn(vcc));
defparam \reset_reg[16] .is_wysiwyg = "true";
defparam \reset_reg[16] .power_up = "low";

dffeas \reset_reg[11] (
	.clk(clk),
	.d(\reset_reg[2]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(reset_reg_11),
	.prn(vcc));
defparam \reset_reg[11] .is_wysiwyg = "true";
defparam \reset_reg[11] .power_up = "low";

dffeas \reset_reg[9] (
	.clk(clk),
	.d(\reset_reg[2]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(reset_reg_9),
	.prn(vcc));
defparam \reset_reg[9] .is_wysiwyg = "true";
defparam \reset_reg[9] .power_up = "low";

dffeas \reset_reg[12] (
	.clk(clk),
	.d(\reset_reg[2]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(reset_reg_12),
	.prn(vcc));
defparam \reset_reg[12] .is_wysiwyg = "true";
defparam \reset_reg[12] .power_up = "low";

dffeas \reset_reg[8] (
	.clk(clk),
	.d(\reset_reg[2]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(reset_reg_8),
	.prn(vcc));
defparam \reset_reg[8] .is_wysiwyg = "true";
defparam \reset_reg[8] .power_up = "low";

dffeas \reset_reg[10] (
	.clk(clk),
	.d(\reset_reg[2]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(reset_reg_10),
	.prn(vcc));
defparam \reset_reg[10] .is_wysiwyg = "true";
defparam \reset_reg[10] .power_up = "low";

dffeas \reset_reg[15] (
	.clk(clk),
	.d(\reset_reg[2]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(reset_reg_15),
	.prn(vcc));
defparam \reset_reg[15] .is_wysiwyg = "true";
defparam \reset_reg[15] .power_up = "low";

dffeas \reset_reg[0] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\reset_reg[0]~q ),
	.prn(vcc));
defparam \reset_reg[0] .is_wysiwyg = "true";
defparam \reset_reg[0] .power_up = "low";

dffeas \reset_reg[1] (
	.clk(clk),
	.d(\reset_reg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\reset_reg[1]~q ),
	.prn(vcc));
defparam \reset_reg[1] .is_wysiwyg = "true";
defparam \reset_reg[1] .power_up = "low";

dffeas \reset_reg[2] (
	.clk(clk),
	.d(\reset_reg[1]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\reset_reg[2]~q ),
	.prn(vcc));
defparam \reset_reg[2] .is_wysiwyg = "true";
defparam \reset_reg[2] .power_up = "low";

endmodule

module ddr3_int_alt_ddrx_input_if (
	clk_0,
	pipe_10_0,
	pipe_12_0,
	pipe_11_0,
	pipe_32_0,
	pipe_12_2,
	pipe_12_3,
	pipe_12_1,
	pipe_10_2,
	pipe_10_3,
	pipe_10_1,
	pipe_11_2,
	pipe_11_3,
	pipe_11_1,
	pipe_29_0,
	pipe_28_0,
	pipe_33_0,
	pipe_12_4,
	pipe_11_4,
	pipe_10_4,
	pipe_25_5,
	pipe_25_0,
	pipe_26_5,
	pipe_26_0,
	pipe_24_5,
	pipe_24_0,
	pipe_22_5,
	pipe_22_0,
	pipe_23_5,
	pipe_23_0,
	pipe_21_5,
	pipe_21_0,
	pipe_19_5,
	pipe_19_0,
	pipe_20_5,
	pipe_20_0,
	pipe_15_5,
	pipe_15_0,
	pipe_13_5,
	pipe_13_0,
	pipe_14_5,
	pipe_14_0,
	pipe_18_5,
	pipe_18_0,
	pipe_16_5,
	pipe_16_0,
	pipe_17_5,
	pipe_17_0,
	pipe_12_5,
	pipe_11_5,
	pipe_10_5,
	pipe_25_3,
	pipe_26_3,
	pipe_24_3,
	pipe_22_3,
	pipe_23_3,
	pipe_21_3,
	pipe_19_3,
	pipe_20_3,
	pipe_15_3,
	pipe_13_3,
	pipe_14_3,
	pipe_18_3,
	pipe_16_3,
	pipe_17_3,
	pipe_25_4,
	pipe_26_4,
	pipe_24_4,
	pipe_22_4,
	pipe_23_4,
	pipe_21_4,
	pipe_19_4,
	pipe_20_4,
	pipe_15_4,
	pipe_13_4,
	pipe_14_4,
	pipe_18_4,
	pipe_16_4,
	pipe_17_4,
	pipe_12_6,
	pipe_11_6,
	pipe_10_6,
	pipe_25_6,
	pipe_26_6,
	pipe_24_6,
	pipe_22_6,
	pipe_23_6,
	pipe_21_6,
	pipe_19_6,
	pipe_20_6,
	pipe_15_6,
	pipe_13_6,
	pipe_14_6,
	pipe_18_6,
	pipe_16_6,
	pipe_17_6,
	pipe_26_7,
	pipe_24_7,
	pipe_25_7,
	pipe_23_7,
	pipe_21_7,
	pipe_22_7,
	pipe_20_7,
	pipe_18_7,
	pipe_19_7,
	pipe_17_7,
	pipe_15_7,
	pipe_16_7,
	pipe_11_7,
	pipe_10_7,
	pipe_14_7,
	pipe_12_7,
	pipe_13_7,
	pipe_25_2,
	pipe_26_2,
	pipe_24_2,
	pipe_22_2,
	pipe_23_2,
	pipe_21_2,
	pipe_19_2,
	pipe_20_2,
	pipe_15_2,
	pipe_13_2,
	pipe_14_2,
	pipe_18_2,
	pipe_16_2,
	pipe_17_2,
	pipe_25_1,
	pipe_26_1,
	pipe_24_1,
	pipe_22_1,
	pipe_23_1,
	pipe_21_1,
	pipe_19_1,
	pipe_20_1,
	pipe_15_1,
	pipe_13_1,
	pipe_14_1,
	pipe_18_1,
	pipe_16_1,
	pipe_17_1,
	pipe_2_0,
	q_b_132,
	q_b_140,
	q_b_128,
	q_b_136,
	q_b_133,
	q_b_141,
	q_b_129,
	q_b_137,
	q_b_134,
	q_b_142,
	q_b_130,
	q_b_138,
	q_b_135,
	q_b_143,
	q_b_131,
	q_b_139,
	q_b_96,
	q_b_32,
	q_b_64,
	q_b_0,
	q_b_97,
	q_b_33,
	q_b_65,
	q_b_1,
	q_b_98,
	q_b_34,
	q_b_66,
	q_b_2,
	q_b_99,
	q_b_35,
	q_b_67,
	q_b_3,
	q_b_100,
	q_b_36,
	q_b_68,
	q_b_4,
	q_b_101,
	q_b_37,
	q_b_69,
	q_b_5,
	q_b_102,
	q_b_38,
	q_b_70,
	q_b_6,
	q_b_103,
	q_b_39,
	q_b_71,
	q_b_7,
	q_b_104,
	q_b_40,
	q_b_72,
	q_b_8,
	q_b_105,
	q_b_41,
	q_b_73,
	q_b_9,
	q_b_106,
	q_b_42,
	q_b_74,
	q_b_10,
	q_b_107,
	q_b_43,
	q_b_75,
	q_b_11,
	q_b_108,
	q_b_44,
	q_b_76,
	q_b_12,
	q_b_109,
	q_b_45,
	q_b_77,
	q_b_13,
	q_b_110,
	q_b_46,
	q_b_78,
	q_b_14,
	q_b_111,
	q_b_47,
	q_b_79,
	q_b_15,
	q_b_112,
	q_b_48,
	q_b_80,
	q_b_16,
	q_b_113,
	q_b_49,
	q_b_81,
	q_b_17,
	q_b_114,
	q_b_50,
	q_b_82,
	q_b_18,
	q_b_115,
	q_b_51,
	q_b_83,
	q_b_19,
	q_b_116,
	q_b_52,
	q_b_84,
	q_b_20,
	q_b_117,
	q_b_53,
	q_b_85,
	q_b_21,
	q_b_118,
	q_b_54,
	q_b_86,
	q_b_22,
	q_b_119,
	q_b_55,
	q_b_87,
	q_b_23,
	q_b_120,
	q_b_56,
	q_b_88,
	q_b_24,
	q_b_121,
	q_b_57,
	q_b_89,
	q_b_25,
	q_b_122,
	q_b_58,
	q_b_90,
	q_b_26,
	q_b_123,
	q_b_59,
	q_b_91,
	q_b_27,
	q_b_124,
	q_b_60,
	q_b_92,
	q_b_28,
	q_b_125,
	q_b_61,
	q_b_93,
	q_b_29,
	q_b_126,
	q_b_62,
	q_b_94,
	q_b_30,
	q_b_127,
	q_b_63,
	q_b_95,
	q_b_31,
	pipe_3_0,
	pipe_4_0,
	pipe_5_0,
	pipe_6_0,
	pipe_7_0,
	pipe_8_0,
	pipe_9_0,
	hold_ready,
	pipefull_7,
	ready_out,
	ctl_init_fail,
	ctl_init_success,
	local_init_done1,
	internal_ready,
	avalon_write_req,
	reset_reg_4,
	fetch,
	read_req,
	write_req,
	pipefull_6,
	reset_reg_5,
	ctl_reset_n,
	ecc_wdata_fifo_read,
	reset_reg_3,
	always38,
	pipefull_0,
	pipefull_5,
	pipefull_1,
	pipefull_4,
	pipefull_2,
	pipefull_3,
	GND_port,
	local_size_1,
	local_address_0,
	local_size_0,
	local_size_6,
	local_size_5,
	local_size_4,
	local_size_2,
	local_size_3,
	local_read_req,
	local_write_req,
	local_burstbegin,
	local_address_8,
	local_address_10,
	local_address_9,
	local_address_23,
	local_address_24,
	local_address_22,
	local_address_20,
	local_address_21,
	local_address_19,
	local_address_17,
	local_address_18,
	local_address_13,
	local_address_11,
	local_address_12,
	local_address_16,
	local_address_14,
	local_address_15,
	local_address_1,
	local_address_2,
	local_address_3,
	local_address_4,
	local_address_5,
	local_address_7,
	local_address_6,
	local_be_4,
	local_be_12,
	local_be_0,
	local_be_8,
	local_be_5,
	local_be_13,
	local_be_1,
	local_be_9,
	local_be_6,
	local_be_14,
	local_be_2,
	local_be_10,
	local_be_7,
	local_be_15,
	local_be_3,
	local_be_11,
	local_wdata_96,
	local_wdata_32,
	local_wdata_64,
	local_wdata_0,
	local_wdata_97,
	local_wdata_33,
	local_wdata_65,
	local_wdata_1,
	local_wdata_98,
	local_wdata_34,
	local_wdata_66,
	local_wdata_2,
	local_wdata_99,
	local_wdata_35,
	local_wdata_67,
	local_wdata_3,
	local_wdata_100,
	local_wdata_36,
	local_wdata_68,
	local_wdata_4,
	local_wdata_101,
	local_wdata_37,
	local_wdata_69,
	local_wdata_5,
	local_wdata_102,
	local_wdata_38,
	local_wdata_70,
	local_wdata_6,
	local_wdata_103,
	local_wdata_39,
	local_wdata_71,
	local_wdata_7,
	local_wdata_104,
	local_wdata_40,
	local_wdata_72,
	local_wdata_8,
	local_wdata_105,
	local_wdata_41,
	local_wdata_73,
	local_wdata_9,
	local_wdata_106,
	local_wdata_42,
	local_wdata_74,
	local_wdata_10,
	local_wdata_107,
	local_wdata_43,
	local_wdata_75,
	local_wdata_11,
	local_wdata_108,
	local_wdata_44,
	local_wdata_76,
	local_wdata_12,
	local_wdata_109,
	local_wdata_45,
	local_wdata_77,
	local_wdata_13,
	local_wdata_110,
	local_wdata_46,
	local_wdata_78,
	local_wdata_14,
	local_wdata_111,
	local_wdata_47,
	local_wdata_79,
	local_wdata_15,
	local_wdata_112,
	local_wdata_48,
	local_wdata_80,
	local_wdata_16,
	local_wdata_113,
	local_wdata_49,
	local_wdata_81,
	local_wdata_17,
	local_wdata_114,
	local_wdata_50,
	local_wdata_82,
	local_wdata_18,
	local_wdata_115,
	local_wdata_51,
	local_wdata_83,
	local_wdata_19,
	local_wdata_116,
	local_wdata_52,
	local_wdata_84,
	local_wdata_20,
	local_wdata_117,
	local_wdata_53,
	local_wdata_85,
	local_wdata_21,
	local_wdata_118,
	local_wdata_54,
	local_wdata_86,
	local_wdata_22,
	local_wdata_119,
	local_wdata_55,
	local_wdata_87,
	local_wdata_23,
	local_wdata_120,
	local_wdata_56,
	local_wdata_88,
	local_wdata_24,
	local_wdata_121,
	local_wdata_57,
	local_wdata_89,
	local_wdata_25,
	local_wdata_122,
	local_wdata_58,
	local_wdata_90,
	local_wdata_26,
	local_wdata_123,
	local_wdata_59,
	local_wdata_91,
	local_wdata_27,
	local_wdata_124,
	local_wdata_60,
	local_wdata_92,
	local_wdata_28,
	local_wdata_125,
	local_wdata_61,
	local_wdata_93,
	local_wdata_29,
	local_wdata_126,
	local_wdata_62,
	local_wdata_94,
	local_wdata_30,
	local_wdata_127,
	local_wdata_63,
	local_wdata_95,
	local_wdata_31)/* synthesis synthesis_greybox=0 */;
input 	clk_0;
output 	pipe_10_0;
output 	pipe_12_0;
output 	pipe_11_0;
output 	pipe_32_0;
output 	pipe_12_2;
output 	pipe_12_3;
output 	pipe_12_1;
output 	pipe_10_2;
output 	pipe_10_3;
output 	pipe_10_1;
output 	pipe_11_2;
output 	pipe_11_3;
output 	pipe_11_1;
output 	pipe_29_0;
output 	pipe_28_0;
output 	pipe_33_0;
output 	pipe_12_4;
output 	pipe_11_4;
output 	pipe_10_4;
output 	pipe_25_5;
output 	pipe_25_0;
output 	pipe_26_5;
output 	pipe_26_0;
output 	pipe_24_5;
output 	pipe_24_0;
output 	pipe_22_5;
output 	pipe_22_0;
output 	pipe_23_5;
output 	pipe_23_0;
output 	pipe_21_5;
output 	pipe_21_0;
output 	pipe_19_5;
output 	pipe_19_0;
output 	pipe_20_5;
output 	pipe_20_0;
output 	pipe_15_5;
output 	pipe_15_0;
output 	pipe_13_5;
output 	pipe_13_0;
output 	pipe_14_5;
output 	pipe_14_0;
output 	pipe_18_5;
output 	pipe_18_0;
output 	pipe_16_5;
output 	pipe_16_0;
output 	pipe_17_5;
output 	pipe_17_0;
output 	pipe_12_5;
output 	pipe_11_5;
output 	pipe_10_5;
output 	pipe_25_3;
output 	pipe_26_3;
output 	pipe_24_3;
output 	pipe_22_3;
output 	pipe_23_3;
output 	pipe_21_3;
output 	pipe_19_3;
output 	pipe_20_3;
output 	pipe_15_3;
output 	pipe_13_3;
output 	pipe_14_3;
output 	pipe_18_3;
output 	pipe_16_3;
output 	pipe_17_3;
output 	pipe_25_4;
output 	pipe_26_4;
output 	pipe_24_4;
output 	pipe_22_4;
output 	pipe_23_4;
output 	pipe_21_4;
output 	pipe_19_4;
output 	pipe_20_4;
output 	pipe_15_4;
output 	pipe_13_4;
output 	pipe_14_4;
output 	pipe_18_4;
output 	pipe_16_4;
output 	pipe_17_4;
output 	pipe_12_6;
output 	pipe_11_6;
output 	pipe_10_6;
output 	pipe_25_6;
output 	pipe_26_6;
output 	pipe_24_6;
output 	pipe_22_6;
output 	pipe_23_6;
output 	pipe_21_6;
output 	pipe_19_6;
output 	pipe_20_6;
output 	pipe_15_6;
output 	pipe_13_6;
output 	pipe_14_6;
output 	pipe_18_6;
output 	pipe_16_6;
output 	pipe_17_6;
output 	pipe_26_7;
output 	pipe_24_7;
output 	pipe_25_7;
output 	pipe_23_7;
output 	pipe_21_7;
output 	pipe_22_7;
output 	pipe_20_7;
output 	pipe_18_7;
output 	pipe_19_7;
output 	pipe_17_7;
output 	pipe_15_7;
output 	pipe_16_7;
output 	pipe_11_7;
output 	pipe_10_7;
output 	pipe_14_7;
output 	pipe_12_7;
output 	pipe_13_7;
output 	pipe_25_2;
output 	pipe_26_2;
output 	pipe_24_2;
output 	pipe_22_2;
output 	pipe_23_2;
output 	pipe_21_2;
output 	pipe_19_2;
output 	pipe_20_2;
output 	pipe_15_2;
output 	pipe_13_2;
output 	pipe_14_2;
output 	pipe_18_2;
output 	pipe_16_2;
output 	pipe_17_2;
output 	pipe_25_1;
output 	pipe_26_1;
output 	pipe_24_1;
output 	pipe_22_1;
output 	pipe_23_1;
output 	pipe_21_1;
output 	pipe_19_1;
output 	pipe_20_1;
output 	pipe_15_1;
output 	pipe_13_1;
output 	pipe_14_1;
output 	pipe_18_1;
output 	pipe_16_1;
output 	pipe_17_1;
output 	pipe_2_0;
output 	q_b_132;
output 	q_b_140;
output 	q_b_128;
output 	q_b_136;
output 	q_b_133;
output 	q_b_141;
output 	q_b_129;
output 	q_b_137;
output 	q_b_134;
output 	q_b_142;
output 	q_b_130;
output 	q_b_138;
output 	q_b_135;
output 	q_b_143;
output 	q_b_131;
output 	q_b_139;
output 	q_b_96;
output 	q_b_32;
output 	q_b_64;
output 	q_b_0;
output 	q_b_97;
output 	q_b_33;
output 	q_b_65;
output 	q_b_1;
output 	q_b_98;
output 	q_b_34;
output 	q_b_66;
output 	q_b_2;
output 	q_b_99;
output 	q_b_35;
output 	q_b_67;
output 	q_b_3;
output 	q_b_100;
output 	q_b_36;
output 	q_b_68;
output 	q_b_4;
output 	q_b_101;
output 	q_b_37;
output 	q_b_69;
output 	q_b_5;
output 	q_b_102;
output 	q_b_38;
output 	q_b_70;
output 	q_b_6;
output 	q_b_103;
output 	q_b_39;
output 	q_b_71;
output 	q_b_7;
output 	q_b_104;
output 	q_b_40;
output 	q_b_72;
output 	q_b_8;
output 	q_b_105;
output 	q_b_41;
output 	q_b_73;
output 	q_b_9;
output 	q_b_106;
output 	q_b_42;
output 	q_b_74;
output 	q_b_10;
output 	q_b_107;
output 	q_b_43;
output 	q_b_75;
output 	q_b_11;
output 	q_b_108;
output 	q_b_44;
output 	q_b_76;
output 	q_b_12;
output 	q_b_109;
output 	q_b_45;
output 	q_b_77;
output 	q_b_13;
output 	q_b_110;
output 	q_b_46;
output 	q_b_78;
output 	q_b_14;
output 	q_b_111;
output 	q_b_47;
output 	q_b_79;
output 	q_b_15;
output 	q_b_112;
output 	q_b_48;
output 	q_b_80;
output 	q_b_16;
output 	q_b_113;
output 	q_b_49;
output 	q_b_81;
output 	q_b_17;
output 	q_b_114;
output 	q_b_50;
output 	q_b_82;
output 	q_b_18;
output 	q_b_115;
output 	q_b_51;
output 	q_b_83;
output 	q_b_19;
output 	q_b_116;
output 	q_b_52;
output 	q_b_84;
output 	q_b_20;
output 	q_b_117;
output 	q_b_53;
output 	q_b_85;
output 	q_b_21;
output 	q_b_118;
output 	q_b_54;
output 	q_b_86;
output 	q_b_22;
output 	q_b_119;
output 	q_b_55;
output 	q_b_87;
output 	q_b_23;
output 	q_b_120;
output 	q_b_56;
output 	q_b_88;
output 	q_b_24;
output 	q_b_121;
output 	q_b_57;
output 	q_b_89;
output 	q_b_25;
output 	q_b_122;
output 	q_b_58;
output 	q_b_90;
output 	q_b_26;
output 	q_b_123;
output 	q_b_59;
output 	q_b_91;
output 	q_b_27;
output 	q_b_124;
output 	q_b_60;
output 	q_b_92;
output 	q_b_28;
output 	q_b_125;
output 	q_b_61;
output 	q_b_93;
output 	q_b_29;
output 	q_b_126;
output 	q_b_62;
output 	q_b_94;
output 	q_b_30;
output 	q_b_127;
output 	q_b_63;
output 	q_b_95;
output 	q_b_31;
output 	pipe_3_0;
output 	pipe_4_0;
output 	pipe_5_0;
output 	pipe_6_0;
output 	pipe_7_0;
output 	pipe_8_0;
output 	pipe_9_0;
output 	hold_ready;
output 	pipefull_7;
output 	ready_out;
input 	ctl_init_fail;
input 	ctl_init_success;
output 	local_init_done1;
output 	internal_ready;
output 	avalon_write_req;
input 	reset_reg_4;
input 	fetch;
output 	read_req;
output 	write_req;
output 	pipefull_6;
input 	reset_reg_5;
input 	[4:0] ctl_reset_n;
input 	ecc_wdata_fifo_read;
input 	reset_reg_3;
input 	always38;
output 	pipefull_0;
output 	pipefull_5;
output 	pipefull_1;
output 	pipefull_4;
output 	pipefull_2;
output 	pipefull_3;
input 	GND_port;
input 	local_size_1;
input 	local_address_0;
input 	local_size_0;
input 	local_size_6;
input 	local_size_5;
input 	local_size_4;
input 	local_size_2;
input 	local_size_3;
input 	local_read_req;
input 	local_write_req;
input 	local_burstbegin;
input 	local_address_8;
input 	local_address_10;
input 	local_address_9;
input 	local_address_23;
input 	local_address_24;
input 	local_address_22;
input 	local_address_20;
input 	local_address_21;
input 	local_address_19;
input 	local_address_17;
input 	local_address_18;
input 	local_address_13;
input 	local_address_11;
input 	local_address_12;
input 	local_address_16;
input 	local_address_14;
input 	local_address_15;
input 	local_address_1;
input 	local_address_2;
input 	local_address_3;
input 	local_address_4;
input 	local_address_5;
input 	local_address_7;
input 	local_address_6;
input 	local_be_4;
input 	local_be_12;
input 	local_be_0;
input 	local_be_8;
input 	local_be_5;
input 	local_be_13;
input 	local_be_1;
input 	local_be_9;
input 	local_be_6;
input 	local_be_14;
input 	local_be_2;
input 	local_be_10;
input 	local_be_7;
input 	local_be_15;
input 	local_be_3;
input 	local_be_11;
input 	local_wdata_96;
input 	local_wdata_32;
input 	local_wdata_64;
input 	local_wdata_0;
input 	local_wdata_97;
input 	local_wdata_33;
input 	local_wdata_65;
input 	local_wdata_1;
input 	local_wdata_98;
input 	local_wdata_34;
input 	local_wdata_66;
input 	local_wdata_2;
input 	local_wdata_99;
input 	local_wdata_35;
input 	local_wdata_67;
input 	local_wdata_3;
input 	local_wdata_100;
input 	local_wdata_36;
input 	local_wdata_68;
input 	local_wdata_4;
input 	local_wdata_101;
input 	local_wdata_37;
input 	local_wdata_69;
input 	local_wdata_5;
input 	local_wdata_102;
input 	local_wdata_38;
input 	local_wdata_70;
input 	local_wdata_6;
input 	local_wdata_103;
input 	local_wdata_39;
input 	local_wdata_71;
input 	local_wdata_7;
input 	local_wdata_104;
input 	local_wdata_40;
input 	local_wdata_72;
input 	local_wdata_8;
input 	local_wdata_105;
input 	local_wdata_41;
input 	local_wdata_73;
input 	local_wdata_9;
input 	local_wdata_106;
input 	local_wdata_42;
input 	local_wdata_74;
input 	local_wdata_10;
input 	local_wdata_107;
input 	local_wdata_43;
input 	local_wdata_75;
input 	local_wdata_11;
input 	local_wdata_108;
input 	local_wdata_44;
input 	local_wdata_76;
input 	local_wdata_12;
input 	local_wdata_109;
input 	local_wdata_45;
input 	local_wdata_77;
input 	local_wdata_13;
input 	local_wdata_110;
input 	local_wdata_46;
input 	local_wdata_78;
input 	local_wdata_14;
input 	local_wdata_111;
input 	local_wdata_47;
input 	local_wdata_79;
input 	local_wdata_15;
input 	local_wdata_112;
input 	local_wdata_48;
input 	local_wdata_80;
input 	local_wdata_16;
input 	local_wdata_113;
input 	local_wdata_49;
input 	local_wdata_81;
input 	local_wdata_17;
input 	local_wdata_114;
input 	local_wdata_50;
input 	local_wdata_82;
input 	local_wdata_18;
input 	local_wdata_115;
input 	local_wdata_51;
input 	local_wdata_83;
input 	local_wdata_19;
input 	local_wdata_116;
input 	local_wdata_52;
input 	local_wdata_84;
input 	local_wdata_20;
input 	local_wdata_117;
input 	local_wdata_53;
input 	local_wdata_85;
input 	local_wdata_21;
input 	local_wdata_118;
input 	local_wdata_54;
input 	local_wdata_86;
input 	local_wdata_22;
input 	local_wdata_119;
input 	local_wdata_55;
input 	local_wdata_87;
input 	local_wdata_23;
input 	local_wdata_120;
input 	local_wdata_56;
input 	local_wdata_88;
input 	local_wdata_24;
input 	local_wdata_121;
input 	local_wdata_57;
input 	local_wdata_89;
input 	local_wdata_25;
input 	local_wdata_122;
input 	local_wdata_58;
input 	local_wdata_90;
input 	local_wdata_26;
input 	local_wdata_123;
input 	local_wdata_59;
input 	local_wdata_91;
input 	local_wdata_27;
input 	local_wdata_124;
input 	local_wdata_60;
input 	local_wdata_92;
input 	local_wdata_28;
input 	local_wdata_125;
input 	local_wdata_61;
input 	local_wdata_93;
input 	local_wdata_29;
input 	local_wdata_126;
input 	local_wdata_62;
input 	local_wdata_94;
input 	local_wdata_30;
input 	local_wdata_127;
input 	local_wdata_63;
input 	local_wdata_95;
input 	local_wdata_31;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \cmd_gen_inst|buf_bank_addr[0]~q ;
wire \cmd_gen_inst|buf_bank_addr[2]~q ;
wire \cmd_gen_inst|buf_bank_addr[1]~q ;
wire \cmd_gen_inst|buf_col_addr[3]~q ;
wire \cmd_gen_inst|buf_col_addr[4]~q ;
wire \cmd_gen_inst|buf_col_addr[5]~q ;
wire \cmd_gen_inst|buf_col_addr[6]~q ;
wire \cmd_gen_inst|buf_col_addr[7]~q ;
wire \cmd_gen_inst|buf_col_addr[9]~q ;
wire \cmd_gen_inst|buf_col_addr[8]~q ;
wire \cmd_gen_inst|buf_row_addr[12]~q ;
wire \cmd_gen_inst|buf_row_addr[13]~q ;
wire \cmd_gen_inst|buf_row_addr[11]~q ;
wire \cmd_gen_inst|buf_row_addr[9]~q ;
wire \cmd_gen_inst|buf_row_addr[10]~q ;
wire \cmd_gen_inst|buf_row_addr[8]~q ;
wire \cmd_gen_inst|buf_row_addr[6]~q ;
wire \cmd_gen_inst|buf_row_addr[7]~q ;
wire \cmd_gen_inst|buf_row_addr[2]~q ;
wire \cmd_gen_inst|buf_row_addr[0]~q ;
wire \cmd_gen_inst|buf_row_addr[1]~q ;
wire \cmd_gen_inst|buf_row_addr[5]~q ;
wire \cmd_gen_inst|buf_row_addr[3]~q ;
wire \cmd_gen_inst|buf_row_addr[4]~q ;
wire \wdata_fifo_inst|wdata_fifo|auto_generated|dffe_af~q ;
wire \avalon_if_inst|avalon_read_req~combout ;
wire \prolong_burstbegin~q ;
wire \cmd_gen_inst|generating~q ;
wire \prolong_burstbegin~0_combout ;
wire \cmd_gen_inst|bank_addr[0]~0_combout ;
wire \cmd_gen_inst|bank_addr[2]~1_combout ;
wire \cmd_gen_inst|bank_addr[1]~2_combout ;
wire \cmd_gen_inst|size[1]~0_combout ;
wire \cmd_gen_inst|size[0]~1_combout ;
wire \cmd_gen_inst|row_addr[12]~0_combout ;
wire \cmd_gen_inst|row_addr[13]~1_combout ;
wire \cmd_gen_inst|row_addr[11]~2_combout ;
wire \cmd_gen_inst|row_addr[9]~3_combout ;
wire \cmd_gen_inst|row_addr[10]~4_combout ;
wire \cmd_gen_inst|row_addr[8]~5_combout ;
wire \cmd_gen_inst|row_addr[6]~6_combout ;
wire \cmd_gen_inst|row_addr[7]~7_combout ;
wire \cmd_gen_inst|row_addr[2]~8_combout ;
wire \cmd_gen_inst|row_addr[0]~9_combout ;
wire \cmd_gen_inst|row_addr[1]~10_combout ;
wire \cmd_gen_inst|row_addr[5]~11_combout ;
wire \cmd_gen_inst|row_addr[3]~12_combout ;
wire \cmd_gen_inst|row_addr[4]~13_combout ;
wire \cmd_gen_inst|col_addr[2]~0_combout ;
wire \cmd_gen_inst|col_addr[3]~1_combout ;
wire \cmd_gen_inst|col_addr[4]~2_combout ;
wire \cmd_gen_inst|col_addr[5]~3_combout ;
wire \cmd_gen_inst|col_addr[6]~4_combout ;
wire \cmd_gen_inst|col_addr[7]~5_combout ;
wire \cmd_gen_inst|col_addr[8]~6_combout ;
wire \cmd_gen_inst|col_addr[9]~7_combout ;
wire \gate_ready_in_reset~q ;


ddr3_int_alt_ddrx_cmd_queue cmd_queue_inst(
	.ctl_clk(clk_0),
	.pipe_10_0(pipe_10_0),
	.pipe_12_0(pipe_12_0),
	.pipe_11_0(pipe_11_0),
	.pipe_32_0(pipe_32_0),
	.pipe_12_2(pipe_12_2),
	.pipe_12_3(pipe_12_3),
	.pipe_12_1(pipe_12_1),
	.pipe_10_2(pipe_10_2),
	.pipe_10_3(pipe_10_3),
	.pipe_10_1(pipe_10_1),
	.pipe_11_2(pipe_11_2),
	.pipe_11_3(pipe_11_3),
	.pipe_11_1(pipe_11_1),
	.pipe_29_0(pipe_29_0),
	.pipe_28_0(pipe_28_0),
	.pipe_33_0(pipe_33_0),
	.pipe_12_4(pipe_12_4),
	.pipe_11_4(pipe_11_4),
	.pipe_10_4(pipe_10_4),
	.buf_bank_addr_0(\cmd_gen_inst|buf_bank_addr[0]~q ),
	.buf_bank_addr_2(\cmd_gen_inst|buf_bank_addr[2]~q ),
	.buf_bank_addr_1(\cmd_gen_inst|buf_bank_addr[1]~q ),
	.pipe_25_5(pipe_25_5),
	.pipe_25_0(pipe_25_0),
	.pipe_26_5(pipe_26_5),
	.pipe_26_0(pipe_26_0),
	.pipe_24_5(pipe_24_5),
	.pipe_24_0(pipe_24_0),
	.pipe_22_5(pipe_22_5),
	.pipe_22_0(pipe_22_0),
	.pipe_23_5(pipe_23_5),
	.pipe_23_0(pipe_23_0),
	.pipe_21_5(pipe_21_5),
	.pipe_21_0(pipe_21_0),
	.pipe_19_5(pipe_19_5),
	.pipe_19_0(pipe_19_0),
	.pipe_20_5(pipe_20_5),
	.pipe_20_0(pipe_20_0),
	.pipe_15_5(pipe_15_5),
	.pipe_15_0(pipe_15_0),
	.pipe_13_5(pipe_13_5),
	.pipe_13_0(pipe_13_0),
	.pipe_14_5(pipe_14_5),
	.pipe_14_0(pipe_14_0),
	.pipe_18_5(pipe_18_5),
	.pipe_18_0(pipe_18_0),
	.pipe_16_5(pipe_16_5),
	.pipe_16_0(pipe_16_0),
	.pipe_17_5(pipe_17_5),
	.pipe_17_0(pipe_17_0),
	.pipe_12_5(pipe_12_5),
	.pipe_11_5(pipe_11_5),
	.pipe_10_5(pipe_10_5),
	.pipe_25_3(pipe_25_3),
	.pipe_26_3(pipe_26_3),
	.pipe_24_3(pipe_24_3),
	.pipe_22_3(pipe_22_3),
	.pipe_23_3(pipe_23_3),
	.pipe_21_3(pipe_21_3),
	.pipe_19_3(pipe_19_3),
	.pipe_20_3(pipe_20_3),
	.pipe_15_3(pipe_15_3),
	.pipe_13_3(pipe_13_3),
	.pipe_14_3(pipe_14_3),
	.pipe_18_3(pipe_18_3),
	.pipe_16_3(pipe_16_3),
	.pipe_17_3(pipe_17_3),
	.pipe_25_4(pipe_25_4),
	.pipe_26_4(pipe_26_4),
	.pipe_24_4(pipe_24_4),
	.pipe_22_4(pipe_22_4),
	.pipe_23_4(pipe_23_4),
	.pipe_21_4(pipe_21_4),
	.pipe_19_4(pipe_19_4),
	.pipe_20_4(pipe_20_4),
	.pipe_15_4(pipe_15_4),
	.pipe_13_4(pipe_13_4),
	.pipe_14_4(pipe_14_4),
	.pipe_18_4(pipe_18_4),
	.pipe_16_4(pipe_16_4),
	.pipe_17_4(pipe_17_4),
	.pipe_12_6(pipe_12_6),
	.pipe_11_6(pipe_11_6),
	.pipe_10_6(pipe_10_6),
	.pipe_25_6(pipe_25_6),
	.pipe_26_6(pipe_26_6),
	.pipe_24_6(pipe_24_6),
	.pipe_22_6(pipe_22_6),
	.pipe_23_6(pipe_23_6),
	.pipe_21_6(pipe_21_6),
	.pipe_19_6(pipe_19_6),
	.pipe_20_6(pipe_20_6),
	.pipe_15_6(pipe_15_6),
	.pipe_13_6(pipe_13_6),
	.pipe_14_6(pipe_14_6),
	.pipe_18_6(pipe_18_6),
	.pipe_16_6(pipe_16_6),
	.pipe_17_6(pipe_17_6),
	.pipe_26_7(pipe_26_7),
	.pipe_24_7(pipe_24_7),
	.pipe_25_7(pipe_25_7),
	.pipe_23_7(pipe_23_7),
	.pipe_21_7(pipe_21_7),
	.pipe_22_7(pipe_22_7),
	.pipe_20_7(pipe_20_7),
	.pipe_18_7(pipe_18_7),
	.pipe_19_7(pipe_19_7),
	.pipe_17_7(pipe_17_7),
	.pipe_15_7(pipe_15_7),
	.pipe_16_7(pipe_16_7),
	.pipe_11_7(pipe_11_7),
	.pipe_10_7(pipe_10_7),
	.pipe_14_7(pipe_14_7),
	.pipe_12_7(pipe_12_7),
	.pipe_13_7(pipe_13_7),
	.pipe_25_2(pipe_25_2),
	.pipe_26_2(pipe_26_2),
	.pipe_24_2(pipe_24_2),
	.pipe_22_2(pipe_22_2),
	.pipe_23_2(pipe_23_2),
	.pipe_21_2(pipe_21_2),
	.pipe_19_2(pipe_19_2),
	.pipe_20_2(pipe_20_2),
	.pipe_15_2(pipe_15_2),
	.pipe_13_2(pipe_13_2),
	.pipe_14_2(pipe_14_2),
	.pipe_18_2(pipe_18_2),
	.pipe_16_2(pipe_16_2),
	.pipe_17_2(pipe_17_2),
	.pipe_25_1(pipe_25_1),
	.pipe_26_1(pipe_26_1),
	.pipe_24_1(pipe_24_1),
	.pipe_22_1(pipe_22_1),
	.pipe_23_1(pipe_23_1),
	.pipe_21_1(pipe_21_1),
	.pipe_19_1(pipe_19_1),
	.pipe_20_1(pipe_20_1),
	.pipe_15_1(pipe_15_1),
	.pipe_13_1(pipe_13_1),
	.pipe_14_1(pipe_14_1),
	.pipe_18_1(pipe_18_1),
	.pipe_16_1(pipe_16_1),
	.pipe_17_1(pipe_17_1),
	.buf_col_addr_3(\cmd_gen_inst|buf_col_addr[3]~q ),
	.buf_col_addr_4(\cmd_gen_inst|buf_col_addr[4]~q ),
	.buf_col_addr_5(\cmd_gen_inst|buf_col_addr[5]~q ),
	.buf_col_addr_6(\cmd_gen_inst|buf_col_addr[6]~q ),
	.buf_col_addr_7(\cmd_gen_inst|buf_col_addr[7]~q ),
	.buf_col_addr_9(\cmd_gen_inst|buf_col_addr[9]~q ),
	.buf_col_addr_8(\cmd_gen_inst|buf_col_addr[8]~q ),
	.buf_row_addr_12(\cmd_gen_inst|buf_row_addr[12]~q ),
	.buf_row_addr_13(\cmd_gen_inst|buf_row_addr[13]~q ),
	.buf_row_addr_11(\cmd_gen_inst|buf_row_addr[11]~q ),
	.buf_row_addr_9(\cmd_gen_inst|buf_row_addr[9]~q ),
	.buf_row_addr_10(\cmd_gen_inst|buf_row_addr[10]~q ),
	.buf_row_addr_8(\cmd_gen_inst|buf_row_addr[8]~q ),
	.buf_row_addr_6(\cmd_gen_inst|buf_row_addr[6]~q ),
	.buf_row_addr_7(\cmd_gen_inst|buf_row_addr[7]~q ),
	.buf_row_addr_2(\cmd_gen_inst|buf_row_addr[2]~q ),
	.buf_row_addr_0(\cmd_gen_inst|buf_row_addr[0]~q ),
	.buf_row_addr_1(\cmd_gen_inst|buf_row_addr[1]~q ),
	.buf_row_addr_5(\cmd_gen_inst|buf_row_addr[5]~q ),
	.buf_row_addr_3(\cmd_gen_inst|buf_row_addr[3]~q ),
	.buf_row_addr_4(\cmd_gen_inst|buf_row_addr[4]~q ),
	.pipe_2_0(pipe_2_0),
	.pipe_3_0(pipe_3_0),
	.pipe_4_0(pipe_4_0),
	.pipe_5_0(pipe_5_0),
	.pipe_6_0(pipe_6_0),
	.pipe_7_0(pipe_7_0),
	.pipe_8_0(pipe_8_0),
	.pipe_9_0(pipe_9_0),
	.pipefull_7(pipefull_7),
	.generating(\cmd_gen_inst|generating~q ),
	.fetch(fetch),
	.read_req(read_req),
	.write_req(write_req),
	.pipefull_6(pipefull_6),
	.ctl_reset_n(reset_reg_5),
	.always38(always38),
	.pipefull_0(pipefull_0),
	.pipefull_5(pipefull_5),
	.pipefull_1(pipefull_1),
	.pipefull_4(pipefull_4),
	.pipefull_2(pipefull_2),
	.pipefull_3(pipefull_3),
	.bank_addr_0(\cmd_gen_inst|bank_addr[0]~0_combout ),
	.bank_addr_2(\cmd_gen_inst|bank_addr[2]~1_combout ),
	.bank_addr_1(\cmd_gen_inst|bank_addr[1]~2_combout ),
	.size_1(\cmd_gen_inst|size[1]~0_combout ),
	.size_0(\cmd_gen_inst|size[0]~1_combout ),
	.row_addr_12(\cmd_gen_inst|row_addr[12]~0_combout ),
	.row_addr_13(\cmd_gen_inst|row_addr[13]~1_combout ),
	.row_addr_11(\cmd_gen_inst|row_addr[11]~2_combout ),
	.row_addr_9(\cmd_gen_inst|row_addr[9]~3_combout ),
	.row_addr_10(\cmd_gen_inst|row_addr[10]~4_combout ),
	.row_addr_8(\cmd_gen_inst|row_addr[8]~5_combout ),
	.row_addr_6(\cmd_gen_inst|row_addr[6]~6_combout ),
	.row_addr_7(\cmd_gen_inst|row_addr[7]~7_combout ),
	.row_addr_2(\cmd_gen_inst|row_addr[2]~8_combout ),
	.row_addr_0(\cmd_gen_inst|row_addr[0]~9_combout ),
	.row_addr_1(\cmd_gen_inst|row_addr[1]~10_combout ),
	.row_addr_5(\cmd_gen_inst|row_addr[5]~11_combout ),
	.row_addr_3(\cmd_gen_inst|row_addr[3]~12_combout ),
	.row_addr_4(\cmd_gen_inst|row_addr[4]~13_combout ),
	.col_addr_2(\cmd_gen_inst|col_addr[2]~0_combout ),
	.col_addr_3(\cmd_gen_inst|col_addr[3]~1_combout ),
	.col_addr_4(\cmd_gen_inst|col_addr[4]~2_combout ),
	.col_addr_5(\cmd_gen_inst|col_addr[5]~3_combout ),
	.col_addr_6(\cmd_gen_inst|col_addr[6]~4_combout ),
	.col_addr_7(\cmd_gen_inst|col_addr[7]~5_combout ),
	.col_addr_8(\cmd_gen_inst|col_addr[8]~6_combout ),
	.col_addr_9(\cmd_gen_inst|col_addr[9]~7_combout ),
	.local_address_0(local_address_0),
	.local_address_8(local_address_8),
	.local_address_10(local_address_10),
	.local_address_9(local_address_9),
	.local_address_23(local_address_23),
	.local_address_24(local_address_24),
	.local_address_22(local_address_22),
	.local_address_20(local_address_20),
	.local_address_21(local_address_21),
	.local_address_19(local_address_19),
	.local_address_17(local_address_17),
	.local_address_18(local_address_18),
	.local_address_13(local_address_13),
	.local_address_11(local_address_11),
	.local_address_12(local_address_12),
	.local_address_16(local_address_16),
	.local_address_14(local_address_14),
	.local_address_15(local_address_15),
	.local_address_1(local_address_1),
	.local_address_2(local_address_2),
	.local_address_3(local_address_3),
	.local_address_4(local_address_4),
	.local_address_5(local_address_5),
	.local_address_7(local_address_7),
	.local_address_6(local_address_6));

ddr3_int_alt_ddrx_avalon_if avalon_if_inst(
	.hold_ready(hold_ready),
	.pipefull_7(pipefull_7),
	.gate_ready_in_reset(\gate_ready_in_reset~q ),
	.dffe_af(\wdata_fifo_inst|wdata_fifo|auto_generated|dffe_af~q ),
	.avalon_read_req1(\avalon_if_inst|avalon_read_req~combout ),
	.avalon_write_req1(avalon_write_req),
	.local_read_req(local_read_req),
	.local_write_req(local_write_req));

ddr3_int_alt_ddrx_cmd_gen cmd_gen_inst(
	.ctl_clk(clk_0),
	.buf_bank_addr_0(\cmd_gen_inst|buf_bank_addr[0]~q ),
	.buf_bank_addr_2(\cmd_gen_inst|buf_bank_addr[2]~q ),
	.buf_bank_addr_1(\cmd_gen_inst|buf_bank_addr[1]~q ),
	.buf_col_addr_3(\cmd_gen_inst|buf_col_addr[3]~q ),
	.buf_col_addr_4(\cmd_gen_inst|buf_col_addr[4]~q ),
	.buf_col_addr_5(\cmd_gen_inst|buf_col_addr[5]~q ),
	.buf_col_addr_6(\cmd_gen_inst|buf_col_addr[6]~q ),
	.buf_col_addr_7(\cmd_gen_inst|buf_col_addr[7]~q ),
	.buf_col_addr_9(\cmd_gen_inst|buf_col_addr[9]~q ),
	.buf_col_addr_8(\cmd_gen_inst|buf_col_addr[8]~q ),
	.buf_row_addr_12(\cmd_gen_inst|buf_row_addr[12]~q ),
	.buf_row_addr_13(\cmd_gen_inst|buf_row_addr[13]~q ),
	.buf_row_addr_11(\cmd_gen_inst|buf_row_addr[11]~q ),
	.buf_row_addr_9(\cmd_gen_inst|buf_row_addr[9]~q ),
	.buf_row_addr_10(\cmd_gen_inst|buf_row_addr[10]~q ),
	.buf_row_addr_8(\cmd_gen_inst|buf_row_addr[8]~q ),
	.buf_row_addr_6(\cmd_gen_inst|buf_row_addr[6]~q ),
	.buf_row_addr_7(\cmd_gen_inst|buf_row_addr[7]~q ),
	.buf_row_addr_2(\cmd_gen_inst|buf_row_addr[2]~q ),
	.buf_row_addr_0(\cmd_gen_inst|buf_row_addr[0]~q ),
	.buf_row_addr_1(\cmd_gen_inst|buf_row_addr[1]~q ),
	.buf_row_addr_5(\cmd_gen_inst|buf_row_addr[5]~q ),
	.buf_row_addr_3(\cmd_gen_inst|buf_row_addr[3]~q ),
	.buf_row_addr_4(\cmd_gen_inst|buf_row_addr[4]~q ),
	.hold_ready1(hold_ready),
	.pipefull_7(pipefull_7),
	.gate_ready_in_reset(\gate_ready_in_reset~q ),
	.dffe_af(\wdata_fifo_inst|wdata_fifo|auto_generated|dffe_af~q ),
	.ready_out1(ready_out),
	.internal_ready(internal_ready),
	.local_read_req(\avalon_if_inst|avalon_read_req~combout ),
	.local_write_req(avalon_write_req),
	.prolong_burstbegin(\prolong_burstbegin~q ),
	.generating1(\cmd_gen_inst|generating~q ),
	.ctl_reset_n(reset_reg_4),
	.read_req(read_req),
	.write_req(write_req),
	.bank_addr_0(\cmd_gen_inst|bank_addr[0]~0_combout ),
	.bank_addr_2(\cmd_gen_inst|bank_addr[2]~1_combout ),
	.bank_addr_1(\cmd_gen_inst|bank_addr[1]~2_combout ),
	.size_1(\cmd_gen_inst|size[1]~0_combout ),
	.size_0(\cmd_gen_inst|size[0]~1_combout ),
	.row_addr_12(\cmd_gen_inst|row_addr[12]~0_combout ),
	.row_addr_13(\cmd_gen_inst|row_addr[13]~1_combout ),
	.row_addr_11(\cmd_gen_inst|row_addr[11]~2_combout ),
	.row_addr_9(\cmd_gen_inst|row_addr[9]~3_combout ),
	.row_addr_10(\cmd_gen_inst|row_addr[10]~4_combout ),
	.row_addr_8(\cmd_gen_inst|row_addr[8]~5_combout ),
	.row_addr_6(\cmd_gen_inst|row_addr[6]~6_combout ),
	.row_addr_7(\cmd_gen_inst|row_addr[7]~7_combout ),
	.row_addr_2(\cmd_gen_inst|row_addr[2]~8_combout ),
	.row_addr_0(\cmd_gen_inst|row_addr[0]~9_combout ),
	.row_addr_1(\cmd_gen_inst|row_addr[1]~10_combout ),
	.row_addr_5(\cmd_gen_inst|row_addr[5]~11_combout ),
	.row_addr_3(\cmd_gen_inst|row_addr[3]~12_combout ),
	.row_addr_4(\cmd_gen_inst|row_addr[4]~13_combout ),
	.col_addr_2(\cmd_gen_inst|col_addr[2]~0_combout ),
	.col_addr_3(\cmd_gen_inst|col_addr[3]~1_combout ),
	.col_addr_4(\cmd_gen_inst|col_addr[4]~2_combout ),
	.col_addr_5(\cmd_gen_inst|col_addr[5]~3_combout ),
	.col_addr_6(\cmd_gen_inst|col_addr[6]~4_combout ),
	.col_addr_7(\cmd_gen_inst|col_addr[7]~5_combout ),
	.col_addr_8(\cmd_gen_inst|col_addr[8]~6_combout ),
	.col_addr_9(\cmd_gen_inst|col_addr[9]~7_combout ),
	.GND_port(GND_port),
	.local_size_1(local_size_1),
	.local_address_0(local_address_0),
	.local_size_0(local_size_0),
	.local_size_6(local_size_6),
	.local_size_5(local_size_5),
	.local_size_4(local_size_4),
	.local_size_2(local_size_2),
	.local_size_3(local_size_3),
	.local_read_req1(local_read_req),
	.local_write_req1(local_write_req),
	.local_burstbegin(local_burstbegin),
	.local_address_8(local_address_8),
	.local_address_10(local_address_10),
	.local_address_9(local_address_9),
	.local_address_23(local_address_23),
	.local_address_24(local_address_24),
	.local_address_22(local_address_22),
	.local_address_20(local_address_20),
	.local_address_21(local_address_21),
	.local_address_19(local_address_19),
	.local_address_17(local_address_17),
	.local_address_18(local_address_18),
	.local_address_13(local_address_13),
	.local_address_11(local_address_11),
	.local_address_12(local_address_12),
	.local_address_16(local_address_16),
	.local_address_14(local_address_14),
	.local_address_15(local_address_15),
	.local_address_1(local_address_1),
	.local_address_2(local_address_2),
	.local_address_3(local_address_3),
	.local_address_4(local_address_4),
	.local_address_5(local_address_5),
	.local_address_7(local_address_7),
	.local_address_6(local_address_6));

ddr3_int_alt_ddrx_wdata_fifo wdata_fifo_inst(
	.clk_0(clk_0),
	.q_b_132(q_b_132),
	.q_b_140(q_b_140),
	.q_b_128(q_b_128),
	.q_b_136(q_b_136),
	.q_b_133(q_b_133),
	.q_b_141(q_b_141),
	.q_b_129(q_b_129),
	.q_b_137(q_b_137),
	.q_b_134(q_b_134),
	.q_b_142(q_b_142),
	.q_b_130(q_b_130),
	.q_b_138(q_b_138),
	.q_b_135(q_b_135),
	.q_b_143(q_b_143),
	.q_b_131(q_b_131),
	.q_b_139(q_b_139),
	.q_b_96(q_b_96),
	.q_b_32(q_b_32),
	.q_b_64(q_b_64),
	.q_b_0(q_b_0),
	.q_b_97(q_b_97),
	.q_b_33(q_b_33),
	.q_b_65(q_b_65),
	.q_b_1(q_b_1),
	.q_b_98(q_b_98),
	.q_b_34(q_b_34),
	.q_b_66(q_b_66),
	.q_b_2(q_b_2),
	.q_b_99(q_b_99),
	.q_b_35(q_b_35),
	.q_b_67(q_b_67),
	.q_b_3(q_b_3),
	.q_b_100(q_b_100),
	.q_b_36(q_b_36),
	.q_b_68(q_b_68),
	.q_b_4(q_b_4),
	.q_b_101(q_b_101),
	.q_b_37(q_b_37),
	.q_b_69(q_b_69),
	.q_b_5(q_b_5),
	.q_b_102(q_b_102),
	.q_b_38(q_b_38),
	.q_b_70(q_b_70),
	.q_b_6(q_b_6),
	.q_b_103(q_b_103),
	.q_b_39(q_b_39),
	.q_b_71(q_b_71),
	.q_b_7(q_b_7),
	.q_b_104(q_b_104),
	.q_b_40(q_b_40),
	.q_b_72(q_b_72),
	.q_b_8(q_b_8),
	.q_b_105(q_b_105),
	.q_b_41(q_b_41),
	.q_b_73(q_b_73),
	.q_b_9(q_b_9),
	.q_b_106(q_b_106),
	.q_b_42(q_b_42),
	.q_b_74(q_b_74),
	.q_b_10(q_b_10),
	.q_b_107(q_b_107),
	.q_b_43(q_b_43),
	.q_b_75(q_b_75),
	.q_b_11(q_b_11),
	.q_b_108(q_b_108),
	.q_b_44(q_b_44),
	.q_b_76(q_b_76),
	.q_b_12(q_b_12),
	.q_b_109(q_b_109),
	.q_b_45(q_b_45),
	.q_b_77(q_b_77),
	.q_b_13(q_b_13),
	.q_b_110(q_b_110),
	.q_b_46(q_b_46),
	.q_b_78(q_b_78),
	.q_b_14(q_b_14),
	.q_b_111(q_b_111),
	.q_b_47(q_b_47),
	.q_b_79(q_b_79),
	.q_b_15(q_b_15),
	.q_b_112(q_b_112),
	.q_b_48(q_b_48),
	.q_b_80(q_b_80),
	.q_b_16(q_b_16),
	.q_b_113(q_b_113),
	.q_b_49(q_b_49),
	.q_b_81(q_b_81),
	.q_b_17(q_b_17),
	.q_b_114(q_b_114),
	.q_b_50(q_b_50),
	.q_b_82(q_b_82),
	.q_b_18(q_b_18),
	.q_b_115(q_b_115),
	.q_b_51(q_b_51),
	.q_b_83(q_b_83),
	.q_b_19(q_b_19),
	.q_b_116(q_b_116),
	.q_b_52(q_b_52),
	.q_b_84(q_b_84),
	.q_b_20(q_b_20),
	.q_b_117(q_b_117),
	.q_b_53(q_b_53),
	.q_b_85(q_b_85),
	.q_b_21(q_b_21),
	.q_b_118(q_b_118),
	.q_b_54(q_b_54),
	.q_b_86(q_b_86),
	.q_b_22(q_b_22),
	.q_b_119(q_b_119),
	.q_b_55(q_b_55),
	.q_b_87(q_b_87),
	.q_b_23(q_b_23),
	.q_b_120(q_b_120),
	.q_b_56(q_b_56),
	.q_b_88(q_b_88),
	.q_b_24(q_b_24),
	.q_b_121(q_b_121),
	.q_b_57(q_b_57),
	.q_b_89(q_b_89),
	.q_b_25(q_b_25),
	.q_b_122(q_b_122),
	.q_b_58(q_b_58),
	.q_b_90(q_b_90),
	.q_b_26(q_b_26),
	.q_b_123(q_b_123),
	.q_b_59(q_b_59),
	.q_b_91(q_b_91),
	.q_b_27(q_b_27),
	.q_b_124(q_b_124),
	.q_b_60(q_b_60),
	.q_b_92(q_b_92),
	.q_b_28(q_b_28),
	.q_b_125(q_b_125),
	.q_b_61(q_b_61),
	.q_b_93(q_b_93),
	.q_b_29(q_b_29),
	.q_b_126(q_b_126),
	.q_b_62(q_b_62),
	.q_b_94(q_b_94),
	.q_b_30(q_b_30),
	.q_b_127(q_b_127),
	.q_b_63(q_b_63),
	.q_b_95(q_b_95),
	.q_b_31(q_b_31),
	.dffe_af(\wdata_fifo_inst|wdata_fifo|auto_generated|dffe_af~q ),
	.ready_out(ready_out),
	.avalon_write_req(avalon_write_req),
	.ecc_wdata_fifo_read(ecc_wdata_fifo_read),
	.reset_reg_3(reset_reg_3),
	.local_write_req(local_write_req),
	.local_be_4(local_be_4),
	.local_be_12(local_be_12),
	.local_be_0(local_be_0),
	.local_be_8(local_be_8),
	.local_be_5(local_be_5),
	.local_be_13(local_be_13),
	.local_be_1(local_be_1),
	.local_be_9(local_be_9),
	.local_be_6(local_be_6),
	.local_be_14(local_be_14),
	.local_be_2(local_be_2),
	.local_be_10(local_be_10),
	.local_be_7(local_be_7),
	.local_be_15(local_be_15),
	.local_be_3(local_be_3),
	.local_be_11(local_be_11),
	.local_wdata_96(local_wdata_96),
	.local_wdata_32(local_wdata_32),
	.local_wdata_64(local_wdata_64),
	.local_wdata_0(local_wdata_0),
	.local_wdata_97(local_wdata_97),
	.local_wdata_33(local_wdata_33),
	.local_wdata_65(local_wdata_65),
	.local_wdata_1(local_wdata_1),
	.local_wdata_98(local_wdata_98),
	.local_wdata_34(local_wdata_34),
	.local_wdata_66(local_wdata_66),
	.local_wdata_2(local_wdata_2),
	.local_wdata_99(local_wdata_99),
	.local_wdata_35(local_wdata_35),
	.local_wdata_67(local_wdata_67),
	.local_wdata_3(local_wdata_3),
	.local_wdata_100(local_wdata_100),
	.local_wdata_36(local_wdata_36),
	.local_wdata_68(local_wdata_68),
	.local_wdata_4(local_wdata_4),
	.local_wdata_101(local_wdata_101),
	.local_wdata_37(local_wdata_37),
	.local_wdata_69(local_wdata_69),
	.local_wdata_5(local_wdata_5),
	.local_wdata_102(local_wdata_102),
	.local_wdata_38(local_wdata_38),
	.local_wdata_70(local_wdata_70),
	.local_wdata_6(local_wdata_6),
	.local_wdata_103(local_wdata_103),
	.local_wdata_39(local_wdata_39),
	.local_wdata_71(local_wdata_71),
	.local_wdata_7(local_wdata_7),
	.local_wdata_104(local_wdata_104),
	.local_wdata_40(local_wdata_40),
	.local_wdata_72(local_wdata_72),
	.local_wdata_8(local_wdata_8),
	.local_wdata_105(local_wdata_105),
	.local_wdata_41(local_wdata_41),
	.local_wdata_73(local_wdata_73),
	.local_wdata_9(local_wdata_9),
	.local_wdata_106(local_wdata_106),
	.local_wdata_42(local_wdata_42),
	.local_wdata_74(local_wdata_74),
	.local_wdata_10(local_wdata_10),
	.local_wdata_107(local_wdata_107),
	.local_wdata_43(local_wdata_43),
	.local_wdata_75(local_wdata_75),
	.local_wdata_11(local_wdata_11),
	.local_wdata_108(local_wdata_108),
	.local_wdata_44(local_wdata_44),
	.local_wdata_76(local_wdata_76),
	.local_wdata_12(local_wdata_12),
	.local_wdata_109(local_wdata_109),
	.local_wdata_45(local_wdata_45),
	.local_wdata_77(local_wdata_77),
	.local_wdata_13(local_wdata_13),
	.local_wdata_110(local_wdata_110),
	.local_wdata_46(local_wdata_46),
	.local_wdata_78(local_wdata_78),
	.local_wdata_14(local_wdata_14),
	.local_wdata_111(local_wdata_111),
	.local_wdata_47(local_wdata_47),
	.local_wdata_79(local_wdata_79),
	.local_wdata_15(local_wdata_15),
	.local_wdata_112(local_wdata_112),
	.local_wdata_48(local_wdata_48),
	.local_wdata_80(local_wdata_80),
	.local_wdata_16(local_wdata_16),
	.local_wdata_113(local_wdata_113),
	.local_wdata_49(local_wdata_49),
	.local_wdata_81(local_wdata_81),
	.local_wdata_17(local_wdata_17),
	.local_wdata_114(local_wdata_114),
	.local_wdata_50(local_wdata_50),
	.local_wdata_82(local_wdata_82),
	.local_wdata_18(local_wdata_18),
	.local_wdata_115(local_wdata_115),
	.local_wdata_51(local_wdata_51),
	.local_wdata_83(local_wdata_83),
	.local_wdata_19(local_wdata_19),
	.local_wdata_116(local_wdata_116),
	.local_wdata_52(local_wdata_52),
	.local_wdata_84(local_wdata_84),
	.local_wdata_20(local_wdata_20),
	.local_wdata_117(local_wdata_117),
	.local_wdata_53(local_wdata_53),
	.local_wdata_85(local_wdata_85),
	.local_wdata_21(local_wdata_21),
	.local_wdata_118(local_wdata_118),
	.local_wdata_54(local_wdata_54),
	.local_wdata_86(local_wdata_86),
	.local_wdata_22(local_wdata_22),
	.local_wdata_119(local_wdata_119),
	.local_wdata_55(local_wdata_55),
	.local_wdata_87(local_wdata_87),
	.local_wdata_23(local_wdata_23),
	.local_wdata_120(local_wdata_120),
	.local_wdata_56(local_wdata_56),
	.local_wdata_88(local_wdata_88),
	.local_wdata_24(local_wdata_24),
	.local_wdata_121(local_wdata_121),
	.local_wdata_57(local_wdata_57),
	.local_wdata_89(local_wdata_89),
	.local_wdata_25(local_wdata_25),
	.local_wdata_122(local_wdata_122),
	.local_wdata_58(local_wdata_58),
	.local_wdata_90(local_wdata_90),
	.local_wdata_26(local_wdata_26),
	.local_wdata_123(local_wdata_123),
	.local_wdata_59(local_wdata_59),
	.local_wdata_91(local_wdata_91),
	.local_wdata_27(local_wdata_27),
	.local_wdata_124(local_wdata_124),
	.local_wdata_60(local_wdata_60),
	.local_wdata_92(local_wdata_92),
	.local_wdata_28(local_wdata_28),
	.local_wdata_125(local_wdata_125),
	.local_wdata_61(local_wdata_61),
	.local_wdata_93(local_wdata_93),
	.local_wdata_29(local_wdata_29),
	.local_wdata_126(local_wdata_126),
	.local_wdata_62(local_wdata_62),
	.local_wdata_94(local_wdata_94),
	.local_wdata_30(local_wdata_30),
	.local_wdata_127(local_wdata_127),
	.local_wdata_63(local_wdata_63),
	.local_wdata_95(local_wdata_95),
	.local_wdata_31(local_wdata_31));

dffeas prolong_burstbegin(
	.clk(clk_0),
	.d(\prolong_burstbegin~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\prolong_burstbegin~q ),
	.prn(vcc));
defparam prolong_burstbegin.is_wysiwyg = "true";
defparam prolong_burstbegin.power_up = "low";

arriaii_lcell_comb \prolong_burstbegin~0 (
	.dataa(!ready_out),
	.datab(!local_write_req),
	.datac(!local_burstbegin),
	.datad(!\prolong_burstbegin~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\prolong_burstbegin~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \prolong_burstbegin~0 .extended_lut = "off";
defparam \prolong_burstbegin~0 .lut_mask = 64'h02EE02EE02EE02EE;
defparam \prolong_burstbegin~0 .shared_arith = "off";

arriaii_lcell_comb local_init_done(
	.dataa(!ctl_init_fail),
	.datab(!ctl_init_success),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(local_init_done1),
	.sumout(),
	.cout(),
	.shareout());
defparam local_init_done.extended_lut = "off";
defparam local_init_done.lut_mask = 64'h2222222222222222;
defparam local_init_done.shared_arith = "off";

arriaii_lcell_comb \internal_ready~0 (
	.dataa(!pipefull_7),
	.datab(!\gate_ready_in_reset~q ),
	.datac(!\wdata_fifo_inst|wdata_fifo|auto_generated|dffe_af~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(internal_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \internal_ready~0 .extended_lut = "off";
defparam \internal_ready~0 .lut_mask = 64'h2020202020202020;
defparam \internal_ready~0 .shared_arith = "off";

dffeas gate_ready_in_reset(
	.clk(clk_0),
	.d(vcc),
	.asdata(vcc),
	.clrn(ctl_reset_n[4]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\gate_ready_in_reset~q ),
	.prn(vcc));
defparam gate_ready_in_reset.is_wysiwyg = "true";
defparam gate_ready_in_reset.power_up = "low";

endmodule

module ddr3_int_alt_ddrx_avalon_if (
	hold_ready,
	pipefull_7,
	gate_ready_in_reset,
	dffe_af,
	avalon_read_req1,
	avalon_write_req1,
	local_read_req,
	local_write_req)/* synthesis synthesis_greybox=0 */;
input 	hold_ready;
input 	pipefull_7;
input 	gate_ready_in_reset;
input 	dffe_af;
output 	avalon_read_req1;
output 	avalon_write_req1;
input 	local_read_req;
input 	local_write_req;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



arriaii_lcell_comb avalon_read_req(
	.dataa(!hold_ready),
	.datab(!pipefull_7),
	.datac(!gate_ready_in_reset),
	.datad(!dffe_af),
	.datae(!local_read_req),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(avalon_read_req1),
	.sumout(),
	.cout(),
	.shareout());
defparam avalon_read_req.extended_lut = "off";
defparam avalon_read_req.lut_mask = 64'h0000080000000800;
defparam avalon_read_req.shared_arith = "off";

arriaii_lcell_comb avalon_write_req(
	.dataa(!hold_ready),
	.datab(!pipefull_7),
	.datac(!gate_ready_in_reset),
	.datad(!dffe_af),
	.datae(!local_write_req),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(avalon_write_req1),
	.sumout(),
	.cout(),
	.shareout());
defparam avalon_write_req.extended_lut = "off";
defparam avalon_write_req.lut_mask = 64'h0000080000000800;
defparam avalon_write_req.shared_arith = "off";

endmodule

module ddr3_int_alt_ddrx_cmd_gen (
	ctl_clk,
	buf_bank_addr_0,
	buf_bank_addr_2,
	buf_bank_addr_1,
	buf_col_addr_3,
	buf_col_addr_4,
	buf_col_addr_5,
	buf_col_addr_6,
	buf_col_addr_7,
	buf_col_addr_9,
	buf_col_addr_8,
	buf_row_addr_12,
	buf_row_addr_13,
	buf_row_addr_11,
	buf_row_addr_9,
	buf_row_addr_10,
	buf_row_addr_8,
	buf_row_addr_6,
	buf_row_addr_7,
	buf_row_addr_2,
	buf_row_addr_0,
	buf_row_addr_1,
	buf_row_addr_5,
	buf_row_addr_3,
	buf_row_addr_4,
	hold_ready1,
	pipefull_7,
	gate_ready_in_reset,
	dffe_af,
	ready_out1,
	internal_ready,
	local_read_req,
	local_write_req,
	prolong_burstbegin,
	generating1,
	ctl_reset_n,
	read_req,
	write_req,
	bank_addr_0,
	bank_addr_2,
	bank_addr_1,
	size_1,
	size_0,
	row_addr_12,
	row_addr_13,
	row_addr_11,
	row_addr_9,
	row_addr_10,
	row_addr_8,
	row_addr_6,
	row_addr_7,
	row_addr_2,
	row_addr_0,
	row_addr_1,
	row_addr_5,
	row_addr_3,
	row_addr_4,
	col_addr_2,
	col_addr_3,
	col_addr_4,
	col_addr_5,
	col_addr_6,
	col_addr_7,
	col_addr_8,
	col_addr_9,
	GND_port,
	local_size_1,
	local_address_0,
	local_size_0,
	local_size_6,
	local_size_5,
	local_size_4,
	local_size_2,
	local_size_3,
	local_read_req1,
	local_write_req1,
	local_burstbegin,
	local_address_8,
	local_address_10,
	local_address_9,
	local_address_23,
	local_address_24,
	local_address_22,
	local_address_20,
	local_address_21,
	local_address_19,
	local_address_17,
	local_address_18,
	local_address_13,
	local_address_11,
	local_address_12,
	local_address_16,
	local_address_14,
	local_address_15,
	local_address_1,
	local_address_2,
	local_address_3,
	local_address_4,
	local_address_5,
	local_address_7,
	local_address_6)/* synthesis synthesis_greybox=0 */;
input 	ctl_clk;
output 	buf_bank_addr_0;
output 	buf_bank_addr_2;
output 	buf_bank_addr_1;
output 	buf_col_addr_3;
output 	buf_col_addr_4;
output 	buf_col_addr_5;
output 	buf_col_addr_6;
output 	buf_col_addr_7;
output 	buf_col_addr_9;
output 	buf_col_addr_8;
output 	buf_row_addr_12;
output 	buf_row_addr_13;
output 	buf_row_addr_11;
output 	buf_row_addr_9;
output 	buf_row_addr_10;
output 	buf_row_addr_8;
output 	buf_row_addr_6;
output 	buf_row_addr_7;
output 	buf_row_addr_2;
output 	buf_row_addr_0;
output 	buf_row_addr_1;
output 	buf_row_addr_5;
output 	buf_row_addr_3;
output 	buf_row_addr_4;
output 	hold_ready1;
input 	pipefull_7;
input 	gate_ready_in_reset;
input 	dffe_af;
output 	ready_out1;
input 	internal_ready;
input 	local_read_req;
input 	local_write_req;
input 	prolong_burstbegin;
output 	generating1;
input 	ctl_reset_n;
output 	read_req;
output 	write_req;
output 	bank_addr_0;
output 	bank_addr_2;
output 	bank_addr_1;
output 	size_1;
output 	size_0;
output 	row_addr_12;
output 	row_addr_13;
output 	row_addr_11;
output 	row_addr_9;
output 	row_addr_10;
output 	row_addr_8;
output 	row_addr_6;
output 	row_addr_7;
output 	row_addr_2;
output 	row_addr_0;
output 	row_addr_1;
output 	row_addr_5;
output 	row_addr_3;
output 	row_addr_4;
output 	col_addr_2;
output 	col_addr_3;
output 	col_addr_4;
output 	col_addr_5;
output 	col_addr_6;
output 	col_addr_7;
output 	col_addr_8;
output 	col_addr_9;
input 	GND_port;
input 	local_size_1;
input 	local_address_0;
input 	local_size_0;
input 	local_size_6;
input 	local_size_5;
input 	local_size_4;
input 	local_size_2;
input 	local_size_3;
input 	local_read_req1;
input 	local_write_req1;
input 	local_burstbegin;
input 	local_address_8;
input 	local_address_10;
input 	local_address_9;
input 	local_address_23;
input 	local_address_24;
input 	local_address_22;
input 	local_address_20;
input 	local_address_21;
input 	local_address_19;
input 	local_address_17;
input 	local_address_18;
input 	local_address_13;
input 	local_address_11;
input 	local_address_12;
input 	local_address_16;
input 	local_address_14;
input 	local_address_15;
input 	local_address_1;
input 	local_address_2;
input 	local_address_3;
input 	local_address_4;
input 	local_address_5;
input 	local_address_7;
input 	local_address_6;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \buf_bank_addr[0]~_wirecell_combout ;
wire \copy~0_combout ;
wire \buf_read_req~q ;
wire \LessThan8~0_combout ;
wire \require_gen~0_combout ;
wire \registered~q ;
wire \pass_write~0_combout ;
wire \pass_write~q ;
wire \write_req~0_combout ;
wire \buf_col_addr[4]~0_combout ;
wire \buf_bank_addr[1]~0_combout ;
wire \buf_bank_addr[1]~1_combout ;
wire \buf_bank_addr~2_combout ;
wire \buf_bank_addr~3_combout ;
wire \Add78~1_sumout ;
wire \buf_col_addr[4]~1_combout ;
wire \Add78~2 ;
wire \Add78~5_sumout ;
wire \Add78~6 ;
wire \Add78~9_sumout ;
wire \Add78~10 ;
wire \Add78~13_sumout ;
wire \Add78~14 ;
wire \Add78~17_sumout ;
wire \Add78~18 ;
wire \Add78~22 ;
wire \Add78~25_sumout ;
wire \Add78~21_sumout ;
wire \Add76~2 ;
wire \Add76~6 ;
wire \Add76~10 ;
wire \Add76~14 ;
wire \Add76~18 ;
wire \Add76~22 ;
wire \Add76~26 ;
wire \Add76~30 ;
wire \Add76~34 ;
wire \Add76~38 ;
wire \Add76~42 ;
wire \Add76~46 ;
wire \Add76~49_sumout ;
wire \buf_row_addr[0]~0_combout ;
wire \buf_row_addr[0]~1_combout ;
wire \buf_row_addr[0]~2_combout ;
wire \buf_row_addr[0]~3_combout ;
wire \buf_row_addr[0]~5_combout ;
wire \buf_row_addr[0]~4_combout ;
wire \Add76~50 ;
wire \Add76~53_sumout ;
wire \Add76~45_sumout ;
wire \Add76~37_sumout ;
wire \Add76~41_sumout ;
wire \Add76~33_sumout ;
wire \Add76~25_sumout ;
wire \Add76~29_sumout ;
wire \Add76~9_sumout ;
wire \Add76~1_sumout ;
wire \Add76~5_sumout ;
wire \Add76~21_sumout ;
wire \Add76~13_sumout ;
wire \Add76~17_sumout ;
wire \Add73~1_sumout ;
wire \buf_size[0]~q ;
wire \Add73~2 ;
wire \Add73~5_sumout ;
wire \buf_size[1]~_wirecell_combout ;
wire \Add73~6 ;
wire \Add73~10 ;
wire \Add73~14 ;
wire \Add73~17_sumout ;
wire \Add73~13_sumout ;
wire \Add74~1_combout ;
wire \buf_size[3]~q ;
wire \Add74~2_combout ;
wire \buf_size[4]~q ;
wire \Add73~18 ;
wire \Add73~22 ;
wire \Add73~25_sumout ;
wire \Add73~21_sumout ;
wire \Add74~4_combout ;
wire \buf_size[5]~q ;
wire \Add74~3_combout ;
wire \buf_size[6]~q ;
wire \buf_size[6]~0_combout ;
wire \buf_size[6]~1_combout ;
wire \buf_size[6]~2_combout ;
wire \buf_size[1]~q ;
wire \LessThan7~0_combout ;
wire \buf_write_req~q ;
wire \hold_ready~0_combout ;
wire \hold_ready~1_combout ;
wire \generating~0_combout ;
wire \Add73~9_sumout ;
wire \Add74~0_combout ;
wire \buf_size[2]~q ;
wire \LessThan9~0_combout ;


dffeas \buf_bank_addr[0] (
	.clk(ctl_clk),
	.d(local_address_8),
	.asdata(\buf_bank_addr[0]~_wirecell_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\copy~0_combout ),
	.ena(\buf_bank_addr[1]~1_combout ),
	.q(buf_bank_addr_0),
	.prn(vcc));
defparam \buf_bank_addr[0] .is_wysiwyg = "true";
defparam \buf_bank_addr[0] .power_up = "low";

dffeas \buf_bank_addr[2] (
	.clk(ctl_clk),
	.d(local_address_10),
	.asdata(\buf_bank_addr~2_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\copy~0_combout ),
	.ena(\buf_bank_addr[1]~1_combout ),
	.q(buf_bank_addr_2),
	.prn(vcc));
defparam \buf_bank_addr[2] .is_wysiwyg = "true";
defparam \buf_bank_addr[2] .power_up = "low";

dffeas \buf_bank_addr[1] (
	.clk(ctl_clk),
	.d(local_address_9),
	.asdata(\buf_bank_addr~3_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\copy~0_combout ),
	.ena(\buf_bank_addr[1]~1_combout ),
	.q(buf_bank_addr_1),
	.prn(vcc));
defparam \buf_bank_addr[1] .is_wysiwyg = "true";
defparam \buf_bank_addr[1] .power_up = "low";

dffeas \buf_col_addr[3] (
	.clk(ctl_clk),
	.d(local_address_1),
	.asdata(\Add78~1_sumout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\copy~0_combout ),
	.ena(\buf_col_addr[4]~1_combout ),
	.q(buf_col_addr_3),
	.prn(vcc));
defparam \buf_col_addr[3] .is_wysiwyg = "true";
defparam \buf_col_addr[3] .power_up = "low";

dffeas \buf_col_addr[4] (
	.clk(ctl_clk),
	.d(local_address_2),
	.asdata(\Add78~5_sumout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\copy~0_combout ),
	.ena(\buf_col_addr[4]~1_combout ),
	.q(buf_col_addr_4),
	.prn(vcc));
defparam \buf_col_addr[4] .is_wysiwyg = "true";
defparam \buf_col_addr[4] .power_up = "low";

dffeas \buf_col_addr[5] (
	.clk(ctl_clk),
	.d(local_address_3),
	.asdata(\Add78~9_sumout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\copy~0_combout ),
	.ena(\buf_col_addr[4]~1_combout ),
	.q(buf_col_addr_5),
	.prn(vcc));
defparam \buf_col_addr[5] .is_wysiwyg = "true";
defparam \buf_col_addr[5] .power_up = "low";

dffeas \buf_col_addr[6] (
	.clk(ctl_clk),
	.d(local_address_4),
	.asdata(\Add78~13_sumout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\copy~0_combout ),
	.ena(\buf_col_addr[4]~1_combout ),
	.q(buf_col_addr_6),
	.prn(vcc));
defparam \buf_col_addr[6] .is_wysiwyg = "true";
defparam \buf_col_addr[6] .power_up = "low";

dffeas \buf_col_addr[7] (
	.clk(ctl_clk),
	.d(local_address_5),
	.asdata(\Add78~17_sumout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\copy~0_combout ),
	.ena(\buf_col_addr[4]~1_combout ),
	.q(buf_col_addr_7),
	.prn(vcc));
defparam \buf_col_addr[7] .is_wysiwyg = "true";
defparam \buf_col_addr[7] .power_up = "low";

dffeas \buf_col_addr[9] (
	.clk(ctl_clk),
	.d(local_address_7),
	.asdata(\Add78~25_sumout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\copy~0_combout ),
	.ena(\buf_col_addr[4]~1_combout ),
	.q(buf_col_addr_9),
	.prn(vcc));
defparam \buf_col_addr[9] .is_wysiwyg = "true";
defparam \buf_col_addr[9] .power_up = "low";

dffeas \buf_col_addr[8] (
	.clk(ctl_clk),
	.d(local_address_6),
	.asdata(\Add78~21_sumout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\copy~0_combout ),
	.ena(\buf_col_addr[4]~1_combout ),
	.q(buf_col_addr_8),
	.prn(vcc));
defparam \buf_col_addr[8] .is_wysiwyg = "true";
defparam \buf_col_addr[8] .power_up = "low";

dffeas \buf_row_addr[12] (
	.clk(ctl_clk),
	.d(\Add76~49_sumout ),
	.asdata(local_address_23),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\buf_row_addr[0]~3_combout ),
	.sload(\copy~0_combout ),
	.ena(\buf_row_addr[0]~4_combout ),
	.q(buf_row_addr_12),
	.prn(vcc));
defparam \buf_row_addr[12] .is_wysiwyg = "true";
defparam \buf_row_addr[12] .power_up = "low";

dffeas \buf_row_addr[13] (
	.clk(ctl_clk),
	.d(\Add76~53_sumout ),
	.asdata(local_address_24),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\buf_row_addr[0]~3_combout ),
	.sload(\copy~0_combout ),
	.ena(\buf_row_addr[0]~4_combout ),
	.q(buf_row_addr_13),
	.prn(vcc));
defparam \buf_row_addr[13] .is_wysiwyg = "true";
defparam \buf_row_addr[13] .power_up = "low";

dffeas \buf_row_addr[11] (
	.clk(ctl_clk),
	.d(\Add76~45_sumout ),
	.asdata(local_address_22),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\buf_row_addr[0]~3_combout ),
	.sload(\copy~0_combout ),
	.ena(\buf_row_addr[0]~4_combout ),
	.q(buf_row_addr_11),
	.prn(vcc));
defparam \buf_row_addr[11] .is_wysiwyg = "true";
defparam \buf_row_addr[11] .power_up = "low";

dffeas \buf_row_addr[9] (
	.clk(ctl_clk),
	.d(\Add76~37_sumout ),
	.asdata(local_address_20),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\buf_row_addr[0]~3_combout ),
	.sload(\copy~0_combout ),
	.ena(\buf_row_addr[0]~4_combout ),
	.q(buf_row_addr_9),
	.prn(vcc));
defparam \buf_row_addr[9] .is_wysiwyg = "true";
defparam \buf_row_addr[9] .power_up = "low";

dffeas \buf_row_addr[10] (
	.clk(ctl_clk),
	.d(\Add76~41_sumout ),
	.asdata(local_address_21),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\buf_row_addr[0]~3_combout ),
	.sload(\copy~0_combout ),
	.ena(\buf_row_addr[0]~4_combout ),
	.q(buf_row_addr_10),
	.prn(vcc));
defparam \buf_row_addr[10] .is_wysiwyg = "true";
defparam \buf_row_addr[10] .power_up = "low";

dffeas \buf_row_addr[8] (
	.clk(ctl_clk),
	.d(\Add76~33_sumout ),
	.asdata(local_address_19),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\buf_row_addr[0]~3_combout ),
	.sload(\copy~0_combout ),
	.ena(\buf_row_addr[0]~4_combout ),
	.q(buf_row_addr_8),
	.prn(vcc));
defparam \buf_row_addr[8] .is_wysiwyg = "true";
defparam \buf_row_addr[8] .power_up = "low";

dffeas \buf_row_addr[6] (
	.clk(ctl_clk),
	.d(\Add76~25_sumout ),
	.asdata(local_address_17),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\buf_row_addr[0]~3_combout ),
	.sload(\copy~0_combout ),
	.ena(\buf_row_addr[0]~4_combout ),
	.q(buf_row_addr_6),
	.prn(vcc));
defparam \buf_row_addr[6] .is_wysiwyg = "true";
defparam \buf_row_addr[6] .power_up = "low";

dffeas \buf_row_addr[7] (
	.clk(ctl_clk),
	.d(\Add76~29_sumout ),
	.asdata(local_address_18),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\buf_row_addr[0]~3_combout ),
	.sload(\copy~0_combout ),
	.ena(\buf_row_addr[0]~4_combout ),
	.q(buf_row_addr_7),
	.prn(vcc));
defparam \buf_row_addr[7] .is_wysiwyg = "true";
defparam \buf_row_addr[7] .power_up = "low";

dffeas \buf_row_addr[2] (
	.clk(ctl_clk),
	.d(\Add76~9_sumout ),
	.asdata(local_address_13),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\buf_row_addr[0]~3_combout ),
	.sload(\copy~0_combout ),
	.ena(\buf_row_addr[0]~4_combout ),
	.q(buf_row_addr_2),
	.prn(vcc));
defparam \buf_row_addr[2] .is_wysiwyg = "true";
defparam \buf_row_addr[2] .power_up = "low";

dffeas \buf_row_addr[0] (
	.clk(ctl_clk),
	.d(\Add76~1_sumout ),
	.asdata(local_address_11),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\buf_row_addr[0]~3_combout ),
	.sload(\copy~0_combout ),
	.ena(\buf_row_addr[0]~4_combout ),
	.q(buf_row_addr_0),
	.prn(vcc));
defparam \buf_row_addr[0] .is_wysiwyg = "true";
defparam \buf_row_addr[0] .power_up = "low";

dffeas \buf_row_addr[1] (
	.clk(ctl_clk),
	.d(\Add76~5_sumout ),
	.asdata(local_address_12),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\buf_row_addr[0]~3_combout ),
	.sload(\copy~0_combout ),
	.ena(\buf_row_addr[0]~4_combout ),
	.q(buf_row_addr_1),
	.prn(vcc));
defparam \buf_row_addr[1] .is_wysiwyg = "true";
defparam \buf_row_addr[1] .power_up = "low";

dffeas \buf_row_addr[5] (
	.clk(ctl_clk),
	.d(\Add76~21_sumout ),
	.asdata(local_address_16),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\buf_row_addr[0]~3_combout ),
	.sload(\copy~0_combout ),
	.ena(\buf_row_addr[0]~4_combout ),
	.q(buf_row_addr_5),
	.prn(vcc));
defparam \buf_row_addr[5] .is_wysiwyg = "true";
defparam \buf_row_addr[5] .power_up = "low";

dffeas \buf_row_addr[3] (
	.clk(ctl_clk),
	.d(\Add76~13_sumout ),
	.asdata(local_address_14),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\buf_row_addr[0]~3_combout ),
	.sload(\copy~0_combout ),
	.ena(\buf_row_addr[0]~4_combout ),
	.q(buf_row_addr_3),
	.prn(vcc));
defparam \buf_row_addr[3] .is_wysiwyg = "true";
defparam \buf_row_addr[3] .power_up = "low";

dffeas \buf_row_addr[4] (
	.clk(ctl_clk),
	.d(\Add76~17_sumout ),
	.asdata(local_address_15),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\buf_row_addr[0]~3_combout ),
	.sload(\copy~0_combout ),
	.ena(\buf_row_addr[0]~4_combout ),
	.q(buf_row_addr_4),
	.prn(vcc));
defparam \buf_row_addr[4] .is_wysiwyg = "true";
defparam \buf_row_addr[4] .power_up = "low";

dffeas hold_ready(
	.clk(ctl_clk),
	.d(\hold_ready~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(hold_ready1),
	.prn(vcc));
defparam hold_ready.is_wysiwyg = "true";
defparam hold_ready.power_up = "low";

arriaii_lcell_comb ready_out(
	.dataa(!hold_ready1),
	.datab(!pipefull_7),
	.datac(!gate_ready_in_reset),
	.datad(!dffe_af),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ready_out1),
	.sumout(),
	.cout(),
	.shareout());
defparam ready_out.extended_lut = "off";
defparam ready_out.lut_mask = 64'h0800080008000800;
defparam ready_out.shared_arith = "off";

dffeas generating(
	.clk(ctl_clk),
	.d(\generating~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(generating1),
	.prn(vcc));
defparam generating.is_wysiwyg = "true";
defparam generating.power_up = "low";

arriaii_lcell_comb \read_req~0 (
	.dataa(!hold_ready1),
	.datab(!internal_ready),
	.datac(!local_read_req1),
	.datad(!\buf_read_req~q ),
	.datae(!generating1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read_req),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_req~0 .extended_lut = "off";
defparam \read_req~0 .lut_mask = 64'h0202003302020033;
defparam \read_req~0 .shared_arith = "off";

arriaii_lcell_comb \write_req~1 (
	.dataa(!internal_ready),
	.datab(!local_write_req),
	.datac(!local_burstbegin),
	.datad(!prolong_burstbegin),
	.datae(!generating1),
	.dataf(!\write_req~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write_req),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_req~1 .extended_lut = "off";
defparam \write_req~1 .lut_mask = 64'h0333000003335555;
defparam \write_req~1 .shared_arith = "off";

arriaii_lcell_comb \bank_addr[0]~0 (
	.dataa(!generating1),
	.datab(!buf_bank_addr_0),
	.datac(!local_address_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(bank_addr_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \bank_addr[0]~0 .extended_lut = "off";
defparam \bank_addr[0]~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \bank_addr[0]~0 .shared_arith = "off";

arriaii_lcell_comb \bank_addr[2]~1 (
	.dataa(!generating1),
	.datab(!buf_bank_addr_2),
	.datac(!local_address_10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(bank_addr_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \bank_addr[2]~1 .extended_lut = "off";
defparam \bank_addr[2]~1 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \bank_addr[2]~1 .shared_arith = "off";

arriaii_lcell_comb \bank_addr[1]~2 (
	.dataa(!generating1),
	.datab(!buf_bank_addr_1),
	.datac(!local_address_9),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(bank_addr_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \bank_addr[1]~2 .extended_lut = "off";
defparam \bank_addr[1]~2 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \bank_addr[1]~2 .shared_arith = "off";

arriaii_lcell_comb \size[1]~0 (
	.dataa(!local_size_1),
	.datab(!local_address_0),
	.datac(!\LessThan8~0_combout ),
	.datad(!generating1),
	.datae(!\LessThan9~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(size_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \size[1]~0 .extended_lut = "off";
defparam \size[1]~0 .lut_mask = 64'hC4FFC400C4FFC400;
defparam \size[1]~0 .shared_arith = "off";

arriaii_lcell_comb \size[0]~1 (
	.dataa(!local_size_1),
	.datab(!local_address_0),
	.datac(!\LessThan8~0_combout ),
	.datad(!generating1),
	.datae(!\LessThan9~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(size_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \size[0]~1 .extended_lut = "off";
defparam \size[0]~1 .lut_mask = 64'h3B003BFF3B003BFF;
defparam \size[0]~1 .shared_arith = "off";

arriaii_lcell_comb \row_addr[12]~0 (
	.dataa(!generating1),
	.datab(!buf_row_addr_12),
	.datac(!local_address_23),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(row_addr_12),
	.sumout(),
	.cout(),
	.shareout());
defparam \row_addr[12]~0 .extended_lut = "off";
defparam \row_addr[12]~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \row_addr[12]~0 .shared_arith = "off";

arriaii_lcell_comb \row_addr[13]~1 (
	.dataa(!generating1),
	.datab(!buf_row_addr_13),
	.datac(!local_address_24),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(row_addr_13),
	.sumout(),
	.cout(),
	.shareout());
defparam \row_addr[13]~1 .extended_lut = "off";
defparam \row_addr[13]~1 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \row_addr[13]~1 .shared_arith = "off";

arriaii_lcell_comb \row_addr[11]~2 (
	.dataa(!generating1),
	.datab(!buf_row_addr_11),
	.datac(!local_address_22),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(row_addr_11),
	.sumout(),
	.cout(),
	.shareout());
defparam \row_addr[11]~2 .extended_lut = "off";
defparam \row_addr[11]~2 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \row_addr[11]~2 .shared_arith = "off";

arriaii_lcell_comb \row_addr[9]~3 (
	.dataa(!generating1),
	.datab(!buf_row_addr_9),
	.datac(!local_address_20),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(row_addr_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \row_addr[9]~3 .extended_lut = "off";
defparam \row_addr[9]~3 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \row_addr[9]~3 .shared_arith = "off";

arriaii_lcell_comb \row_addr[10]~4 (
	.dataa(!generating1),
	.datab(!buf_row_addr_10),
	.datac(!local_address_21),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(row_addr_10),
	.sumout(),
	.cout(),
	.shareout());
defparam \row_addr[10]~4 .extended_lut = "off";
defparam \row_addr[10]~4 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \row_addr[10]~4 .shared_arith = "off";

arriaii_lcell_comb \row_addr[8]~5 (
	.dataa(!generating1),
	.datab(!buf_row_addr_8),
	.datac(!local_address_19),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(row_addr_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \row_addr[8]~5 .extended_lut = "off";
defparam \row_addr[8]~5 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \row_addr[8]~5 .shared_arith = "off";

arriaii_lcell_comb \row_addr[6]~6 (
	.dataa(!generating1),
	.datab(!buf_row_addr_6),
	.datac(!local_address_17),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(row_addr_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \row_addr[6]~6 .extended_lut = "off";
defparam \row_addr[6]~6 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \row_addr[6]~6 .shared_arith = "off";

arriaii_lcell_comb \row_addr[7]~7 (
	.dataa(!generating1),
	.datab(!buf_row_addr_7),
	.datac(!local_address_18),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(row_addr_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \row_addr[7]~7 .extended_lut = "off";
defparam \row_addr[7]~7 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \row_addr[7]~7 .shared_arith = "off";

arriaii_lcell_comb \row_addr[2]~8 (
	.dataa(!generating1),
	.datab(!buf_row_addr_2),
	.datac(!local_address_13),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(row_addr_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \row_addr[2]~8 .extended_lut = "off";
defparam \row_addr[2]~8 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \row_addr[2]~8 .shared_arith = "off";

arriaii_lcell_comb \row_addr[0]~9 (
	.dataa(!generating1),
	.datab(!buf_row_addr_0),
	.datac(!local_address_11),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(row_addr_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \row_addr[0]~9 .extended_lut = "off";
defparam \row_addr[0]~9 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \row_addr[0]~9 .shared_arith = "off";

arriaii_lcell_comb \row_addr[1]~10 (
	.dataa(!generating1),
	.datab(!buf_row_addr_1),
	.datac(!local_address_12),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(row_addr_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \row_addr[1]~10 .extended_lut = "off";
defparam \row_addr[1]~10 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \row_addr[1]~10 .shared_arith = "off";

arriaii_lcell_comb \row_addr[5]~11 (
	.dataa(!generating1),
	.datab(!buf_row_addr_5),
	.datac(!local_address_16),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(row_addr_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \row_addr[5]~11 .extended_lut = "off";
defparam \row_addr[5]~11 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \row_addr[5]~11 .shared_arith = "off";

arriaii_lcell_comb \row_addr[3]~12 (
	.dataa(!generating1),
	.datab(!buf_row_addr_3),
	.datac(!local_address_14),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(row_addr_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \row_addr[3]~12 .extended_lut = "off";
defparam \row_addr[3]~12 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \row_addr[3]~12 .shared_arith = "off";

arriaii_lcell_comb \row_addr[4]~13 (
	.dataa(!generating1),
	.datab(!buf_row_addr_4),
	.datac(!local_address_15),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(row_addr_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \row_addr[4]~13 .extended_lut = "off";
defparam \row_addr[4]~13 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \row_addr[4]~13 .shared_arith = "off";

arriaii_lcell_comb \col_addr[2]~0 (
	.dataa(!local_address_0),
	.datab(!generating1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(col_addr_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \col_addr[2]~0 .extended_lut = "off";
defparam \col_addr[2]~0 .lut_mask = 64'h4444444444444444;
defparam \col_addr[2]~0 .shared_arith = "off";

arriaii_lcell_comb \col_addr[3]~1 (
	.dataa(!generating1),
	.datab(!buf_col_addr_3),
	.datac(!local_address_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(col_addr_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \col_addr[3]~1 .extended_lut = "off";
defparam \col_addr[3]~1 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \col_addr[3]~1 .shared_arith = "off";

arriaii_lcell_comb \col_addr[4]~2 (
	.dataa(!generating1),
	.datab(!buf_col_addr_4),
	.datac(!local_address_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(col_addr_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \col_addr[4]~2 .extended_lut = "off";
defparam \col_addr[4]~2 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \col_addr[4]~2 .shared_arith = "off";

arriaii_lcell_comb \col_addr[5]~3 (
	.dataa(!generating1),
	.datab(!buf_col_addr_5),
	.datac(!local_address_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(col_addr_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \col_addr[5]~3 .extended_lut = "off";
defparam \col_addr[5]~3 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \col_addr[5]~3 .shared_arith = "off";

arriaii_lcell_comb \col_addr[6]~4 (
	.dataa(!generating1),
	.datab(!buf_col_addr_6),
	.datac(!local_address_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(col_addr_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \col_addr[6]~4 .extended_lut = "off";
defparam \col_addr[6]~4 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \col_addr[6]~4 .shared_arith = "off";

arriaii_lcell_comb \col_addr[7]~5 (
	.dataa(!generating1),
	.datab(!buf_col_addr_7),
	.datac(!local_address_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(col_addr_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \col_addr[7]~5 .extended_lut = "off";
defparam \col_addr[7]~5 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \col_addr[7]~5 .shared_arith = "off";

arriaii_lcell_comb \col_addr[8]~6 (
	.dataa(!generating1),
	.datab(!buf_col_addr_8),
	.datac(!local_address_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(col_addr_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \col_addr[8]~6 .extended_lut = "off";
defparam \col_addr[8]~6 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \col_addr[8]~6 .shared_arith = "off";

arriaii_lcell_comb \col_addr[9]~7 (
	.dataa(!generating1),
	.datab(!buf_col_addr_9),
	.datac(!local_address_7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(col_addr_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \col_addr[9]~7 .extended_lut = "off";
defparam \col_addr[9]~7 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \col_addr[9]~7 .shared_arith = "off";

arriaii_lcell_comb \buf_bank_addr[0]~_wirecell (
	.dataa(!buf_bank_addr_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\buf_bank_addr[0]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \buf_bank_addr[0]~_wirecell .extended_lut = "off";
defparam \buf_bank_addr[0]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \buf_bank_addr[0]~_wirecell .shared_arith = "off";

arriaii_lcell_comb \copy~0 (
	.dataa(!internal_ready),
	.datab(!local_read_req),
	.datac(!local_write_req),
	.datad(!local_burstbegin),
	.datae(!prolong_burstbegin),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\copy~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \copy~0 .extended_lut = "off";
defparam \copy~0 .lut_mask = 64'h1115151511151515;
defparam \copy~0 .shared_arith = "off";

dffeas buf_read_req(
	.clk(ctl_clk),
	.d(local_read_req),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\copy~0_combout ),
	.q(\buf_read_req~q ),
	.prn(vcc));
defparam buf_read_req.is_wysiwyg = "true";
defparam buf_read_req.power_up = "low";

arriaii_lcell_comb \LessThan8~0 (
	.dataa(!local_size_6),
	.datab(!local_size_5),
	.datac(!local_size_4),
	.datad(!local_size_2),
	.datae(!local_size_3),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan8~0 .extended_lut = "off";
defparam \LessThan8~0 .lut_mask = 64'h8000000080000000;
defparam \LessThan8~0 .shared_arith = "off";

arriaii_lcell_comb \require_gen~0 (
	.dataa(!local_size_1),
	.datab(!local_address_0),
	.datac(!local_size_0),
	.datad(!\LessThan8~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\require_gen~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \require_gen~0 .extended_lut = "off";
defparam \require_gen~0 .lut_mask = 64'hFF15FF15FF15FF15;
defparam \require_gen~0 .shared_arith = "off";

dffeas registered(
	.clk(ctl_clk),
	.d(\require_gen~0_combout ),
	.asdata(GND_port),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\copy~0_combout ),
	.ena(vcc),
	.q(\registered~q ),
	.prn(vcc));
defparam registered.is_wysiwyg = "true";
defparam registered.power_up = "low";

arriaii_lcell_comb \pass_write~0 (
	.dataa(!local_address_0),
	.datab(!\require_gen~0_combout ),
	.datac(!local_write_req),
	.datad(!\copy~0_combout ),
	.datae(!\pass_write~q ),
	.dataf(!\registered~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pass_write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pass_write~0 .extended_lut = "off";
defparam \pass_write~0 .lut_mask = 64'h0F1DF0D10011FFDD;
defparam \pass_write~0 .shared_arith = "off";

dffeas pass_write(
	.clk(ctl_clk),
	.d(\pass_write~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pass_write~q ),
	.prn(vcc));
defparam pass_write.is_wysiwyg = "true";
defparam pass_write.power_up = "low";

arriaii_lcell_comb \write_req~0 (
	.dataa(!hold_ready1),
	.datab(!local_write_req1),
	.datac(!\pass_write~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write_req~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_req~0 .extended_lut = "off";
defparam \write_req~0 .lut_mask = 64'h0202020202020202;
defparam \write_req~0 .shared_arith = "off";

arriaii_lcell_comb \buf_col_addr[4]~0 (
	.dataa(!internal_ready),
	.datab(!\buf_read_req~q ),
	.datac(!generating1),
	.datad(!\write_req~0_combout ),
	.datae(!\registered~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\buf_col_addr[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \buf_col_addr[4]~0 .extended_lut = "off";
defparam \buf_col_addr[4]~0 .lut_mask = 64'hFEFA0000FEFA0000;
defparam \buf_col_addr[4]~0 .shared_arith = "off";

arriaii_lcell_comb \buf_bank_addr[1]~0 (
	.dataa(!buf_col_addr_6),
	.datab(!buf_col_addr_7),
	.datac(!buf_col_addr_9),
	.datad(!buf_col_addr_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\buf_bank_addr[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \buf_bank_addr[1]~0 .extended_lut = "off";
defparam \buf_bank_addr[1]~0 .lut_mask = 64'h0001000100010001;
defparam \buf_bank_addr[1]~0 .shared_arith = "off";

arriaii_lcell_comb \buf_bank_addr[1]~1 (
	.dataa(!\copy~0_combout ),
	.datab(!\buf_col_addr[4]~0_combout ),
	.datac(!buf_col_addr_3),
	.datad(!buf_col_addr_4),
	.datae(!buf_col_addr_5),
	.dataf(!\buf_bank_addr[1]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\buf_bank_addr[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \buf_bank_addr[1]~1 .extended_lut = "off";
defparam \buf_bank_addr[1]~1 .lut_mask = 64'h555555555555555D;
defparam \buf_bank_addr[1]~1 .shared_arith = "off";

arriaii_lcell_comb \buf_bank_addr~2 (
	.dataa(!buf_bank_addr_0),
	.datab(!buf_bank_addr_2),
	.datac(!buf_bank_addr_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\buf_bank_addr~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \buf_bank_addr~2 .extended_lut = "off";
defparam \buf_bank_addr~2 .lut_mask = 64'h3636363636363636;
defparam \buf_bank_addr~2 .shared_arith = "off";

arriaii_lcell_comb \buf_bank_addr~3 (
	.dataa(!buf_bank_addr_0),
	.datab(!buf_bank_addr_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\buf_bank_addr~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \buf_bank_addr~3 .extended_lut = "off";
defparam \buf_bank_addr~3 .lut_mask = 64'h6666666666666666;
defparam \buf_bank_addr~3 .shared_arith = "off";

arriaii_lcell_comb \Add78~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!buf_col_addr_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add78~1_sumout ),
	.cout(\Add78~2 ),
	.shareout());
defparam \Add78~1 .extended_lut = "off";
defparam \Add78~1 .lut_mask = 64'h00000000000000FF;
defparam \Add78~1 .shared_arith = "off";

arriaii_lcell_comb \buf_col_addr[4]~1 (
	.dataa(!\copy~0_combout ),
	.datab(!\buf_col_addr[4]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\buf_col_addr[4]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \buf_col_addr[4]~1 .extended_lut = "off";
defparam \buf_col_addr[4]~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \buf_col_addr[4]~1 .shared_arith = "off";

arriaii_lcell_comb \Add78~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!buf_col_addr_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add78~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add78~5_sumout ),
	.cout(\Add78~6 ),
	.shareout());
defparam \Add78~5 .extended_lut = "off";
defparam \Add78~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add78~5 .shared_arith = "off";

arriaii_lcell_comb \Add78~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!buf_col_addr_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add78~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add78~9_sumout ),
	.cout(\Add78~10 ),
	.shareout());
defparam \Add78~9 .extended_lut = "off";
defparam \Add78~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add78~9 .shared_arith = "off";

arriaii_lcell_comb \Add78~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!buf_col_addr_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add78~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add78~13_sumout ),
	.cout(\Add78~14 ),
	.shareout());
defparam \Add78~13 .extended_lut = "off";
defparam \Add78~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add78~13 .shared_arith = "off";

arriaii_lcell_comb \Add78~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!buf_col_addr_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add78~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add78~17_sumout ),
	.cout(\Add78~18 ),
	.shareout());
defparam \Add78~17 .extended_lut = "off";
defparam \Add78~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add78~17 .shared_arith = "off";

arriaii_lcell_comb \Add78~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!buf_col_addr_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add78~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add78~21_sumout ),
	.cout(\Add78~22 ),
	.shareout());
defparam \Add78~21 .extended_lut = "off";
defparam \Add78~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add78~21 .shared_arith = "off";

arriaii_lcell_comb \Add78~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!buf_col_addr_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add78~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add78~25_sumout ),
	.cout(),
	.shareout());
defparam \Add78~25 .extended_lut = "off";
defparam \Add78~25 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add78~25 .shared_arith = "off";

arriaii_lcell_comb \Add76~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!buf_row_addr_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add76~1_sumout ),
	.cout(\Add76~2 ),
	.shareout());
defparam \Add76~1 .extended_lut = "off";
defparam \Add76~1 .lut_mask = 64'h00000000000000FF;
defparam \Add76~1 .shared_arith = "off";

arriaii_lcell_comb \Add76~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!buf_row_addr_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add76~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add76~5_sumout ),
	.cout(\Add76~6 ),
	.shareout());
defparam \Add76~5 .extended_lut = "off";
defparam \Add76~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add76~5 .shared_arith = "off";

arriaii_lcell_comb \Add76~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!buf_row_addr_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add76~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add76~9_sumout ),
	.cout(\Add76~10 ),
	.shareout());
defparam \Add76~9 .extended_lut = "off";
defparam \Add76~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add76~9 .shared_arith = "off";

arriaii_lcell_comb \Add76~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!buf_row_addr_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add76~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add76~13_sumout ),
	.cout(\Add76~14 ),
	.shareout());
defparam \Add76~13 .extended_lut = "off";
defparam \Add76~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add76~13 .shared_arith = "off";

arriaii_lcell_comb \Add76~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!buf_row_addr_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add76~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add76~17_sumout ),
	.cout(\Add76~18 ),
	.shareout());
defparam \Add76~17 .extended_lut = "off";
defparam \Add76~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add76~17 .shared_arith = "off";

arriaii_lcell_comb \Add76~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!buf_row_addr_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add76~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add76~21_sumout ),
	.cout(\Add76~22 ),
	.shareout());
defparam \Add76~21 .extended_lut = "off";
defparam \Add76~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add76~21 .shared_arith = "off";

arriaii_lcell_comb \Add76~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!buf_row_addr_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add76~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add76~25_sumout ),
	.cout(\Add76~26 ),
	.shareout());
defparam \Add76~25 .extended_lut = "off";
defparam \Add76~25 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add76~25 .shared_arith = "off";

arriaii_lcell_comb \Add76~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!buf_row_addr_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add76~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add76~29_sumout ),
	.cout(\Add76~30 ),
	.shareout());
defparam \Add76~29 .extended_lut = "off";
defparam \Add76~29 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add76~29 .shared_arith = "off";

arriaii_lcell_comb \Add76~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!buf_row_addr_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add76~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add76~33_sumout ),
	.cout(\Add76~34 ),
	.shareout());
defparam \Add76~33 .extended_lut = "off";
defparam \Add76~33 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add76~33 .shared_arith = "off";

arriaii_lcell_comb \Add76~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!buf_row_addr_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add76~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add76~37_sumout ),
	.cout(\Add76~38 ),
	.shareout());
defparam \Add76~37 .extended_lut = "off";
defparam \Add76~37 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add76~37 .shared_arith = "off";

arriaii_lcell_comb \Add76~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!buf_row_addr_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add76~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add76~41_sumout ),
	.cout(\Add76~42 ),
	.shareout());
defparam \Add76~41 .extended_lut = "off";
defparam \Add76~41 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add76~41 .shared_arith = "off";

arriaii_lcell_comb \Add76~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!buf_row_addr_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add76~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add76~45_sumout ),
	.cout(\Add76~46 ),
	.shareout());
defparam \Add76~45 .extended_lut = "off";
defparam \Add76~45 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add76~45 .shared_arith = "off";

arriaii_lcell_comb \Add76~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!buf_row_addr_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add76~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add76~49_sumout ),
	.cout(\Add76~50 ),
	.shareout());
defparam \Add76~49 .extended_lut = "off";
defparam \Add76~49 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add76~49 .shared_arith = "off";

arriaii_lcell_comb \buf_row_addr[0]~0 (
	.dataa(!buf_row_addr_12),
	.datab(!buf_row_addr_13),
	.datac(!buf_row_addr_2),
	.datad(!buf_row_addr_0),
	.datae(!buf_row_addr_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\buf_row_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \buf_row_addr[0]~0 .extended_lut = "off";
defparam \buf_row_addr[0]~0 .lut_mask = 64'h0000000100000001;
defparam \buf_row_addr[0]~0 .shared_arith = "off";

arriaii_lcell_comb \buf_row_addr[0]~1 (
	.dataa(!buf_row_addr_9),
	.datab(!buf_row_addr_10),
	.datac(!buf_row_addr_8),
	.datad(!buf_row_addr_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\buf_row_addr[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \buf_row_addr[0]~1 .extended_lut = "off";
defparam \buf_row_addr[0]~1 .lut_mask = 64'h0001000100010001;
defparam \buf_row_addr[0]~1 .shared_arith = "off";

arriaii_lcell_comb \buf_row_addr[0]~2 (
	.dataa(!buf_row_addr_11),
	.datab(!buf_row_addr_6),
	.datac(!buf_row_addr_5),
	.datad(!\buf_row_addr[0]~0_combout ),
	.datae(!\buf_row_addr[0]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\buf_row_addr[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \buf_row_addr[0]~2 .extended_lut = "off";
defparam \buf_row_addr[0]~2 .lut_mask = 64'h0000000100000001;
defparam \buf_row_addr[0]~2 .shared_arith = "off";

arriaii_lcell_comb \buf_row_addr[0]~3 (
	.dataa(!\copy~0_combout ),
	.datab(!buf_row_addr_3),
	.datac(!buf_row_addr_4),
	.datad(!\buf_row_addr[0]~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\buf_row_addr[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \buf_row_addr[0]~3 .extended_lut = "off";
defparam \buf_row_addr[0]~3 .lut_mask = 64'h0002000200020002;
defparam \buf_row_addr[0]~3 .shared_arith = "off";

arriaii_lcell_comb \buf_row_addr[0]~5 (
	.dataa(!buf_bank_addr_1),
	.datab(!buf_col_addr_3),
	.datac(!buf_col_addr_4),
	.datad(!buf_col_addr_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\buf_row_addr[0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \buf_row_addr[0]~5 .extended_lut = "off";
defparam \buf_row_addr[0]~5 .lut_mask = 64'h0001000100010001;
defparam \buf_row_addr[0]~5 .shared_arith = "off";

arriaii_lcell_comb \buf_row_addr[0]~4 (
	.dataa(!\copy~0_combout ),
	.datab(!buf_bank_addr_0),
	.datac(!buf_bank_addr_2),
	.datad(!\buf_col_addr[4]~0_combout ),
	.datae(!\buf_bank_addr[1]~0_combout ),
	.dataf(!\buf_row_addr[0]~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\buf_row_addr[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \buf_row_addr[0]~4 .extended_lut = "off";
defparam \buf_row_addr[0]~4 .lut_mask = 64'h5555555555555755;
defparam \buf_row_addr[0]~4 .shared_arith = "off";

arriaii_lcell_comb \Add76~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!buf_row_addr_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add76~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add76~53_sumout ),
	.cout(),
	.shareout());
defparam \Add76~53 .extended_lut = "off";
defparam \Add76~53 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add76~53 .shared_arith = "off";

arriaii_lcell_comb \Add73~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!local_size_0),
	.datae(gnd),
	.dataf(!local_address_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add73~1_sumout ),
	.cout(\Add73~2 ),
	.shareout());
defparam \Add73~1 .extended_lut = "off";
defparam \Add73~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add73~1 .shared_arith = "off";

dffeas \buf_size[0] (
	.clk(ctl_clk),
	.d(\Add73~1_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\copy~0_combout ),
	.q(\buf_size[0]~q ),
	.prn(vcc));
defparam \buf_size[0] .is_wysiwyg = "true";
defparam \buf_size[0] .power_up = "low";

arriaii_lcell_comb \Add73~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!local_size_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add73~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add73~5_sumout ),
	.cout(\Add73~6 ),
	.shareout());
defparam \Add73~5 .extended_lut = "off";
defparam \Add73~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add73~5 .shared_arith = "off";

arriaii_lcell_comb \buf_size[1]~_wirecell (
	.dataa(!\buf_size[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\buf_size[1]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \buf_size[1]~_wirecell .extended_lut = "off";
defparam \buf_size[1]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \buf_size[1]~_wirecell .shared_arith = "off";

arriaii_lcell_comb \Add73~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!local_size_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add73~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add73~9_sumout ),
	.cout(\Add73~10 ),
	.shareout());
defparam \Add73~9 .extended_lut = "off";
defparam \Add73~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add73~9 .shared_arith = "off";

arriaii_lcell_comb \Add73~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!local_size_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add73~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add73~13_sumout ),
	.cout(\Add73~14 ),
	.shareout());
defparam \Add73~13 .extended_lut = "off";
defparam \Add73~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add73~13 .shared_arith = "off";

arriaii_lcell_comb \Add73~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!local_size_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add73~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add73~17_sumout ),
	.cout(\Add73~18 ),
	.shareout());
defparam \Add73~17 .extended_lut = "off";
defparam \Add73~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add73~17 .shared_arith = "off";

arriaii_lcell_comb \Add74~1 (
	.dataa(!\buf_size[2]~q ),
	.datab(!\buf_size[1]~q ),
	.datac(!\buf_size[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add74~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add74~1 .extended_lut = "off";
defparam \Add74~1 .lut_mask = 64'h8787878787878787;
defparam \Add74~1 .shared_arith = "off";

dffeas \buf_size[3] (
	.clk(ctl_clk),
	.d(\Add73~13_sumout ),
	.asdata(\Add74~1_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\copy~0_combout ),
	.ena(\buf_size[6]~2_combout ),
	.q(\buf_size[3]~q ),
	.prn(vcc));
defparam \buf_size[3] .is_wysiwyg = "true";
defparam \buf_size[3] .power_up = "low";

arriaii_lcell_comb \Add74~2 (
	.dataa(!\buf_size[2]~q ),
	.datab(!\buf_size[1]~q ),
	.datac(!\buf_size[3]~q ),
	.datad(!\buf_size[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add74~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add74~2 .extended_lut = "off";
defparam \Add74~2 .lut_mask = 64'h807F807F807F807F;
defparam \Add74~2 .shared_arith = "off";

dffeas \buf_size[4] (
	.clk(ctl_clk),
	.d(\Add73~17_sumout ),
	.asdata(\Add74~2_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\copy~0_combout ),
	.ena(\buf_size[6]~2_combout ),
	.q(\buf_size[4]~q ),
	.prn(vcc));
defparam \buf_size[4] .is_wysiwyg = "true";
defparam \buf_size[4] .power_up = "low";

arriaii_lcell_comb \Add73~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!local_size_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add73~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add73~21_sumout ),
	.cout(\Add73~22 ),
	.shareout());
defparam \Add73~21 .extended_lut = "off";
defparam \Add73~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add73~21 .shared_arith = "off";

arriaii_lcell_comb \Add73~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!local_size_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add73~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add73~25_sumout ),
	.cout(),
	.shareout());
defparam \Add73~25 .extended_lut = "off";
defparam \Add73~25 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add73~25 .shared_arith = "off";

arriaii_lcell_comb \Add74~4 (
	.dataa(!\buf_size[2]~q ),
	.datab(!\buf_size[1]~q ),
	.datac(!\buf_size[3]~q ),
	.datad(!\buf_size[4]~q ),
	.datae(!\buf_size[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add74~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add74~4 .extended_lut = "off";
defparam \Add74~4 .lut_mask = 64'h80007FFF80007FFF;
defparam \Add74~4 .shared_arith = "off";

dffeas \buf_size[5] (
	.clk(ctl_clk),
	.d(\Add73~21_sumout ),
	.asdata(\Add74~4_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\copy~0_combout ),
	.ena(\buf_size[6]~2_combout ),
	.q(\buf_size[5]~q ),
	.prn(vcc));
defparam \buf_size[5] .is_wysiwyg = "true";
defparam \buf_size[5] .power_up = "low";

arriaii_lcell_comb \Add74~3 (
	.dataa(!\buf_size[2]~q ),
	.datab(!\buf_size[1]~q ),
	.datac(!\buf_size[3]~q ),
	.datad(!\buf_size[4]~q ),
	.datae(!\buf_size[6]~q ),
	.dataf(!\buf_size[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add74~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add74~3 .extended_lut = "off";
defparam \Add74~3 .lut_mask = 64'h80007FFF0000FFFF;
defparam \Add74~3 .shared_arith = "off";

dffeas \buf_size[6] (
	.clk(ctl_clk),
	.d(\Add73~25_sumout ),
	.asdata(\Add74~3_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\copy~0_combout ),
	.ena(\buf_size[6]~2_combout ),
	.q(\buf_size[6]~q ),
	.prn(vcc));
defparam \buf_size[6] .is_wysiwyg = "true";
defparam \buf_size[6] .power_up = "low";

arriaii_lcell_comb \buf_size[6]~0 (
	.dataa(!\buf_size[3]~q ),
	.datab(!\buf_size[4]~q ),
	.datac(!\buf_size[6]~q ),
	.datad(!\buf_size[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\buf_size[6]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \buf_size[6]~0 .extended_lut = "off";
defparam \buf_size[6]~0 .lut_mask = 64'h8000800080008000;
defparam \buf_size[6]~0 .shared_arith = "off";

arriaii_lcell_comb \buf_size[6]~1 (
	.dataa(!\buf_size[2]~q ),
	.datab(!\buf_size[0]~q ),
	.datac(!\buf_size[1]~q ),
	.datad(!\buf_size[6]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\buf_size[6]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \buf_size[6]~1 .extended_lut = "off";
defparam \buf_size[6]~1 .lut_mask = 64'h00A800A800A800A8;
defparam \buf_size[6]~1 .shared_arith = "off";

arriaii_lcell_comb \buf_size[6]~2 (
	.dataa(!internal_ready),
	.datab(!\copy~0_combout ),
	.datac(!\buf_read_req~q ),
	.datad(!\write_req~0_combout ),
	.datae(!\buf_size[6]~1_combout ),
	.dataf(!\registered~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\buf_size[6]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \buf_size[6]~2 .extended_lut = "off";
defparam \buf_size[6]~2 .lut_mask = 64'h3777333333333333;
defparam \buf_size[6]~2 .shared_arith = "off";

dffeas \buf_size[1] (
	.clk(ctl_clk),
	.d(\Add73~5_sumout ),
	.asdata(\buf_size[1]~_wirecell_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\copy~0_combout ),
	.ena(\buf_size[6]~2_combout ),
	.q(\buf_size[1]~q ),
	.prn(vcc));
defparam \buf_size[1] .is_wysiwyg = "true";
defparam \buf_size[1] .power_up = "low";

arriaii_lcell_comb \LessThan7~0 (
	.dataa(!\buf_size[2]~q ),
	.datab(!\buf_size[0]~q ),
	.datac(!\buf_size[1]~q ),
	.datad(!\buf_size[6]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan7~0 .extended_lut = "off";
defparam \LessThan7~0 .lut_mask = 64'h00EA00EA00EA00EA;
defparam \LessThan7~0 .shared_arith = "off";

dffeas buf_write_req(
	.clk(ctl_clk),
	.d(local_write_req),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\copy~0_combout ),
	.q(\buf_write_req~q ),
	.prn(vcc));
defparam buf_write_req.is_wysiwyg = "true";
defparam buf_write_req.power_up = "low";

arriaii_lcell_comb \hold_ready~0 (
	.dataa(!hold_ready1),
	.datab(!internal_ready),
	.datac(!\buf_read_req~q ),
	.datad(!\buf_write_req~q ),
	.datae(!generating1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\hold_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \hold_ready~0 .extended_lut = "off";
defparam \hold_ready~0 .lut_mask = 64'h5500540055005400;
defparam \hold_ready~0 .shared_arith = "off";

arriaii_lcell_comb \hold_ready~1 (
	.dataa(!\require_gen~0_combout ),
	.datab(!\copy~0_combout ),
	.datac(!\buf_read_req~q ),
	.datad(!\LessThan7~0_combout ),
	.datae(!\hold_ready~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\hold_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \hold_ready~1 .extended_lut = "off";
defparam \hold_ready~1 .lut_mask = 64'h1F11FFFF1F11FFFF;
defparam \hold_ready~1 .shared_arith = "off";

arriaii_lcell_comb \generating~0 (
	.dataa(!internal_ready),
	.datab(!\buf_read_req~q ),
	.datac(!\LessThan7~0_combout ),
	.datad(!generating1),
	.datae(!\write_req~0_combout ),
	.dataf(!\registered~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\generating~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \generating~0 .extended_lut = "off";
defparam \generating~0 .lut_mask = 64'h00FE00FAFFFFFFFF;
defparam \generating~0 .shared_arith = "off";

arriaii_lcell_comb \Add74~0 (
	.dataa(!\buf_size[2]~q ),
	.datab(!\buf_size[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add74~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add74~0 .extended_lut = "off";
defparam \Add74~0 .lut_mask = 64'h9999999999999999;
defparam \Add74~0 .shared_arith = "off";

dffeas \buf_size[2] (
	.clk(ctl_clk),
	.d(\Add73~9_sumout ),
	.asdata(\Add74~0_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\copy~0_combout ),
	.ena(\buf_size[6]~2_combout ),
	.q(\buf_size[2]~q ),
	.prn(vcc));
defparam \buf_size[2] .is_wysiwyg = "true";
defparam \buf_size[2] .power_up = "low";

arriaii_lcell_comb \LessThan9~0 (
	.dataa(!\buf_size[2]~q ),
	.datab(!\buf_size[1]~q ),
	.datac(!\buf_size[3]~q ),
	.datad(!\buf_size[4]~q ),
	.datae(!\buf_size[6]~q ),
	.dataf(!\buf_size[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan9~0 .extended_lut = "off";
defparam \LessThan9~0 .lut_mask = 64'h2000000000000000;
defparam \LessThan9~0 .shared_arith = "off";

endmodule

module ddr3_int_alt_ddrx_cmd_queue (
	ctl_clk,
	pipe_10_0,
	pipe_12_0,
	pipe_11_0,
	pipe_32_0,
	pipe_12_2,
	pipe_12_3,
	pipe_12_1,
	pipe_10_2,
	pipe_10_3,
	pipe_10_1,
	pipe_11_2,
	pipe_11_3,
	pipe_11_1,
	pipe_29_0,
	pipe_28_0,
	pipe_33_0,
	pipe_12_4,
	pipe_11_4,
	pipe_10_4,
	buf_bank_addr_0,
	buf_bank_addr_2,
	buf_bank_addr_1,
	pipe_25_5,
	pipe_25_0,
	pipe_26_5,
	pipe_26_0,
	pipe_24_5,
	pipe_24_0,
	pipe_22_5,
	pipe_22_0,
	pipe_23_5,
	pipe_23_0,
	pipe_21_5,
	pipe_21_0,
	pipe_19_5,
	pipe_19_0,
	pipe_20_5,
	pipe_20_0,
	pipe_15_5,
	pipe_15_0,
	pipe_13_5,
	pipe_13_0,
	pipe_14_5,
	pipe_14_0,
	pipe_18_5,
	pipe_18_0,
	pipe_16_5,
	pipe_16_0,
	pipe_17_5,
	pipe_17_0,
	pipe_12_5,
	pipe_11_5,
	pipe_10_5,
	pipe_25_3,
	pipe_26_3,
	pipe_24_3,
	pipe_22_3,
	pipe_23_3,
	pipe_21_3,
	pipe_19_3,
	pipe_20_3,
	pipe_15_3,
	pipe_13_3,
	pipe_14_3,
	pipe_18_3,
	pipe_16_3,
	pipe_17_3,
	pipe_25_4,
	pipe_26_4,
	pipe_24_4,
	pipe_22_4,
	pipe_23_4,
	pipe_21_4,
	pipe_19_4,
	pipe_20_4,
	pipe_15_4,
	pipe_13_4,
	pipe_14_4,
	pipe_18_4,
	pipe_16_4,
	pipe_17_4,
	pipe_12_6,
	pipe_11_6,
	pipe_10_6,
	pipe_25_6,
	pipe_26_6,
	pipe_24_6,
	pipe_22_6,
	pipe_23_6,
	pipe_21_6,
	pipe_19_6,
	pipe_20_6,
	pipe_15_6,
	pipe_13_6,
	pipe_14_6,
	pipe_18_6,
	pipe_16_6,
	pipe_17_6,
	pipe_26_7,
	pipe_24_7,
	pipe_25_7,
	pipe_23_7,
	pipe_21_7,
	pipe_22_7,
	pipe_20_7,
	pipe_18_7,
	pipe_19_7,
	pipe_17_7,
	pipe_15_7,
	pipe_16_7,
	pipe_11_7,
	pipe_10_7,
	pipe_14_7,
	pipe_12_7,
	pipe_13_7,
	pipe_25_2,
	pipe_26_2,
	pipe_24_2,
	pipe_22_2,
	pipe_23_2,
	pipe_21_2,
	pipe_19_2,
	pipe_20_2,
	pipe_15_2,
	pipe_13_2,
	pipe_14_2,
	pipe_18_2,
	pipe_16_2,
	pipe_17_2,
	pipe_25_1,
	pipe_26_1,
	pipe_24_1,
	pipe_22_1,
	pipe_23_1,
	pipe_21_1,
	pipe_19_1,
	pipe_20_1,
	pipe_15_1,
	pipe_13_1,
	pipe_14_1,
	pipe_18_1,
	pipe_16_1,
	pipe_17_1,
	buf_col_addr_3,
	buf_col_addr_4,
	buf_col_addr_5,
	buf_col_addr_6,
	buf_col_addr_7,
	buf_col_addr_9,
	buf_col_addr_8,
	buf_row_addr_12,
	buf_row_addr_13,
	buf_row_addr_11,
	buf_row_addr_9,
	buf_row_addr_10,
	buf_row_addr_8,
	buf_row_addr_6,
	buf_row_addr_7,
	buf_row_addr_2,
	buf_row_addr_0,
	buf_row_addr_1,
	buf_row_addr_5,
	buf_row_addr_3,
	buf_row_addr_4,
	pipe_2_0,
	pipe_3_0,
	pipe_4_0,
	pipe_5_0,
	pipe_6_0,
	pipe_7_0,
	pipe_8_0,
	pipe_9_0,
	pipefull_7,
	generating,
	fetch,
	read_req,
	write_req,
	pipefull_6,
	ctl_reset_n,
	always38,
	pipefull_0,
	pipefull_5,
	pipefull_1,
	pipefull_4,
	pipefull_2,
	pipefull_3,
	bank_addr_0,
	bank_addr_2,
	bank_addr_1,
	size_1,
	size_0,
	row_addr_12,
	row_addr_13,
	row_addr_11,
	row_addr_9,
	row_addr_10,
	row_addr_8,
	row_addr_6,
	row_addr_7,
	row_addr_2,
	row_addr_0,
	row_addr_1,
	row_addr_5,
	row_addr_3,
	row_addr_4,
	col_addr_2,
	col_addr_3,
	col_addr_4,
	col_addr_5,
	col_addr_6,
	col_addr_7,
	col_addr_8,
	col_addr_9,
	local_address_0,
	local_address_8,
	local_address_10,
	local_address_9,
	local_address_23,
	local_address_24,
	local_address_22,
	local_address_20,
	local_address_21,
	local_address_19,
	local_address_17,
	local_address_18,
	local_address_13,
	local_address_11,
	local_address_12,
	local_address_16,
	local_address_14,
	local_address_15,
	local_address_1,
	local_address_2,
	local_address_3,
	local_address_4,
	local_address_5,
	local_address_7,
	local_address_6)/* synthesis synthesis_greybox=0 */;
input 	ctl_clk;
output 	pipe_10_0;
output 	pipe_12_0;
output 	pipe_11_0;
output 	pipe_32_0;
output 	pipe_12_2;
output 	pipe_12_3;
output 	pipe_12_1;
output 	pipe_10_2;
output 	pipe_10_3;
output 	pipe_10_1;
output 	pipe_11_2;
output 	pipe_11_3;
output 	pipe_11_1;
output 	pipe_29_0;
output 	pipe_28_0;
output 	pipe_33_0;
output 	pipe_12_4;
output 	pipe_11_4;
output 	pipe_10_4;
input 	buf_bank_addr_0;
input 	buf_bank_addr_2;
input 	buf_bank_addr_1;
output 	pipe_25_5;
output 	pipe_25_0;
output 	pipe_26_5;
output 	pipe_26_0;
output 	pipe_24_5;
output 	pipe_24_0;
output 	pipe_22_5;
output 	pipe_22_0;
output 	pipe_23_5;
output 	pipe_23_0;
output 	pipe_21_5;
output 	pipe_21_0;
output 	pipe_19_5;
output 	pipe_19_0;
output 	pipe_20_5;
output 	pipe_20_0;
output 	pipe_15_5;
output 	pipe_15_0;
output 	pipe_13_5;
output 	pipe_13_0;
output 	pipe_14_5;
output 	pipe_14_0;
output 	pipe_18_5;
output 	pipe_18_0;
output 	pipe_16_5;
output 	pipe_16_0;
output 	pipe_17_5;
output 	pipe_17_0;
output 	pipe_12_5;
output 	pipe_11_5;
output 	pipe_10_5;
output 	pipe_25_3;
output 	pipe_26_3;
output 	pipe_24_3;
output 	pipe_22_3;
output 	pipe_23_3;
output 	pipe_21_3;
output 	pipe_19_3;
output 	pipe_20_3;
output 	pipe_15_3;
output 	pipe_13_3;
output 	pipe_14_3;
output 	pipe_18_3;
output 	pipe_16_3;
output 	pipe_17_3;
output 	pipe_25_4;
output 	pipe_26_4;
output 	pipe_24_4;
output 	pipe_22_4;
output 	pipe_23_4;
output 	pipe_21_4;
output 	pipe_19_4;
output 	pipe_20_4;
output 	pipe_15_4;
output 	pipe_13_4;
output 	pipe_14_4;
output 	pipe_18_4;
output 	pipe_16_4;
output 	pipe_17_4;
output 	pipe_12_6;
output 	pipe_11_6;
output 	pipe_10_6;
output 	pipe_25_6;
output 	pipe_26_6;
output 	pipe_24_6;
output 	pipe_22_6;
output 	pipe_23_6;
output 	pipe_21_6;
output 	pipe_19_6;
output 	pipe_20_6;
output 	pipe_15_6;
output 	pipe_13_6;
output 	pipe_14_6;
output 	pipe_18_6;
output 	pipe_16_6;
output 	pipe_17_6;
output 	pipe_26_7;
output 	pipe_24_7;
output 	pipe_25_7;
output 	pipe_23_7;
output 	pipe_21_7;
output 	pipe_22_7;
output 	pipe_20_7;
output 	pipe_18_7;
output 	pipe_19_7;
output 	pipe_17_7;
output 	pipe_15_7;
output 	pipe_16_7;
output 	pipe_11_7;
output 	pipe_10_7;
output 	pipe_14_7;
output 	pipe_12_7;
output 	pipe_13_7;
output 	pipe_25_2;
output 	pipe_26_2;
output 	pipe_24_2;
output 	pipe_22_2;
output 	pipe_23_2;
output 	pipe_21_2;
output 	pipe_19_2;
output 	pipe_20_2;
output 	pipe_15_2;
output 	pipe_13_2;
output 	pipe_14_2;
output 	pipe_18_2;
output 	pipe_16_2;
output 	pipe_17_2;
output 	pipe_25_1;
output 	pipe_26_1;
output 	pipe_24_1;
output 	pipe_22_1;
output 	pipe_23_1;
output 	pipe_21_1;
output 	pipe_19_1;
output 	pipe_20_1;
output 	pipe_15_1;
output 	pipe_13_1;
output 	pipe_14_1;
output 	pipe_18_1;
output 	pipe_16_1;
output 	pipe_17_1;
input 	buf_col_addr_3;
input 	buf_col_addr_4;
input 	buf_col_addr_5;
input 	buf_col_addr_6;
input 	buf_col_addr_7;
input 	buf_col_addr_9;
input 	buf_col_addr_8;
input 	buf_row_addr_12;
input 	buf_row_addr_13;
input 	buf_row_addr_11;
input 	buf_row_addr_9;
input 	buf_row_addr_10;
input 	buf_row_addr_8;
input 	buf_row_addr_6;
input 	buf_row_addr_7;
input 	buf_row_addr_2;
input 	buf_row_addr_0;
input 	buf_row_addr_1;
input 	buf_row_addr_5;
input 	buf_row_addr_3;
input 	buf_row_addr_4;
output 	pipe_2_0;
output 	pipe_3_0;
output 	pipe_4_0;
output 	pipe_5_0;
output 	pipe_6_0;
output 	pipe_7_0;
output 	pipe_8_0;
output 	pipe_9_0;
output 	pipefull_7;
input 	generating;
input 	fetch;
input 	read_req;
input 	write_req;
output 	pipefull_6;
input 	ctl_reset_n;
input 	always38;
output 	pipefull_0;
output 	pipefull_5;
output 	pipefull_1;
output 	pipefull_4;
output 	pipefull_2;
output 	pipefull_3;
input 	bank_addr_0;
input 	bank_addr_2;
input 	bank_addr_1;
input 	size_1;
input 	size_0;
input 	row_addr_12;
input 	row_addr_13;
input 	row_addr_11;
input 	row_addr_9;
input 	row_addr_10;
input 	row_addr_8;
input 	row_addr_6;
input 	row_addr_7;
input 	row_addr_2;
input 	row_addr_0;
input 	row_addr_1;
input 	row_addr_5;
input 	row_addr_3;
input 	row_addr_4;
input 	col_addr_2;
input 	col_addr_3;
input 	col_addr_4;
input 	col_addr_5;
input 	col_addr_6;
input 	col_addr_7;
input 	col_addr_8;
input 	col_addr_9;
input 	local_address_0;
input 	local_address_8;
input 	local_address_10;
input 	local_address_9;
input 	local_address_23;
input 	local_address_24;
input 	local_address_22;
input 	local_address_20;
input 	local_address_21;
input 	local_address_19;
input 	local_address_17;
input 	local_address_18;
input 	local_address_13;
input 	local_address_11;
input 	local_address_12;
input 	local_address_16;
input 	local_address_14;
input 	local_address_15;
input 	local_address_1;
input 	local_address_2;
input 	local_address_3;
input 	local_address_4;
input 	local_address_5;
input 	local_address_7;
input 	local_address_6;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \pipe~0_combout ;
wire \pipe[0][5]~1_combout ;
wire \pipe~2_combout ;
wire \pipe~3_combout ;
wire \pipe~192_combout ;
wire \pipe[1][11]~7_combout ;
wire \pipe[7][32]~q ;
wire \pipe~180_combout ;
wire \pipe[6][32]~q ;
wire \pipe~168_combout ;
wire \pipe[5][32]~q ;
wire \pipe~156_combout ;
wire \pipe[4][32]~q ;
wire \pipe~151_combout ;
wire \pipe[3][32]~q ;
wire \pipe~146_combout ;
wire \pipe[2][32]~q ;
wire \pipe~21_combout ;
wire \pipe[1][32]~q ;
wire \pipe~4_combout ;
wire \pipe~5_combout ;
wire \pipe~6_combout ;
wire \pipe~8_combout ;
wire \pipe~9_combout ;
wire \pipe~10_combout ;
wire \pipe~11_combout ;
wire \pipe~12_combout ;
wire \pipe~13_combout ;
wire \pipe~14_combout ;
wire \pipe~194_combout ;
wire \pipe[7][29]~q ;
wire \pipe~182_combout ;
wire \pipe[6][29]~q ;
wire \pipe~170_combout ;
wire \pipe[5][29]~q ;
wire \pipe~158_combout ;
wire \pipe[4][29]~q ;
wire \pipe~153_combout ;
wire \pipe[3][29]~q ;
wire \pipe~148_combout ;
wire \pipe[2][29]~q ;
wire \pipe~143_combout ;
wire \pipe[1][29]~q ;
wire \pipe~15_combout ;
wire \pipe~195_combout ;
wire \pipe[7][28]~q ;
wire \pipe~183_combout ;
wire \pipe[6][28]~q ;
wire \pipe~171_combout ;
wire \pipe[5][28]~q ;
wire \pipe~159_combout ;
wire \pipe[4][28]~q ;
wire \pipe~154_combout ;
wire \pipe[3][28]~q ;
wire \pipe~149_combout ;
wire \pipe[2][28]~q ;
wire \pipe~144_combout ;
wire \pipe[1][28]~q ;
wire \pipe~16_combout ;
wire \pipe~196_combout ;
wire \pipe[7][33]~q ;
wire \pipe~184_combout ;
wire \pipe[6][33]~q ;
wire \pipe~172_combout ;
wire \pipe[5][33]~q ;
wire \pipe~160_combout ;
wire \pipe[4][33]~q ;
wire \pipe~155_combout ;
wire \pipe[3][33]~q ;
wire \pipe~150_combout ;
wire \pipe[2][33]~q ;
wire \pipe~145_combout ;
wire \pipe[1][33]~q ;
wire \pipe~17_combout ;
wire \pipe~18_combout ;
wire \pipe~19_combout ;
wire \pipe~20_combout ;
wire \pipe~22_combout ;
wire \pipe~23_combout ;
wire \pipe~24_combout ;
wire \pipe~25_combout ;
wire \pipe~26_combout ;
wire \pipe~27_combout ;
wire \pipe~28_combout ;
wire \pipe~29_combout ;
wire \pipe~30_combout ;
wire \pipe~31_combout ;
wire \pipe~32_combout ;
wire \pipe~33_combout ;
wire \pipe~34_combout ;
wire \pipe~35_combout ;
wire \pipe~36_combout ;
wire \pipe~37_combout ;
wire \pipe~38_combout ;
wire \pipe~39_combout ;
wire \pipe~40_combout ;
wire \pipe~41_combout ;
wire \pipe~42_combout ;
wire \pipe~43_combout ;
wire \pipe~44_combout ;
wire \pipe~45_combout ;
wire \pipe~46_combout ;
wire \pipe~47_combout ;
wire \pipe~48_combout ;
wire \pipe~49_combout ;
wire \pipe~50_combout ;
wire \pipe~51_combout ;
wire \pipe~52_combout ;
wire \pipe~53_combout ;
wire \pipe~54_combout ;
wire \pipe~55_combout ;
wire \pipe~56_combout ;
wire \pipe~57_combout ;
wire \pipe~58_combout ;
wire \pipe~59_combout ;
wire \pipe~60_combout ;
wire \pipe~61_combout ;
wire \pipe~62_combout ;
wire \pipe~63_combout ;
wire \pipe~64_combout ;
wire \pipe~65_combout ;
wire \pipe~66_combout ;
wire \pipe~67_combout ;
wire \pipe~68_combout ;
wire \pipe~69_combout ;
wire \pipe~70_combout ;
wire \pipe~71_combout ;
wire \pipe~72_combout ;
wire \pipe~73_combout ;
wire \pipe~74_combout ;
wire \pipe~75_combout ;
wire \pipe~76_combout ;
wire \pipe~77_combout ;
wire \pipe~78_combout ;
wire \pipe~79_combout ;
wire \pipe~80_combout ;
wire \pipe~81_combout ;
wire \pipe~82_combout ;
wire \pipe~83_combout ;
wire \pipe~84_combout ;
wire \pipe~85_combout ;
wire \pipe~86_combout ;
wire \pipe~87_combout ;
wire \pipe~88_combout ;
wire \pipe~89_combout ;
wire \pipe~90_combout ;
wire \pipe~91_combout ;
wire \pipe~92_combout ;
wire \pipe~93_combout ;
wire \pipe~94_combout ;
wire \pipe~95_combout ;
wire \pipe~96_combout ;
wire \pipe~97_combout ;
wire \pipe~98_combout ;
wire \pipe~99_combout ;
wire \pipe~100_combout ;
wire \pipe~101_combout ;
wire \pipe~102_combout ;
wire \pipe~103_combout ;
wire \pipe~104_combout ;
wire \pipe~105_combout ;
wire \pipe~106_combout ;
wire \pipe~107_combout ;
wire \pipe~108_combout ;
wire \pipe~109_combout ;
wire \pipe~110_combout ;
wire \pipe~111_combout ;
wire \pipe~112_combout ;
wire \pipe~113_combout ;
wire \pipe~114_combout ;
wire \pipe~115_combout ;
wire \pipe~116_combout ;
wire \pipe~117_combout ;
wire \pipe~118_combout ;
wire \pipe~119_combout ;
wire \pipe~120_combout ;
wire \pipe~121_combout ;
wire \pipe~122_combout ;
wire \pipe~123_combout ;
wire \pipe~124_combout ;
wire \pipe~125_combout ;
wire \pipe~126_combout ;
wire \pipe~127_combout ;
wire \pipe~128_combout ;
wire \pipe~129_combout ;
wire \pipe~130_combout ;
wire \pipe~131_combout ;
wire \pipe~132_combout ;
wire \pipe~133_combout ;
wire \pipe~134_combout ;
wire \pipe~135_combout ;
wire \pipe~136_combout ;
wire \pipe~137_combout ;
wire \pipe~138_combout ;
wire \pipe~139_combout ;
wire \pipe~140_combout ;
wire \pipe~141_combout ;
wire \pipe~142_combout ;
wire \pipe~212_combout ;
wire \pipe[7][2]~q ;
wire \pipe~204_combout ;
wire \pipe[6][2]~q ;
wire \pipe~193_combout ;
wire \pipe[5][2]~q ;
wire \pipe~181_combout ;
wire \pipe[4][2]~q ;
wire \pipe~169_combout ;
wire \pipe[3][2]~q ;
wire \pipe~157_combout ;
wire \pipe[2][2]~q ;
wire \pipe~152_combout ;
wire \pipe[1][2]~q ;
wire \pipe~147_combout ;
wire \pipe~227_combout ;
wire \pipe[7][3]~q ;
wire \pipe~220_combout ;
wire \pipe[6][3]~q ;
wire \pipe~213_combout ;
wire \pipe[5][3]~q ;
wire \pipe~205_combout ;
wire \pipe[4][3]~q ;
wire \pipe~197_combout ;
wire \pipe[3][3]~q ;
wire \pipe~185_combout ;
wire \pipe[2][3]~q ;
wire \pipe~173_combout ;
wire \pipe[1][3]~q ;
wire \pipe~161_combout ;
wire \pipe~228_combout ;
wire \pipe[7][4]~q ;
wire \pipe~221_combout ;
wire \pipe[6][4]~q ;
wire \pipe~214_combout ;
wire \pipe[5][4]~q ;
wire \pipe~206_combout ;
wire \pipe[4][4]~q ;
wire \pipe~198_combout ;
wire \pipe[3][4]~q ;
wire \pipe~186_combout ;
wire \pipe[2][4]~q ;
wire \pipe~174_combout ;
wire \pipe[1][4]~q ;
wire \pipe~162_combout ;
wire \pipe~229_combout ;
wire \pipe[7][5]~q ;
wire \pipe~222_combout ;
wire \pipe[6][5]~q ;
wire \pipe~215_combout ;
wire \pipe[5][5]~q ;
wire \pipe~207_combout ;
wire \pipe[4][5]~q ;
wire \pipe~199_combout ;
wire \pipe[3][5]~q ;
wire \pipe~187_combout ;
wire \pipe[2][5]~q ;
wire \pipe~175_combout ;
wire \pipe[1][5]~q ;
wire \pipe~163_combout ;
wire \pipe~230_combout ;
wire \pipe[7][6]~q ;
wire \pipe~223_combout ;
wire \pipe[6][6]~q ;
wire \pipe~216_combout ;
wire \pipe[5][6]~q ;
wire \pipe~208_combout ;
wire \pipe[4][6]~q ;
wire \pipe~200_combout ;
wire \pipe[3][6]~q ;
wire \pipe~188_combout ;
wire \pipe[2][6]~q ;
wire \pipe~176_combout ;
wire \pipe[1][6]~q ;
wire \pipe~164_combout ;
wire \pipe~231_combout ;
wire \pipe[7][7]~q ;
wire \pipe~224_combout ;
wire \pipe[6][7]~q ;
wire \pipe~217_combout ;
wire \pipe[5][7]~q ;
wire \pipe~209_combout ;
wire \pipe[4][7]~q ;
wire \pipe~201_combout ;
wire \pipe[3][7]~q ;
wire \pipe~189_combout ;
wire \pipe[2][7]~q ;
wire \pipe~177_combout ;
wire \pipe[1][7]~q ;
wire \pipe~165_combout ;
wire \pipe~232_combout ;
wire \pipe[7][8]~q ;
wire \pipe~225_combout ;
wire \pipe[6][8]~q ;
wire \pipe~218_combout ;
wire \pipe[5][8]~q ;
wire \pipe~210_combout ;
wire \pipe[4][8]~q ;
wire \pipe~202_combout ;
wire \pipe[3][8]~q ;
wire \pipe~190_combout ;
wire \pipe[2][8]~q ;
wire \pipe~178_combout ;
wire \pipe[1][8]~q ;
wire \pipe~166_combout ;
wire \pipe~233_combout ;
wire \pipe[7][9]~q ;
wire \pipe~226_combout ;
wire \pipe[6][9]~q ;
wire \pipe~219_combout ;
wire \pipe[5][9]~q ;
wire \pipe~211_combout ;
wire \pipe[4][9]~q ;
wire \pipe~203_combout ;
wire \pipe[3][9]~q ;
wire \pipe~191_combout ;
wire \pipe[2][9]~q ;
wire \pipe~179_combout ;
wire \pipe[1][9]~q ;
wire \pipe~167_combout ;
wire \pipefull~0_combout ;
wire \pipefull~1_combout ;
wire \pipefull~2_combout ;
wire \pipefull~3_combout ;
wire \pipefull~4_combout ;
wire \pipefull~5_combout ;
wire \pipefull~6_combout ;
wire \pipefull~7_combout ;


dffeas \pipe[0][10] (
	.clk(ctl_clk),
	.d(\pipe~0_combout ),
	.asdata(bank_addr_0),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[0][5]~1_combout ),
	.q(pipe_10_0),
	.prn(vcc));
defparam \pipe[0][10] .is_wysiwyg = "true";
defparam \pipe[0][10] .power_up = "low";

dffeas \pipe[0][12] (
	.clk(ctl_clk),
	.d(\pipe~2_combout ),
	.asdata(bank_addr_2),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[0][5]~1_combout ),
	.q(pipe_12_0),
	.prn(vcc));
defparam \pipe[0][12] .is_wysiwyg = "true";
defparam \pipe[0][12] .power_up = "low";

dffeas \pipe[0][11] (
	.clk(ctl_clk),
	.d(\pipe~3_combout ),
	.asdata(bank_addr_1),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[0][5]~1_combout ),
	.q(pipe_11_0),
	.prn(vcc));
defparam \pipe[0][11] .is_wysiwyg = "true";
defparam \pipe[0][11] .power_up = "low";

dffeas \pipe[0][32] (
	.clk(ctl_clk),
	.d(\pipe~4_combout ),
	.asdata(write_req),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[0][5]~1_combout ),
	.q(pipe_32_0),
	.prn(vcc));
defparam \pipe[0][32] .is_wysiwyg = "true";
defparam \pipe[0][32] .power_up = "low";

dffeas \pipe[2][12] (
	.clk(ctl_clk),
	.d(\pipe~5_combout ),
	.asdata(\pipe~6_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_12_2),
	.prn(vcc));
defparam \pipe[2][12] .is_wysiwyg = "true";
defparam \pipe[2][12] .power_up = "low";

dffeas \pipe[3][12] (
	.clk(ctl_clk),
	.d(\pipe~8_combout ),
	.asdata(\pipe~5_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_12_3),
	.prn(vcc));
defparam \pipe[3][12] .is_wysiwyg = "true";
defparam \pipe[3][12] .power_up = "low";

dffeas \pipe[1][12] (
	.clk(ctl_clk),
	.d(\pipe~6_combout ),
	.asdata(\pipe~2_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_12_1),
	.prn(vcc));
defparam \pipe[1][12] .is_wysiwyg = "true";
defparam \pipe[1][12] .power_up = "low";

dffeas \pipe[2][10] (
	.clk(ctl_clk),
	.d(\pipe~9_combout ),
	.asdata(\pipe~10_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_10_2),
	.prn(vcc));
defparam \pipe[2][10] .is_wysiwyg = "true";
defparam \pipe[2][10] .power_up = "low";

dffeas \pipe[3][10] (
	.clk(ctl_clk),
	.d(\pipe~11_combout ),
	.asdata(\pipe~9_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_10_3),
	.prn(vcc));
defparam \pipe[3][10] .is_wysiwyg = "true";
defparam \pipe[3][10] .power_up = "low";

dffeas \pipe[1][10] (
	.clk(ctl_clk),
	.d(\pipe~10_combout ),
	.asdata(\pipe~0_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_10_1),
	.prn(vcc));
defparam \pipe[1][10] .is_wysiwyg = "true";
defparam \pipe[1][10] .power_up = "low";

dffeas \pipe[2][11] (
	.clk(ctl_clk),
	.d(\pipe~12_combout ),
	.asdata(\pipe~13_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_11_2),
	.prn(vcc));
defparam \pipe[2][11] .is_wysiwyg = "true";
defparam \pipe[2][11] .power_up = "low";

dffeas \pipe[3][11] (
	.clk(ctl_clk),
	.d(\pipe~14_combout ),
	.asdata(\pipe~12_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_11_3),
	.prn(vcc));
defparam \pipe[3][11] .is_wysiwyg = "true";
defparam \pipe[3][11] .power_up = "low";

dffeas \pipe[1][11] (
	.clk(ctl_clk),
	.d(\pipe~13_combout ),
	.asdata(\pipe~3_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_11_1),
	.prn(vcc));
defparam \pipe[1][11] .is_wysiwyg = "true";
defparam \pipe[1][11] .power_up = "low";

dffeas \pipe[0][29] (
	.clk(ctl_clk),
	.d(\pipe~15_combout ),
	.asdata(size_1),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[0][5]~1_combout ),
	.q(pipe_29_0),
	.prn(vcc));
defparam \pipe[0][29] .is_wysiwyg = "true";
defparam \pipe[0][29] .power_up = "low";

dffeas \pipe[0][28] (
	.clk(ctl_clk),
	.d(\pipe~16_combout ),
	.asdata(size_0),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[0][5]~1_combout ),
	.q(pipe_28_0),
	.prn(vcc));
defparam \pipe[0][28] .is_wysiwyg = "true";
defparam \pipe[0][28] .power_up = "low";

dffeas \pipe[0][33] (
	.clk(ctl_clk),
	.d(\pipe~17_combout ),
	.asdata(read_req),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[0][5]~1_combout ),
	.q(pipe_33_0),
	.prn(vcc));
defparam \pipe[0][33] .is_wysiwyg = "true";
defparam \pipe[0][33] .power_up = "low";

dffeas \pipe[4][12] (
	.clk(ctl_clk),
	.d(\pipe~18_combout ),
	.asdata(\pipe~8_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_12_4),
	.prn(vcc));
defparam \pipe[4][12] .is_wysiwyg = "true";
defparam \pipe[4][12] .power_up = "low";

dffeas \pipe[4][11] (
	.clk(ctl_clk),
	.d(\pipe~19_combout ),
	.asdata(\pipe~14_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_11_4),
	.prn(vcc));
defparam \pipe[4][11] .is_wysiwyg = "true";
defparam \pipe[4][11] .power_up = "low";

dffeas \pipe[4][10] (
	.clk(ctl_clk),
	.d(\pipe~20_combout ),
	.asdata(\pipe~11_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_10_4),
	.prn(vcc));
defparam \pipe[4][10] .is_wysiwyg = "true";
defparam \pipe[4][10] .power_up = "low";

dffeas \pipe[5][25] (
	.clk(ctl_clk),
	.d(\pipe~22_combout ),
	.asdata(\pipe~23_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_25_5),
	.prn(vcc));
defparam \pipe[5][25] .is_wysiwyg = "true";
defparam \pipe[5][25] .power_up = "low";

dffeas \pipe[0][25] (
	.clk(ctl_clk),
	.d(\pipe~24_combout ),
	.asdata(row_addr_12),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[0][5]~1_combout ),
	.q(pipe_25_0),
	.prn(vcc));
defparam \pipe[0][25] .is_wysiwyg = "true";
defparam \pipe[0][25] .power_up = "low";

dffeas \pipe[5][26] (
	.clk(ctl_clk),
	.d(\pipe~25_combout ),
	.asdata(\pipe~26_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_26_5),
	.prn(vcc));
defparam \pipe[5][26] .is_wysiwyg = "true";
defparam \pipe[5][26] .power_up = "low";

dffeas \pipe[0][26] (
	.clk(ctl_clk),
	.d(\pipe~27_combout ),
	.asdata(row_addr_13),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[0][5]~1_combout ),
	.q(pipe_26_0),
	.prn(vcc));
defparam \pipe[0][26] .is_wysiwyg = "true";
defparam \pipe[0][26] .power_up = "low";

dffeas \pipe[5][24] (
	.clk(ctl_clk),
	.d(\pipe~28_combout ),
	.asdata(\pipe~29_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_24_5),
	.prn(vcc));
defparam \pipe[5][24] .is_wysiwyg = "true";
defparam \pipe[5][24] .power_up = "low";

dffeas \pipe[0][24] (
	.clk(ctl_clk),
	.d(\pipe~30_combout ),
	.asdata(row_addr_11),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[0][5]~1_combout ),
	.q(pipe_24_0),
	.prn(vcc));
defparam \pipe[0][24] .is_wysiwyg = "true";
defparam \pipe[0][24] .power_up = "low";

dffeas \pipe[5][22] (
	.clk(ctl_clk),
	.d(\pipe~31_combout ),
	.asdata(\pipe~32_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_22_5),
	.prn(vcc));
defparam \pipe[5][22] .is_wysiwyg = "true";
defparam \pipe[5][22] .power_up = "low";

dffeas \pipe[0][22] (
	.clk(ctl_clk),
	.d(\pipe~33_combout ),
	.asdata(row_addr_9),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[0][5]~1_combout ),
	.q(pipe_22_0),
	.prn(vcc));
defparam \pipe[0][22] .is_wysiwyg = "true";
defparam \pipe[0][22] .power_up = "low";

dffeas \pipe[5][23] (
	.clk(ctl_clk),
	.d(\pipe~34_combout ),
	.asdata(\pipe~35_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_23_5),
	.prn(vcc));
defparam \pipe[5][23] .is_wysiwyg = "true";
defparam \pipe[5][23] .power_up = "low";

dffeas \pipe[0][23] (
	.clk(ctl_clk),
	.d(\pipe~36_combout ),
	.asdata(row_addr_10),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[0][5]~1_combout ),
	.q(pipe_23_0),
	.prn(vcc));
defparam \pipe[0][23] .is_wysiwyg = "true";
defparam \pipe[0][23] .power_up = "low";

dffeas \pipe[5][21] (
	.clk(ctl_clk),
	.d(\pipe~37_combout ),
	.asdata(\pipe~38_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_21_5),
	.prn(vcc));
defparam \pipe[5][21] .is_wysiwyg = "true";
defparam \pipe[5][21] .power_up = "low";

dffeas \pipe[0][21] (
	.clk(ctl_clk),
	.d(\pipe~39_combout ),
	.asdata(row_addr_8),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[0][5]~1_combout ),
	.q(pipe_21_0),
	.prn(vcc));
defparam \pipe[0][21] .is_wysiwyg = "true";
defparam \pipe[0][21] .power_up = "low";

dffeas \pipe[5][19] (
	.clk(ctl_clk),
	.d(\pipe~40_combout ),
	.asdata(\pipe~41_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_19_5),
	.prn(vcc));
defparam \pipe[5][19] .is_wysiwyg = "true";
defparam \pipe[5][19] .power_up = "low";

dffeas \pipe[0][19] (
	.clk(ctl_clk),
	.d(\pipe~42_combout ),
	.asdata(row_addr_6),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[0][5]~1_combout ),
	.q(pipe_19_0),
	.prn(vcc));
defparam \pipe[0][19] .is_wysiwyg = "true";
defparam \pipe[0][19] .power_up = "low";

dffeas \pipe[5][20] (
	.clk(ctl_clk),
	.d(\pipe~43_combout ),
	.asdata(\pipe~44_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_20_5),
	.prn(vcc));
defparam \pipe[5][20] .is_wysiwyg = "true";
defparam \pipe[5][20] .power_up = "low";

dffeas \pipe[0][20] (
	.clk(ctl_clk),
	.d(\pipe~45_combout ),
	.asdata(row_addr_7),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[0][5]~1_combout ),
	.q(pipe_20_0),
	.prn(vcc));
defparam \pipe[0][20] .is_wysiwyg = "true";
defparam \pipe[0][20] .power_up = "low";

dffeas \pipe[5][15] (
	.clk(ctl_clk),
	.d(\pipe~46_combout ),
	.asdata(\pipe~47_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_15_5),
	.prn(vcc));
defparam \pipe[5][15] .is_wysiwyg = "true";
defparam \pipe[5][15] .power_up = "low";

dffeas \pipe[0][15] (
	.clk(ctl_clk),
	.d(\pipe~48_combout ),
	.asdata(row_addr_2),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[0][5]~1_combout ),
	.q(pipe_15_0),
	.prn(vcc));
defparam \pipe[0][15] .is_wysiwyg = "true";
defparam \pipe[0][15] .power_up = "low";

dffeas \pipe[5][13] (
	.clk(ctl_clk),
	.d(\pipe~49_combout ),
	.asdata(\pipe~50_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_13_5),
	.prn(vcc));
defparam \pipe[5][13] .is_wysiwyg = "true";
defparam \pipe[5][13] .power_up = "low";

dffeas \pipe[0][13] (
	.clk(ctl_clk),
	.d(\pipe~51_combout ),
	.asdata(row_addr_0),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[0][5]~1_combout ),
	.q(pipe_13_0),
	.prn(vcc));
defparam \pipe[0][13] .is_wysiwyg = "true";
defparam \pipe[0][13] .power_up = "low";

dffeas \pipe[5][14] (
	.clk(ctl_clk),
	.d(\pipe~52_combout ),
	.asdata(\pipe~53_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_14_5),
	.prn(vcc));
defparam \pipe[5][14] .is_wysiwyg = "true";
defparam \pipe[5][14] .power_up = "low";

dffeas \pipe[0][14] (
	.clk(ctl_clk),
	.d(\pipe~54_combout ),
	.asdata(row_addr_1),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[0][5]~1_combout ),
	.q(pipe_14_0),
	.prn(vcc));
defparam \pipe[0][14] .is_wysiwyg = "true";
defparam \pipe[0][14] .power_up = "low";

dffeas \pipe[5][18] (
	.clk(ctl_clk),
	.d(\pipe~55_combout ),
	.asdata(\pipe~56_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_18_5),
	.prn(vcc));
defparam \pipe[5][18] .is_wysiwyg = "true";
defparam \pipe[5][18] .power_up = "low";

dffeas \pipe[0][18] (
	.clk(ctl_clk),
	.d(\pipe~57_combout ),
	.asdata(row_addr_5),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[0][5]~1_combout ),
	.q(pipe_18_0),
	.prn(vcc));
defparam \pipe[0][18] .is_wysiwyg = "true";
defparam \pipe[0][18] .power_up = "low";

dffeas \pipe[5][16] (
	.clk(ctl_clk),
	.d(\pipe~58_combout ),
	.asdata(\pipe~59_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_16_5),
	.prn(vcc));
defparam \pipe[5][16] .is_wysiwyg = "true";
defparam \pipe[5][16] .power_up = "low";

dffeas \pipe[0][16] (
	.clk(ctl_clk),
	.d(\pipe~60_combout ),
	.asdata(row_addr_3),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[0][5]~1_combout ),
	.q(pipe_16_0),
	.prn(vcc));
defparam \pipe[0][16] .is_wysiwyg = "true";
defparam \pipe[0][16] .power_up = "low";

dffeas \pipe[5][17] (
	.clk(ctl_clk),
	.d(\pipe~61_combout ),
	.asdata(\pipe~62_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_17_5),
	.prn(vcc));
defparam \pipe[5][17] .is_wysiwyg = "true";
defparam \pipe[5][17] .power_up = "low";

dffeas \pipe[0][17] (
	.clk(ctl_clk),
	.d(\pipe~63_combout ),
	.asdata(row_addr_4),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[0][5]~1_combout ),
	.q(pipe_17_0),
	.prn(vcc));
defparam \pipe[0][17] .is_wysiwyg = "true";
defparam \pipe[0][17] .power_up = "low";

dffeas \pipe[5][12] (
	.clk(ctl_clk),
	.d(\pipe~64_combout ),
	.asdata(\pipe~18_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_12_5),
	.prn(vcc));
defparam \pipe[5][12] .is_wysiwyg = "true";
defparam \pipe[5][12] .power_up = "low";

dffeas \pipe[5][11] (
	.clk(ctl_clk),
	.d(\pipe~65_combout ),
	.asdata(\pipe~19_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_11_5),
	.prn(vcc));
defparam \pipe[5][11] .is_wysiwyg = "true";
defparam \pipe[5][11] .power_up = "low";

dffeas \pipe[5][10] (
	.clk(ctl_clk),
	.d(\pipe~66_combout ),
	.asdata(\pipe~20_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_10_5),
	.prn(vcc));
defparam \pipe[5][10] .is_wysiwyg = "true";
defparam \pipe[5][10] .power_up = "low";

dffeas \pipe[3][25] (
	.clk(ctl_clk),
	.d(\pipe~67_combout ),
	.asdata(\pipe~68_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_25_3),
	.prn(vcc));
defparam \pipe[3][25] .is_wysiwyg = "true";
defparam \pipe[3][25] .power_up = "low";

dffeas \pipe[3][26] (
	.clk(ctl_clk),
	.d(\pipe~69_combout ),
	.asdata(\pipe~70_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_26_3),
	.prn(vcc));
defparam \pipe[3][26] .is_wysiwyg = "true";
defparam \pipe[3][26] .power_up = "low";

dffeas \pipe[3][24] (
	.clk(ctl_clk),
	.d(\pipe~71_combout ),
	.asdata(\pipe~72_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_24_3),
	.prn(vcc));
defparam \pipe[3][24] .is_wysiwyg = "true";
defparam \pipe[3][24] .power_up = "low";

dffeas \pipe[3][22] (
	.clk(ctl_clk),
	.d(\pipe~73_combout ),
	.asdata(\pipe~74_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_22_3),
	.prn(vcc));
defparam \pipe[3][22] .is_wysiwyg = "true";
defparam \pipe[3][22] .power_up = "low";

dffeas \pipe[3][23] (
	.clk(ctl_clk),
	.d(\pipe~75_combout ),
	.asdata(\pipe~76_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_23_3),
	.prn(vcc));
defparam \pipe[3][23] .is_wysiwyg = "true";
defparam \pipe[3][23] .power_up = "low";

dffeas \pipe[3][21] (
	.clk(ctl_clk),
	.d(\pipe~77_combout ),
	.asdata(\pipe~78_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_21_3),
	.prn(vcc));
defparam \pipe[3][21] .is_wysiwyg = "true";
defparam \pipe[3][21] .power_up = "low";

dffeas \pipe[3][19] (
	.clk(ctl_clk),
	.d(\pipe~79_combout ),
	.asdata(\pipe~80_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_19_3),
	.prn(vcc));
defparam \pipe[3][19] .is_wysiwyg = "true";
defparam \pipe[3][19] .power_up = "low";

dffeas \pipe[3][20] (
	.clk(ctl_clk),
	.d(\pipe~81_combout ),
	.asdata(\pipe~82_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_20_3),
	.prn(vcc));
defparam \pipe[3][20] .is_wysiwyg = "true";
defparam \pipe[3][20] .power_up = "low";

dffeas \pipe[3][15] (
	.clk(ctl_clk),
	.d(\pipe~83_combout ),
	.asdata(\pipe~84_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_15_3),
	.prn(vcc));
defparam \pipe[3][15] .is_wysiwyg = "true";
defparam \pipe[3][15] .power_up = "low";

dffeas \pipe[3][13] (
	.clk(ctl_clk),
	.d(\pipe~85_combout ),
	.asdata(\pipe~86_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_13_3),
	.prn(vcc));
defparam \pipe[3][13] .is_wysiwyg = "true";
defparam \pipe[3][13] .power_up = "low";

dffeas \pipe[3][14] (
	.clk(ctl_clk),
	.d(\pipe~87_combout ),
	.asdata(\pipe~88_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_14_3),
	.prn(vcc));
defparam \pipe[3][14] .is_wysiwyg = "true";
defparam \pipe[3][14] .power_up = "low";

dffeas \pipe[3][18] (
	.clk(ctl_clk),
	.d(\pipe~89_combout ),
	.asdata(\pipe~90_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_18_3),
	.prn(vcc));
defparam \pipe[3][18] .is_wysiwyg = "true";
defparam \pipe[3][18] .power_up = "low";

dffeas \pipe[3][16] (
	.clk(ctl_clk),
	.d(\pipe~91_combout ),
	.asdata(\pipe~92_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_16_3),
	.prn(vcc));
defparam \pipe[3][16] .is_wysiwyg = "true";
defparam \pipe[3][16] .power_up = "low";

dffeas \pipe[3][17] (
	.clk(ctl_clk),
	.d(\pipe~93_combout ),
	.asdata(\pipe~94_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_17_3),
	.prn(vcc));
defparam \pipe[3][17] .is_wysiwyg = "true";
defparam \pipe[3][17] .power_up = "low";

dffeas \pipe[4][25] (
	.clk(ctl_clk),
	.d(\pipe~23_combout ),
	.asdata(\pipe~67_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_25_4),
	.prn(vcc));
defparam \pipe[4][25] .is_wysiwyg = "true";
defparam \pipe[4][25] .power_up = "low";

dffeas \pipe[4][26] (
	.clk(ctl_clk),
	.d(\pipe~26_combout ),
	.asdata(\pipe~69_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_26_4),
	.prn(vcc));
defparam \pipe[4][26] .is_wysiwyg = "true";
defparam \pipe[4][26] .power_up = "low";

dffeas \pipe[4][24] (
	.clk(ctl_clk),
	.d(\pipe~29_combout ),
	.asdata(\pipe~71_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_24_4),
	.prn(vcc));
defparam \pipe[4][24] .is_wysiwyg = "true";
defparam \pipe[4][24] .power_up = "low";

dffeas \pipe[4][22] (
	.clk(ctl_clk),
	.d(\pipe~32_combout ),
	.asdata(\pipe~73_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_22_4),
	.prn(vcc));
defparam \pipe[4][22] .is_wysiwyg = "true";
defparam \pipe[4][22] .power_up = "low";

dffeas \pipe[4][23] (
	.clk(ctl_clk),
	.d(\pipe~35_combout ),
	.asdata(\pipe~75_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_23_4),
	.prn(vcc));
defparam \pipe[4][23] .is_wysiwyg = "true";
defparam \pipe[4][23] .power_up = "low";

dffeas \pipe[4][21] (
	.clk(ctl_clk),
	.d(\pipe~38_combout ),
	.asdata(\pipe~77_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_21_4),
	.prn(vcc));
defparam \pipe[4][21] .is_wysiwyg = "true";
defparam \pipe[4][21] .power_up = "low";

dffeas \pipe[4][19] (
	.clk(ctl_clk),
	.d(\pipe~41_combout ),
	.asdata(\pipe~79_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_19_4),
	.prn(vcc));
defparam \pipe[4][19] .is_wysiwyg = "true";
defparam \pipe[4][19] .power_up = "low";

dffeas \pipe[4][20] (
	.clk(ctl_clk),
	.d(\pipe~44_combout ),
	.asdata(\pipe~81_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_20_4),
	.prn(vcc));
defparam \pipe[4][20] .is_wysiwyg = "true";
defparam \pipe[4][20] .power_up = "low";

dffeas \pipe[4][15] (
	.clk(ctl_clk),
	.d(\pipe~47_combout ),
	.asdata(\pipe~83_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_15_4),
	.prn(vcc));
defparam \pipe[4][15] .is_wysiwyg = "true";
defparam \pipe[4][15] .power_up = "low";

dffeas \pipe[4][13] (
	.clk(ctl_clk),
	.d(\pipe~50_combout ),
	.asdata(\pipe~85_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_13_4),
	.prn(vcc));
defparam \pipe[4][13] .is_wysiwyg = "true";
defparam \pipe[4][13] .power_up = "low";

dffeas \pipe[4][14] (
	.clk(ctl_clk),
	.d(\pipe~53_combout ),
	.asdata(\pipe~87_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_14_4),
	.prn(vcc));
defparam \pipe[4][14] .is_wysiwyg = "true";
defparam \pipe[4][14] .power_up = "low";

dffeas \pipe[4][18] (
	.clk(ctl_clk),
	.d(\pipe~56_combout ),
	.asdata(\pipe~89_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_18_4),
	.prn(vcc));
defparam \pipe[4][18] .is_wysiwyg = "true";
defparam \pipe[4][18] .power_up = "low";

dffeas \pipe[4][16] (
	.clk(ctl_clk),
	.d(\pipe~59_combout ),
	.asdata(\pipe~91_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_16_4),
	.prn(vcc));
defparam \pipe[4][16] .is_wysiwyg = "true";
defparam \pipe[4][16] .power_up = "low";

dffeas \pipe[4][17] (
	.clk(ctl_clk),
	.d(\pipe~62_combout ),
	.asdata(\pipe~93_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_17_4),
	.prn(vcc));
defparam \pipe[4][17] .is_wysiwyg = "true";
defparam \pipe[4][17] .power_up = "low";

dffeas \pipe[6][12] (
	.clk(ctl_clk),
	.d(\pipe~95_combout ),
	.asdata(\pipe~64_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_12_6),
	.prn(vcc));
defparam \pipe[6][12] .is_wysiwyg = "true";
defparam \pipe[6][12] .power_up = "low";

dffeas \pipe[6][11] (
	.clk(ctl_clk),
	.d(\pipe~96_combout ),
	.asdata(\pipe~65_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_11_6),
	.prn(vcc));
defparam \pipe[6][11] .is_wysiwyg = "true";
defparam \pipe[6][11] .power_up = "low";

dffeas \pipe[6][10] (
	.clk(ctl_clk),
	.d(\pipe~97_combout ),
	.asdata(\pipe~66_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_10_6),
	.prn(vcc));
defparam \pipe[6][10] .is_wysiwyg = "true";
defparam \pipe[6][10] .power_up = "low";

dffeas \pipe[6][25] (
	.clk(ctl_clk),
	.d(\pipe~98_combout ),
	.asdata(\pipe~22_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_25_6),
	.prn(vcc));
defparam \pipe[6][25] .is_wysiwyg = "true";
defparam \pipe[6][25] .power_up = "low";

dffeas \pipe[6][26] (
	.clk(ctl_clk),
	.d(\pipe~99_combout ),
	.asdata(\pipe~25_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_26_6),
	.prn(vcc));
defparam \pipe[6][26] .is_wysiwyg = "true";
defparam \pipe[6][26] .power_up = "low";

dffeas \pipe[6][24] (
	.clk(ctl_clk),
	.d(\pipe~100_combout ),
	.asdata(\pipe~28_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_24_6),
	.prn(vcc));
defparam \pipe[6][24] .is_wysiwyg = "true";
defparam \pipe[6][24] .power_up = "low";

dffeas \pipe[6][22] (
	.clk(ctl_clk),
	.d(\pipe~101_combout ),
	.asdata(\pipe~31_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_22_6),
	.prn(vcc));
defparam \pipe[6][22] .is_wysiwyg = "true";
defparam \pipe[6][22] .power_up = "low";

dffeas \pipe[6][23] (
	.clk(ctl_clk),
	.d(\pipe~102_combout ),
	.asdata(\pipe~34_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_23_6),
	.prn(vcc));
defparam \pipe[6][23] .is_wysiwyg = "true";
defparam \pipe[6][23] .power_up = "low";

dffeas \pipe[6][21] (
	.clk(ctl_clk),
	.d(\pipe~103_combout ),
	.asdata(\pipe~37_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_21_6),
	.prn(vcc));
defparam \pipe[6][21] .is_wysiwyg = "true";
defparam \pipe[6][21] .power_up = "low";

dffeas \pipe[6][19] (
	.clk(ctl_clk),
	.d(\pipe~104_combout ),
	.asdata(\pipe~40_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_19_6),
	.prn(vcc));
defparam \pipe[6][19] .is_wysiwyg = "true";
defparam \pipe[6][19] .power_up = "low";

dffeas \pipe[6][20] (
	.clk(ctl_clk),
	.d(\pipe~105_combout ),
	.asdata(\pipe~43_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_20_6),
	.prn(vcc));
defparam \pipe[6][20] .is_wysiwyg = "true";
defparam \pipe[6][20] .power_up = "low";

dffeas \pipe[6][15] (
	.clk(ctl_clk),
	.d(\pipe~106_combout ),
	.asdata(\pipe~46_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_15_6),
	.prn(vcc));
defparam \pipe[6][15] .is_wysiwyg = "true";
defparam \pipe[6][15] .power_up = "low";

dffeas \pipe[6][13] (
	.clk(ctl_clk),
	.d(\pipe~107_combout ),
	.asdata(\pipe~49_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_13_6),
	.prn(vcc));
defparam \pipe[6][13] .is_wysiwyg = "true";
defparam \pipe[6][13] .power_up = "low";

dffeas \pipe[6][14] (
	.clk(ctl_clk),
	.d(\pipe~108_combout ),
	.asdata(\pipe~52_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_14_6),
	.prn(vcc));
defparam \pipe[6][14] .is_wysiwyg = "true";
defparam \pipe[6][14] .power_up = "low";

dffeas \pipe[6][18] (
	.clk(ctl_clk),
	.d(\pipe~109_combout ),
	.asdata(\pipe~55_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_18_6),
	.prn(vcc));
defparam \pipe[6][18] .is_wysiwyg = "true";
defparam \pipe[6][18] .power_up = "low";

dffeas \pipe[6][16] (
	.clk(ctl_clk),
	.d(\pipe~110_combout ),
	.asdata(\pipe~58_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_16_6),
	.prn(vcc));
defparam \pipe[6][16] .is_wysiwyg = "true";
defparam \pipe[6][16] .power_up = "low";

dffeas \pipe[6][17] (
	.clk(ctl_clk),
	.d(\pipe~111_combout ),
	.asdata(\pipe~61_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_17_6),
	.prn(vcc));
defparam \pipe[6][17] .is_wysiwyg = "true";
defparam \pipe[6][17] .power_up = "low";

dffeas \pipe[7][26] (
	.clk(ctl_clk),
	.d(\pipe~112_combout ),
	.asdata(\pipe~99_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_26_7),
	.prn(vcc));
defparam \pipe[7][26] .is_wysiwyg = "true";
defparam \pipe[7][26] .power_up = "low";

dffeas \pipe[7][24] (
	.clk(ctl_clk),
	.d(\pipe~113_combout ),
	.asdata(\pipe~100_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_24_7),
	.prn(vcc));
defparam \pipe[7][24] .is_wysiwyg = "true";
defparam \pipe[7][24] .power_up = "low";

dffeas \pipe[7][25] (
	.clk(ctl_clk),
	.d(\pipe~114_combout ),
	.asdata(\pipe~98_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_25_7),
	.prn(vcc));
defparam \pipe[7][25] .is_wysiwyg = "true";
defparam \pipe[7][25] .power_up = "low";

dffeas \pipe[7][23] (
	.clk(ctl_clk),
	.d(\pipe~115_combout ),
	.asdata(\pipe~102_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_23_7),
	.prn(vcc));
defparam \pipe[7][23] .is_wysiwyg = "true";
defparam \pipe[7][23] .power_up = "low";

dffeas \pipe[7][21] (
	.clk(ctl_clk),
	.d(\pipe~116_combout ),
	.asdata(\pipe~103_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_21_7),
	.prn(vcc));
defparam \pipe[7][21] .is_wysiwyg = "true";
defparam \pipe[7][21] .power_up = "low";

dffeas \pipe[7][22] (
	.clk(ctl_clk),
	.d(\pipe~117_combout ),
	.asdata(\pipe~101_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_22_7),
	.prn(vcc));
defparam \pipe[7][22] .is_wysiwyg = "true";
defparam \pipe[7][22] .power_up = "low";

dffeas \pipe[7][20] (
	.clk(ctl_clk),
	.d(\pipe~118_combout ),
	.asdata(\pipe~105_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_20_7),
	.prn(vcc));
defparam \pipe[7][20] .is_wysiwyg = "true";
defparam \pipe[7][20] .power_up = "low";

dffeas \pipe[7][18] (
	.clk(ctl_clk),
	.d(\pipe~119_combout ),
	.asdata(\pipe~109_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_18_7),
	.prn(vcc));
defparam \pipe[7][18] .is_wysiwyg = "true";
defparam \pipe[7][18] .power_up = "low";

dffeas \pipe[7][19] (
	.clk(ctl_clk),
	.d(\pipe~120_combout ),
	.asdata(\pipe~104_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_19_7),
	.prn(vcc));
defparam \pipe[7][19] .is_wysiwyg = "true";
defparam \pipe[7][19] .power_up = "low";

dffeas \pipe[7][17] (
	.clk(ctl_clk),
	.d(\pipe~121_combout ),
	.asdata(\pipe~111_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_17_7),
	.prn(vcc));
defparam \pipe[7][17] .is_wysiwyg = "true";
defparam \pipe[7][17] .power_up = "low";

dffeas \pipe[7][15] (
	.clk(ctl_clk),
	.d(\pipe~122_combout ),
	.asdata(\pipe~106_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_15_7),
	.prn(vcc));
defparam \pipe[7][15] .is_wysiwyg = "true";
defparam \pipe[7][15] .power_up = "low";

dffeas \pipe[7][16] (
	.clk(ctl_clk),
	.d(\pipe~123_combout ),
	.asdata(\pipe~110_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_16_7),
	.prn(vcc));
defparam \pipe[7][16] .is_wysiwyg = "true";
defparam \pipe[7][16] .power_up = "low";

dffeas \pipe[7][11] (
	.clk(ctl_clk),
	.d(\pipe~124_combout ),
	.asdata(\pipe~96_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_11_7),
	.prn(vcc));
defparam \pipe[7][11] .is_wysiwyg = "true";
defparam \pipe[7][11] .power_up = "low";

dffeas \pipe[7][10] (
	.clk(ctl_clk),
	.d(\pipe~125_combout ),
	.asdata(\pipe~97_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_10_7),
	.prn(vcc));
defparam \pipe[7][10] .is_wysiwyg = "true";
defparam \pipe[7][10] .power_up = "low";

dffeas \pipe[7][14] (
	.clk(ctl_clk),
	.d(\pipe~126_combout ),
	.asdata(\pipe~108_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_14_7),
	.prn(vcc));
defparam \pipe[7][14] .is_wysiwyg = "true";
defparam \pipe[7][14] .power_up = "low";

dffeas \pipe[7][12] (
	.clk(ctl_clk),
	.d(\pipe~127_combout ),
	.asdata(\pipe~95_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_12_7),
	.prn(vcc));
defparam \pipe[7][12] .is_wysiwyg = "true";
defparam \pipe[7][12] .power_up = "low";

dffeas \pipe[7][13] (
	.clk(ctl_clk),
	.d(\pipe~128_combout ),
	.asdata(\pipe~107_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_13_7),
	.prn(vcc));
defparam \pipe[7][13] .is_wysiwyg = "true";
defparam \pipe[7][13] .power_up = "low";

dffeas \pipe[2][25] (
	.clk(ctl_clk),
	.d(\pipe~68_combout ),
	.asdata(\pipe~129_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_25_2),
	.prn(vcc));
defparam \pipe[2][25] .is_wysiwyg = "true";
defparam \pipe[2][25] .power_up = "low";

dffeas \pipe[2][26] (
	.clk(ctl_clk),
	.d(\pipe~70_combout ),
	.asdata(\pipe~130_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_26_2),
	.prn(vcc));
defparam \pipe[2][26] .is_wysiwyg = "true";
defparam \pipe[2][26] .power_up = "low";

dffeas \pipe[2][24] (
	.clk(ctl_clk),
	.d(\pipe~72_combout ),
	.asdata(\pipe~131_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_24_2),
	.prn(vcc));
defparam \pipe[2][24] .is_wysiwyg = "true";
defparam \pipe[2][24] .power_up = "low";

dffeas \pipe[2][22] (
	.clk(ctl_clk),
	.d(\pipe~74_combout ),
	.asdata(\pipe~132_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_22_2),
	.prn(vcc));
defparam \pipe[2][22] .is_wysiwyg = "true";
defparam \pipe[2][22] .power_up = "low";

dffeas \pipe[2][23] (
	.clk(ctl_clk),
	.d(\pipe~76_combout ),
	.asdata(\pipe~133_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_23_2),
	.prn(vcc));
defparam \pipe[2][23] .is_wysiwyg = "true";
defparam \pipe[2][23] .power_up = "low";

dffeas \pipe[2][21] (
	.clk(ctl_clk),
	.d(\pipe~78_combout ),
	.asdata(\pipe~134_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_21_2),
	.prn(vcc));
defparam \pipe[2][21] .is_wysiwyg = "true";
defparam \pipe[2][21] .power_up = "low";

dffeas \pipe[2][19] (
	.clk(ctl_clk),
	.d(\pipe~80_combout ),
	.asdata(\pipe~135_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_19_2),
	.prn(vcc));
defparam \pipe[2][19] .is_wysiwyg = "true";
defparam \pipe[2][19] .power_up = "low";

dffeas \pipe[2][20] (
	.clk(ctl_clk),
	.d(\pipe~82_combout ),
	.asdata(\pipe~136_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_20_2),
	.prn(vcc));
defparam \pipe[2][20] .is_wysiwyg = "true";
defparam \pipe[2][20] .power_up = "low";

dffeas \pipe[2][15] (
	.clk(ctl_clk),
	.d(\pipe~84_combout ),
	.asdata(\pipe~137_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_15_2),
	.prn(vcc));
defparam \pipe[2][15] .is_wysiwyg = "true";
defparam \pipe[2][15] .power_up = "low";

dffeas \pipe[2][13] (
	.clk(ctl_clk),
	.d(\pipe~86_combout ),
	.asdata(\pipe~138_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_13_2),
	.prn(vcc));
defparam \pipe[2][13] .is_wysiwyg = "true";
defparam \pipe[2][13] .power_up = "low";

dffeas \pipe[2][14] (
	.clk(ctl_clk),
	.d(\pipe~88_combout ),
	.asdata(\pipe~139_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_14_2),
	.prn(vcc));
defparam \pipe[2][14] .is_wysiwyg = "true";
defparam \pipe[2][14] .power_up = "low";

dffeas \pipe[2][18] (
	.clk(ctl_clk),
	.d(\pipe~90_combout ),
	.asdata(\pipe~140_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_18_2),
	.prn(vcc));
defparam \pipe[2][18] .is_wysiwyg = "true";
defparam \pipe[2][18] .power_up = "low";

dffeas \pipe[2][16] (
	.clk(ctl_clk),
	.d(\pipe~92_combout ),
	.asdata(\pipe~141_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_16_2),
	.prn(vcc));
defparam \pipe[2][16] .is_wysiwyg = "true";
defparam \pipe[2][16] .power_up = "low";

dffeas \pipe[2][17] (
	.clk(ctl_clk),
	.d(\pipe~94_combout ),
	.asdata(\pipe~142_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_17_2),
	.prn(vcc));
defparam \pipe[2][17] .is_wysiwyg = "true";
defparam \pipe[2][17] .power_up = "low";

dffeas \pipe[1][25] (
	.clk(ctl_clk),
	.d(\pipe~129_combout ),
	.asdata(\pipe~24_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_25_1),
	.prn(vcc));
defparam \pipe[1][25] .is_wysiwyg = "true";
defparam \pipe[1][25] .power_up = "low";

dffeas \pipe[1][26] (
	.clk(ctl_clk),
	.d(\pipe~130_combout ),
	.asdata(\pipe~27_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_26_1),
	.prn(vcc));
defparam \pipe[1][26] .is_wysiwyg = "true";
defparam \pipe[1][26] .power_up = "low";

dffeas \pipe[1][24] (
	.clk(ctl_clk),
	.d(\pipe~131_combout ),
	.asdata(\pipe~30_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_24_1),
	.prn(vcc));
defparam \pipe[1][24] .is_wysiwyg = "true";
defparam \pipe[1][24] .power_up = "low";

dffeas \pipe[1][22] (
	.clk(ctl_clk),
	.d(\pipe~132_combout ),
	.asdata(\pipe~33_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_22_1),
	.prn(vcc));
defparam \pipe[1][22] .is_wysiwyg = "true";
defparam \pipe[1][22] .power_up = "low";

dffeas \pipe[1][23] (
	.clk(ctl_clk),
	.d(\pipe~133_combout ),
	.asdata(\pipe~36_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_23_1),
	.prn(vcc));
defparam \pipe[1][23] .is_wysiwyg = "true";
defparam \pipe[1][23] .power_up = "low";

dffeas \pipe[1][21] (
	.clk(ctl_clk),
	.d(\pipe~134_combout ),
	.asdata(\pipe~39_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_21_1),
	.prn(vcc));
defparam \pipe[1][21] .is_wysiwyg = "true";
defparam \pipe[1][21] .power_up = "low";

dffeas \pipe[1][19] (
	.clk(ctl_clk),
	.d(\pipe~135_combout ),
	.asdata(\pipe~42_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_19_1),
	.prn(vcc));
defparam \pipe[1][19] .is_wysiwyg = "true";
defparam \pipe[1][19] .power_up = "low";

dffeas \pipe[1][20] (
	.clk(ctl_clk),
	.d(\pipe~136_combout ),
	.asdata(\pipe~45_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_20_1),
	.prn(vcc));
defparam \pipe[1][20] .is_wysiwyg = "true";
defparam \pipe[1][20] .power_up = "low";

dffeas \pipe[1][15] (
	.clk(ctl_clk),
	.d(\pipe~137_combout ),
	.asdata(\pipe~48_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_15_1),
	.prn(vcc));
defparam \pipe[1][15] .is_wysiwyg = "true";
defparam \pipe[1][15] .power_up = "low";

dffeas \pipe[1][13] (
	.clk(ctl_clk),
	.d(\pipe~138_combout ),
	.asdata(\pipe~51_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_13_1),
	.prn(vcc));
defparam \pipe[1][13] .is_wysiwyg = "true";
defparam \pipe[1][13] .power_up = "low";

dffeas \pipe[1][14] (
	.clk(ctl_clk),
	.d(\pipe~139_combout ),
	.asdata(\pipe~54_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_14_1),
	.prn(vcc));
defparam \pipe[1][14] .is_wysiwyg = "true";
defparam \pipe[1][14] .power_up = "low";

dffeas \pipe[1][18] (
	.clk(ctl_clk),
	.d(\pipe~140_combout ),
	.asdata(\pipe~57_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_18_1),
	.prn(vcc));
defparam \pipe[1][18] .is_wysiwyg = "true";
defparam \pipe[1][18] .power_up = "low";

dffeas \pipe[1][16] (
	.clk(ctl_clk),
	.d(\pipe~141_combout ),
	.asdata(\pipe~60_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_16_1),
	.prn(vcc));
defparam \pipe[1][16] .is_wysiwyg = "true";
defparam \pipe[1][16] .power_up = "low";

dffeas \pipe[1][17] (
	.clk(ctl_clk),
	.d(\pipe~142_combout ),
	.asdata(\pipe~63_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(pipe_17_1),
	.prn(vcc));
defparam \pipe[1][17] .is_wysiwyg = "true";
defparam \pipe[1][17] .power_up = "low";

dffeas \pipe[0][2] (
	.clk(ctl_clk),
	.d(\pipe~147_combout ),
	.asdata(col_addr_2),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[0][5]~1_combout ),
	.q(pipe_2_0),
	.prn(vcc));
defparam \pipe[0][2] .is_wysiwyg = "true";
defparam \pipe[0][2] .power_up = "low";

dffeas \pipe[0][3] (
	.clk(ctl_clk),
	.d(\pipe~161_combout ),
	.asdata(col_addr_3),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[0][5]~1_combout ),
	.q(pipe_3_0),
	.prn(vcc));
defparam \pipe[0][3] .is_wysiwyg = "true";
defparam \pipe[0][3] .power_up = "low";

dffeas \pipe[0][4] (
	.clk(ctl_clk),
	.d(\pipe~162_combout ),
	.asdata(col_addr_4),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[0][5]~1_combout ),
	.q(pipe_4_0),
	.prn(vcc));
defparam \pipe[0][4] .is_wysiwyg = "true";
defparam \pipe[0][4] .power_up = "low";

dffeas \pipe[0][5] (
	.clk(ctl_clk),
	.d(\pipe~163_combout ),
	.asdata(col_addr_5),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[0][5]~1_combout ),
	.q(pipe_5_0),
	.prn(vcc));
defparam \pipe[0][5] .is_wysiwyg = "true";
defparam \pipe[0][5] .power_up = "low";

dffeas \pipe[0][6] (
	.clk(ctl_clk),
	.d(\pipe~164_combout ),
	.asdata(col_addr_6),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[0][5]~1_combout ),
	.q(pipe_6_0),
	.prn(vcc));
defparam \pipe[0][6] .is_wysiwyg = "true";
defparam \pipe[0][6] .power_up = "low";

dffeas \pipe[0][7] (
	.clk(ctl_clk),
	.d(\pipe~165_combout ),
	.asdata(col_addr_7),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[0][5]~1_combout ),
	.q(pipe_7_0),
	.prn(vcc));
defparam \pipe[0][7] .is_wysiwyg = "true";
defparam \pipe[0][7] .power_up = "low";

dffeas \pipe[0][8] (
	.clk(ctl_clk),
	.d(\pipe~166_combout ),
	.asdata(col_addr_8),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[0][5]~1_combout ),
	.q(pipe_8_0),
	.prn(vcc));
defparam \pipe[0][8] .is_wysiwyg = "true";
defparam \pipe[0][8] .power_up = "low";

dffeas \pipe[0][9] (
	.clk(ctl_clk),
	.d(\pipe~167_combout ),
	.asdata(col_addr_9),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[0][5]~1_combout ),
	.q(pipe_9_0),
	.prn(vcc));
defparam \pipe[0][9] .is_wysiwyg = "true";
defparam \pipe[0][9] .power_up = "low";

dffeas \pipefull[7] (
	.clk(ctl_clk),
	.d(\pipefull~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(pipefull_7),
	.prn(vcc));
defparam \pipefull[7] .is_wysiwyg = "true";
defparam \pipefull[7] .power_up = "low";

dffeas \pipefull[6] (
	.clk(ctl_clk),
	.d(\pipefull~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(pipefull_6),
	.prn(vcc));
defparam \pipefull[6] .is_wysiwyg = "true";
defparam \pipefull[6] .power_up = "low";

dffeas \pipefull[0] (
	.clk(ctl_clk),
	.d(\pipefull~2_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(pipefull_0),
	.prn(vcc));
defparam \pipefull[0] .is_wysiwyg = "true";
defparam \pipefull[0] .power_up = "low";

dffeas \pipefull[5] (
	.clk(ctl_clk),
	.d(\pipefull~3_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(pipefull_5),
	.prn(vcc));
defparam \pipefull[5] .is_wysiwyg = "true";
defparam \pipefull[5] .power_up = "low";

dffeas \pipefull[1] (
	.clk(ctl_clk),
	.d(\pipefull~4_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(pipefull_1),
	.prn(vcc));
defparam \pipefull[1] .is_wysiwyg = "true";
defparam \pipefull[1] .power_up = "low";

dffeas \pipefull[4] (
	.clk(ctl_clk),
	.d(\pipefull~5_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(pipefull_4),
	.prn(vcc));
defparam \pipefull[4] .is_wysiwyg = "true";
defparam \pipefull[4] .power_up = "low";

dffeas \pipefull[2] (
	.clk(ctl_clk),
	.d(\pipefull~6_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(pipefull_2),
	.prn(vcc));
defparam \pipefull[2] .is_wysiwyg = "true";
defparam \pipefull[2] .power_up = "low";

dffeas \pipefull[3] (
	.clk(ctl_clk),
	.d(\pipefull~7_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(pipefull_3),
	.prn(vcc));
defparam \pipefull[3] .is_wysiwyg = "true";
defparam \pipefull[3] .power_up = "low";

arriaii_lcell_comb \pipe~0 (
	.dataa(!pipefull_0),
	.datab(!pipefull_1),
	.datac(!pipe_10_1),
	.datad(!bank_addr_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~0 .extended_lut = "off";
defparam \pipe~0 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~0 .shared_arith = "off";

arriaii_lcell_comb \pipe[0][5]~1 (
	.dataa(!fetch),
	.datab(!read_req),
	.datac(!write_req),
	.datad(!pipefull_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe[0][5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe[0][5]~1 .extended_lut = "off";
defparam \pipe[0][5]~1 .lut_mask = 64'h7F557F557F557F55;
defparam \pipe[0][5]~1 .shared_arith = "off";

arriaii_lcell_comb \pipe~2 (
	.dataa(!pipefull_0),
	.datab(!pipefull_1),
	.datac(!pipe_12_1),
	.datad(!bank_addr_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~2 .extended_lut = "off";
defparam \pipe~2 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~2 .shared_arith = "off";

arriaii_lcell_comb \pipe~3 (
	.dataa(!pipefull_0),
	.datab(!pipefull_1),
	.datac(!pipe_11_1),
	.datad(!bank_addr_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~3 .extended_lut = "off";
defparam \pipe~3 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~3 .shared_arith = "off";

arriaii_lcell_comb \pipe~192 (
	.dataa(!write_req),
	.datab(!\pipe[7][32]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~192_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~192 .extended_lut = "off";
defparam \pipe~192 .lut_mask = 64'h1111111111111111;
defparam \pipe~192 .shared_arith = "off";

arriaii_lcell_comb \pipe[1][11]~7 (
	.dataa(!fetch),
	.datab(!read_req),
	.datac(!write_req),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe[1][11]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe[1][11]~7 .extended_lut = "off";
defparam \pipe[1][11]~7 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \pipe[1][11]~7 .shared_arith = "off";

dffeas \pipe[7][32] (
	.clk(ctl_clk),
	.d(\pipe~192_combout ),
	.asdata(\pipe~180_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[7][32]~q ),
	.prn(vcc));
defparam \pipe[7][32] .is_wysiwyg = "true";
defparam \pipe[7][32] .power_up = "low";

arriaii_lcell_comb \pipe~180 (
	.dataa(!pipefull_7),
	.datab(!write_req),
	.datac(!pipefull_6),
	.datad(!\pipe[7][32]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~180_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~180 .extended_lut = "off";
defparam \pipe~180 .lut_mask = 64'h02F702F702F702F7;
defparam \pipe~180 .shared_arith = "off";

dffeas \pipe[6][32] (
	.clk(ctl_clk),
	.d(\pipe~180_combout ),
	.asdata(\pipe~168_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[6][32]~q ),
	.prn(vcc));
defparam \pipe[6][32] .is_wysiwyg = "true";
defparam \pipe[6][32] .power_up = "low";

arriaii_lcell_comb \pipe~168 (
	.dataa(!write_req),
	.datab(!pipefull_6),
	.datac(!pipefull_5),
	.datad(!\pipe[6][32]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~168_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~168 .extended_lut = "off";
defparam \pipe~168 .lut_mask = 64'h04F704F704F704F7;
defparam \pipe~168 .shared_arith = "off";

dffeas \pipe[5][32] (
	.clk(ctl_clk),
	.d(\pipe~168_combout ),
	.asdata(\pipe~156_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[5][32]~q ),
	.prn(vcc));
defparam \pipe[5][32] .is_wysiwyg = "true";
defparam \pipe[5][32] .power_up = "low";

arriaii_lcell_comb \pipe~156 (
	.dataa(!write_req),
	.datab(!pipefull_5),
	.datac(!pipefull_4),
	.datad(!\pipe[5][32]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~156_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~156 .extended_lut = "off";
defparam \pipe~156 .lut_mask = 64'h04F704F704F704F7;
defparam \pipe~156 .shared_arith = "off";

dffeas \pipe[4][32] (
	.clk(ctl_clk),
	.d(\pipe~156_combout ),
	.asdata(\pipe~151_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[4][32]~q ),
	.prn(vcc));
defparam \pipe[4][32] .is_wysiwyg = "true";
defparam \pipe[4][32] .power_up = "low";

arriaii_lcell_comb \pipe~151 (
	.dataa(!write_req),
	.datab(!pipefull_4),
	.datac(!pipefull_3),
	.datad(!\pipe[4][32]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~151_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~151 .extended_lut = "off";
defparam \pipe~151 .lut_mask = 64'h04F704F704F704F7;
defparam \pipe~151 .shared_arith = "off";

dffeas \pipe[3][32] (
	.clk(ctl_clk),
	.d(\pipe~151_combout ),
	.asdata(\pipe~146_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[3][32]~q ),
	.prn(vcc));
defparam \pipe[3][32] .is_wysiwyg = "true";
defparam \pipe[3][32] .power_up = "low";

arriaii_lcell_comb \pipe~146 (
	.dataa(!write_req),
	.datab(!pipefull_2),
	.datac(!pipefull_3),
	.datad(!\pipe[3][32]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~146_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~146 .extended_lut = "off";
defparam \pipe~146 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \pipe~146 .shared_arith = "off";

dffeas \pipe[2][32] (
	.clk(ctl_clk),
	.d(\pipe~146_combout ),
	.asdata(\pipe~21_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[2][32]~q ),
	.prn(vcc));
defparam \pipe[2][32] .is_wysiwyg = "true";
defparam \pipe[2][32] .power_up = "low";

arriaii_lcell_comb \pipe~21 (
	.dataa(!write_req),
	.datab(!pipefull_1),
	.datac(!pipefull_2),
	.datad(!\pipe[2][32]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~21 .extended_lut = "off";
defparam \pipe~21 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \pipe~21 .shared_arith = "off";

dffeas \pipe[1][32] (
	.clk(ctl_clk),
	.d(\pipe~21_combout ),
	.asdata(\pipe~4_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[1][32]~q ),
	.prn(vcc));
defparam \pipe[1][32] .is_wysiwyg = "true";
defparam \pipe[1][32] .power_up = "low";

arriaii_lcell_comb \pipe~4 (
	.dataa(!write_req),
	.datab(!pipefull_0),
	.datac(!pipefull_1),
	.datad(!\pipe[1][32]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~4 .extended_lut = "off";
defparam \pipe~4 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \pipe~4 .shared_arith = "off";

arriaii_lcell_comb \pipe~5 (
	.dataa(!pipe_12_3),
	.datab(!pipefull_2),
	.datac(!pipefull_3),
	.datad(!bank_addr_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~5 .extended_lut = "off";
defparam \pipe~5 .lut_mask = 64'h4575457545754575;
defparam \pipe~5 .shared_arith = "off";

arriaii_lcell_comb \pipe~6 (
	.dataa(!pipefull_1),
	.datab(!pipe_12_2),
	.datac(!pipefull_2),
	.datad(!bank_addr_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~6 .extended_lut = "off";
defparam \pipe~6 .lut_mask = 64'h2373237323732373;
defparam \pipe~6 .shared_arith = "off";

arriaii_lcell_comb \pipe~8 (
	.dataa(!pipefull_4),
	.datab(!pipefull_3),
	.datac(!pipe_12_4),
	.datad(!bank_addr_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~8 .extended_lut = "off";
defparam \pipe~8 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~8 .shared_arith = "off";

arriaii_lcell_comb \pipe~9 (
	.dataa(!pipe_10_3),
	.datab(!pipefull_2),
	.datac(!pipefull_3),
	.datad(!bank_addr_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~9 .extended_lut = "off";
defparam \pipe~9 .lut_mask = 64'h4575457545754575;
defparam \pipe~9 .shared_arith = "off";

arriaii_lcell_comb \pipe~10 (
	.dataa(!pipefull_1),
	.datab(!pipe_10_2),
	.datac(!pipefull_2),
	.datad(!bank_addr_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~10 .extended_lut = "off";
defparam \pipe~10 .lut_mask = 64'h2373237323732373;
defparam \pipe~10 .shared_arith = "off";

arriaii_lcell_comb \pipe~11 (
	.dataa(!pipefull_4),
	.datab(!pipefull_3),
	.datac(!pipe_10_4),
	.datad(!bank_addr_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~11 .extended_lut = "off";
defparam \pipe~11 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~11 .shared_arith = "off";

arriaii_lcell_comb \pipe~12 (
	.dataa(!pipe_11_3),
	.datab(!pipefull_2),
	.datac(!pipefull_3),
	.datad(!bank_addr_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~12 .extended_lut = "off";
defparam \pipe~12 .lut_mask = 64'h4575457545754575;
defparam \pipe~12 .shared_arith = "off";

arriaii_lcell_comb \pipe~13 (
	.dataa(!pipefull_1),
	.datab(!pipe_11_2),
	.datac(!pipefull_2),
	.datad(!bank_addr_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~13 .extended_lut = "off";
defparam \pipe~13 .lut_mask = 64'h2373237323732373;
defparam \pipe~13 .shared_arith = "off";

arriaii_lcell_comb \pipe~14 (
	.dataa(!pipefull_4),
	.datab(!pipefull_3),
	.datac(!pipe_11_4),
	.datad(!bank_addr_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~14 .extended_lut = "off";
defparam \pipe~14 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~14 .shared_arith = "off";

arriaii_lcell_comb \pipe~194 (
	.dataa(!size_1),
	.datab(!\pipe[7][29]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~194_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~194 .extended_lut = "off";
defparam \pipe~194 .lut_mask = 64'h1111111111111111;
defparam \pipe~194 .shared_arith = "off";

dffeas \pipe[7][29] (
	.clk(ctl_clk),
	.d(\pipe~194_combout ),
	.asdata(\pipe~182_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[7][29]~q ),
	.prn(vcc));
defparam \pipe[7][29] .is_wysiwyg = "true";
defparam \pipe[7][29] .power_up = "low";

arriaii_lcell_comb \pipe~182 (
	.dataa(!pipefull_7),
	.datab(!pipefull_6),
	.datac(!size_1),
	.datad(!\pipe[7][29]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~182_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~182 .extended_lut = "off";
defparam \pipe~182 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~182 .shared_arith = "off";

dffeas \pipe[6][29] (
	.clk(ctl_clk),
	.d(\pipe~182_combout ),
	.asdata(\pipe~170_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[6][29]~q ),
	.prn(vcc));
defparam \pipe[6][29] .is_wysiwyg = "true";
defparam \pipe[6][29] .power_up = "low";

arriaii_lcell_comb \pipe~170 (
	.dataa(!pipefull_6),
	.datab(!pipefull_5),
	.datac(!size_1),
	.datad(!\pipe[6][29]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~170_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~170 .extended_lut = "off";
defparam \pipe~170 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~170 .shared_arith = "off";

dffeas \pipe[5][29] (
	.clk(ctl_clk),
	.d(\pipe~170_combout ),
	.asdata(\pipe~158_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[5][29]~q ),
	.prn(vcc));
defparam \pipe[5][29] .is_wysiwyg = "true";
defparam \pipe[5][29] .power_up = "low";

arriaii_lcell_comb \pipe~158 (
	.dataa(!pipefull_5),
	.datab(!pipefull_4),
	.datac(!size_1),
	.datad(!\pipe[5][29]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~158_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~158 .extended_lut = "off";
defparam \pipe~158 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~158 .shared_arith = "off";

dffeas \pipe[4][29] (
	.clk(ctl_clk),
	.d(\pipe~158_combout ),
	.asdata(\pipe~153_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[4][29]~q ),
	.prn(vcc));
defparam \pipe[4][29] .is_wysiwyg = "true";
defparam \pipe[4][29] .power_up = "low";

arriaii_lcell_comb \pipe~153 (
	.dataa(!pipefull_4),
	.datab(!pipefull_3),
	.datac(!size_1),
	.datad(!\pipe[4][29]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~153_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~153 .extended_lut = "off";
defparam \pipe~153 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~153 .shared_arith = "off";

dffeas \pipe[3][29] (
	.clk(ctl_clk),
	.d(\pipe~153_combout ),
	.asdata(\pipe~148_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[3][29]~q ),
	.prn(vcc));
defparam \pipe[3][29] .is_wysiwyg = "true";
defparam \pipe[3][29] .power_up = "low";

arriaii_lcell_comb \pipe~148 (
	.dataa(!pipefull_2),
	.datab(!pipefull_3),
	.datac(!size_1),
	.datad(!\pipe[3][29]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~148_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~148 .extended_lut = "off";
defparam \pipe~148 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \pipe~148 .shared_arith = "off";

dffeas \pipe[2][29] (
	.clk(ctl_clk),
	.d(\pipe~148_combout ),
	.asdata(\pipe~143_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[2][29]~q ),
	.prn(vcc));
defparam \pipe[2][29] .is_wysiwyg = "true";
defparam \pipe[2][29] .power_up = "low";

arriaii_lcell_comb \pipe~143 (
	.dataa(!pipefull_1),
	.datab(!pipefull_2),
	.datac(!size_1),
	.datad(!\pipe[2][29]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~143_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~143 .extended_lut = "off";
defparam \pipe~143 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \pipe~143 .shared_arith = "off";

dffeas \pipe[1][29] (
	.clk(ctl_clk),
	.d(\pipe~143_combout ),
	.asdata(\pipe~15_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[1][29]~q ),
	.prn(vcc));
defparam \pipe[1][29] .is_wysiwyg = "true";
defparam \pipe[1][29] .power_up = "low";

arriaii_lcell_comb \pipe~15 (
	.dataa(!pipefull_0),
	.datab(!pipefull_1),
	.datac(!size_1),
	.datad(!\pipe[1][29]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~15 .extended_lut = "off";
defparam \pipe~15 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \pipe~15 .shared_arith = "off";

arriaii_lcell_comb \pipe~195 (
	.dataa(!size_0),
	.datab(!\pipe[7][28]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~195_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~195 .extended_lut = "off";
defparam \pipe~195 .lut_mask = 64'h1111111111111111;
defparam \pipe~195 .shared_arith = "off";

dffeas \pipe[7][28] (
	.clk(ctl_clk),
	.d(\pipe~195_combout ),
	.asdata(\pipe~183_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[7][28]~q ),
	.prn(vcc));
defparam \pipe[7][28] .is_wysiwyg = "true";
defparam \pipe[7][28] .power_up = "low";

arriaii_lcell_comb \pipe~183 (
	.dataa(!pipefull_7),
	.datab(!pipefull_6),
	.datac(!size_0),
	.datad(!\pipe[7][28]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~183_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~183 .extended_lut = "off";
defparam \pipe~183 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~183 .shared_arith = "off";

dffeas \pipe[6][28] (
	.clk(ctl_clk),
	.d(\pipe~183_combout ),
	.asdata(\pipe~171_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[6][28]~q ),
	.prn(vcc));
defparam \pipe[6][28] .is_wysiwyg = "true";
defparam \pipe[6][28] .power_up = "low";

arriaii_lcell_comb \pipe~171 (
	.dataa(!pipefull_6),
	.datab(!pipefull_5),
	.datac(!size_0),
	.datad(!\pipe[6][28]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~171_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~171 .extended_lut = "off";
defparam \pipe~171 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~171 .shared_arith = "off";

dffeas \pipe[5][28] (
	.clk(ctl_clk),
	.d(\pipe~171_combout ),
	.asdata(\pipe~159_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[5][28]~q ),
	.prn(vcc));
defparam \pipe[5][28] .is_wysiwyg = "true";
defparam \pipe[5][28] .power_up = "low";

arriaii_lcell_comb \pipe~159 (
	.dataa(!pipefull_5),
	.datab(!pipefull_4),
	.datac(!size_0),
	.datad(!\pipe[5][28]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~159_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~159 .extended_lut = "off";
defparam \pipe~159 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~159 .shared_arith = "off";

dffeas \pipe[4][28] (
	.clk(ctl_clk),
	.d(\pipe~159_combout ),
	.asdata(\pipe~154_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[4][28]~q ),
	.prn(vcc));
defparam \pipe[4][28] .is_wysiwyg = "true";
defparam \pipe[4][28] .power_up = "low";

arriaii_lcell_comb \pipe~154 (
	.dataa(!pipefull_4),
	.datab(!pipefull_3),
	.datac(!size_0),
	.datad(!\pipe[4][28]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~154_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~154 .extended_lut = "off";
defparam \pipe~154 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~154 .shared_arith = "off";

dffeas \pipe[3][28] (
	.clk(ctl_clk),
	.d(\pipe~154_combout ),
	.asdata(\pipe~149_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[3][28]~q ),
	.prn(vcc));
defparam \pipe[3][28] .is_wysiwyg = "true";
defparam \pipe[3][28] .power_up = "low";

arriaii_lcell_comb \pipe~149 (
	.dataa(!pipefull_2),
	.datab(!pipefull_3),
	.datac(!size_0),
	.datad(!\pipe[3][28]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~149_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~149 .extended_lut = "off";
defparam \pipe~149 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \pipe~149 .shared_arith = "off";

dffeas \pipe[2][28] (
	.clk(ctl_clk),
	.d(\pipe~149_combout ),
	.asdata(\pipe~144_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[2][28]~q ),
	.prn(vcc));
defparam \pipe[2][28] .is_wysiwyg = "true";
defparam \pipe[2][28] .power_up = "low";

arriaii_lcell_comb \pipe~144 (
	.dataa(!pipefull_1),
	.datab(!pipefull_2),
	.datac(!size_0),
	.datad(!\pipe[2][28]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~144_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~144 .extended_lut = "off";
defparam \pipe~144 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \pipe~144 .shared_arith = "off";

dffeas \pipe[1][28] (
	.clk(ctl_clk),
	.d(\pipe~144_combout ),
	.asdata(\pipe~16_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[1][28]~q ),
	.prn(vcc));
defparam \pipe[1][28] .is_wysiwyg = "true";
defparam \pipe[1][28] .power_up = "low";

arriaii_lcell_comb \pipe~16 (
	.dataa(!pipefull_0),
	.datab(!pipefull_1),
	.datac(!size_0),
	.datad(!\pipe[1][28]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~16 .extended_lut = "off";
defparam \pipe~16 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \pipe~16 .shared_arith = "off";

arriaii_lcell_comb \pipe~196 (
	.dataa(!read_req),
	.datab(!\pipe[7][33]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~196_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~196 .extended_lut = "off";
defparam \pipe~196 .lut_mask = 64'h1111111111111111;
defparam \pipe~196 .shared_arith = "off";

dffeas \pipe[7][33] (
	.clk(ctl_clk),
	.d(\pipe~196_combout ),
	.asdata(\pipe~184_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[7][33]~q ),
	.prn(vcc));
defparam \pipe[7][33] .is_wysiwyg = "true";
defparam \pipe[7][33] .power_up = "low";

arriaii_lcell_comb \pipe~184 (
	.dataa(!pipefull_7),
	.datab(!read_req),
	.datac(!pipefull_6),
	.datad(!\pipe[7][33]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~184_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~184 .extended_lut = "off";
defparam \pipe~184 .lut_mask = 64'h02F702F702F702F7;
defparam \pipe~184 .shared_arith = "off";

dffeas \pipe[6][33] (
	.clk(ctl_clk),
	.d(\pipe~184_combout ),
	.asdata(\pipe~172_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[6][33]~q ),
	.prn(vcc));
defparam \pipe[6][33] .is_wysiwyg = "true";
defparam \pipe[6][33] .power_up = "low";

arriaii_lcell_comb \pipe~172 (
	.dataa(!read_req),
	.datab(!pipefull_6),
	.datac(!pipefull_5),
	.datad(!\pipe[6][33]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~172_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~172 .extended_lut = "off";
defparam \pipe~172 .lut_mask = 64'h04F704F704F704F7;
defparam \pipe~172 .shared_arith = "off";

dffeas \pipe[5][33] (
	.clk(ctl_clk),
	.d(\pipe~172_combout ),
	.asdata(\pipe~160_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[5][33]~q ),
	.prn(vcc));
defparam \pipe[5][33] .is_wysiwyg = "true";
defparam \pipe[5][33] .power_up = "low";

arriaii_lcell_comb \pipe~160 (
	.dataa(!read_req),
	.datab(!pipefull_5),
	.datac(!pipefull_4),
	.datad(!\pipe[5][33]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~160_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~160 .extended_lut = "off";
defparam \pipe~160 .lut_mask = 64'h04F704F704F704F7;
defparam \pipe~160 .shared_arith = "off";

dffeas \pipe[4][33] (
	.clk(ctl_clk),
	.d(\pipe~160_combout ),
	.asdata(\pipe~155_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[4][33]~q ),
	.prn(vcc));
defparam \pipe[4][33] .is_wysiwyg = "true";
defparam \pipe[4][33] .power_up = "low";

arriaii_lcell_comb \pipe~155 (
	.dataa(!read_req),
	.datab(!pipefull_4),
	.datac(!pipefull_3),
	.datad(!\pipe[4][33]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~155_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~155 .extended_lut = "off";
defparam \pipe~155 .lut_mask = 64'h04F704F704F704F7;
defparam \pipe~155 .shared_arith = "off";

dffeas \pipe[3][33] (
	.clk(ctl_clk),
	.d(\pipe~155_combout ),
	.asdata(\pipe~150_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[3][33]~q ),
	.prn(vcc));
defparam \pipe[3][33] .is_wysiwyg = "true";
defparam \pipe[3][33] .power_up = "low";

arriaii_lcell_comb \pipe~150 (
	.dataa(!read_req),
	.datab(!pipefull_2),
	.datac(!pipefull_3),
	.datad(!\pipe[3][33]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~150_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~150 .extended_lut = "off";
defparam \pipe~150 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \pipe~150 .shared_arith = "off";

dffeas \pipe[2][33] (
	.clk(ctl_clk),
	.d(\pipe~150_combout ),
	.asdata(\pipe~145_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[2][33]~q ),
	.prn(vcc));
defparam \pipe[2][33] .is_wysiwyg = "true";
defparam \pipe[2][33] .power_up = "low";

arriaii_lcell_comb \pipe~145 (
	.dataa(!read_req),
	.datab(!pipefull_1),
	.datac(!pipefull_2),
	.datad(!\pipe[2][33]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~145_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~145 .extended_lut = "off";
defparam \pipe~145 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \pipe~145 .shared_arith = "off";

dffeas \pipe[1][33] (
	.clk(ctl_clk),
	.d(\pipe~145_combout ),
	.asdata(\pipe~17_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[1][33]~q ),
	.prn(vcc));
defparam \pipe[1][33] .is_wysiwyg = "true";
defparam \pipe[1][33] .power_up = "low";

arriaii_lcell_comb \pipe~17 (
	.dataa(!read_req),
	.datab(!pipefull_0),
	.datac(!pipefull_1),
	.datad(!\pipe[1][33]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~17 .extended_lut = "off";
defparam \pipe~17 .lut_mask = 64'h10DF10DF10DF10DF;
defparam \pipe~17 .shared_arith = "off";

arriaii_lcell_comb \pipe~18 (
	.dataa(!pipefull_5),
	.datab(!pipefull_4),
	.datac(!bank_addr_2),
	.datad(!pipe_12_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~18 .extended_lut = "off";
defparam \pipe~18 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~18 .shared_arith = "off";

arriaii_lcell_comb \pipe~19 (
	.dataa(!pipefull_5),
	.datab(!pipefull_4),
	.datac(!bank_addr_1),
	.datad(!pipe_11_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~19 .extended_lut = "off";
defparam \pipe~19 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~19 .shared_arith = "off";

arriaii_lcell_comb \pipe~20 (
	.dataa(!pipefull_5),
	.datab(!pipefull_4),
	.datac(!bank_addr_0),
	.datad(!pipe_10_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~20 .extended_lut = "off";
defparam \pipe~20 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~20 .shared_arith = "off";

arriaii_lcell_comb \pipe~22 (
	.dataa(!pipefull_6),
	.datab(!pipefull_5),
	.datac(!pipe_25_6),
	.datad(!row_addr_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~22 .extended_lut = "off";
defparam \pipe~22 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~22 .shared_arith = "off";

arriaii_lcell_comb \pipe~23 (
	.dataa(!pipefull_5),
	.datab(!pipefull_4),
	.datac(!pipe_25_5),
	.datad(!row_addr_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~23 .extended_lut = "off";
defparam \pipe~23 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~23 .shared_arith = "off";

arriaii_lcell_comb \pipe~24 (
	.dataa(!pipefull_0),
	.datab(!pipefull_1),
	.datac(!pipe_25_1),
	.datad(!row_addr_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~24 .extended_lut = "off";
defparam \pipe~24 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~24 .shared_arith = "off";

arriaii_lcell_comb \pipe~25 (
	.dataa(!pipefull_6),
	.datab(!pipefull_5),
	.datac(!pipe_26_6),
	.datad(!row_addr_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~25 .extended_lut = "off";
defparam \pipe~25 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~25 .shared_arith = "off";

arriaii_lcell_comb \pipe~26 (
	.dataa(!pipefull_5),
	.datab(!pipefull_4),
	.datac(!pipe_26_5),
	.datad(!row_addr_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~26 .extended_lut = "off";
defparam \pipe~26 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~26 .shared_arith = "off";

arriaii_lcell_comb \pipe~27 (
	.dataa(!pipefull_0),
	.datab(!pipefull_1),
	.datac(!pipe_26_1),
	.datad(!row_addr_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~27 .extended_lut = "off";
defparam \pipe~27 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~27 .shared_arith = "off";

arriaii_lcell_comb \pipe~28 (
	.dataa(!pipefull_6),
	.datab(!pipefull_5),
	.datac(!pipe_24_6),
	.datad(!row_addr_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~28 .extended_lut = "off";
defparam \pipe~28 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~28 .shared_arith = "off";

arriaii_lcell_comb \pipe~29 (
	.dataa(!pipefull_5),
	.datab(!pipefull_4),
	.datac(!pipe_24_5),
	.datad(!row_addr_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~29 .extended_lut = "off";
defparam \pipe~29 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~29 .shared_arith = "off";

arriaii_lcell_comb \pipe~30 (
	.dataa(!pipefull_0),
	.datab(!pipefull_1),
	.datac(!pipe_24_1),
	.datad(!row_addr_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~30 .extended_lut = "off";
defparam \pipe~30 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~30 .shared_arith = "off";

arriaii_lcell_comb \pipe~31 (
	.dataa(!pipefull_6),
	.datab(!pipefull_5),
	.datac(!pipe_22_6),
	.datad(!row_addr_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~31 .extended_lut = "off";
defparam \pipe~31 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~31 .shared_arith = "off";

arriaii_lcell_comb \pipe~32 (
	.dataa(!pipefull_5),
	.datab(!pipefull_4),
	.datac(!pipe_22_5),
	.datad(!row_addr_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~32 .extended_lut = "off";
defparam \pipe~32 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~32 .shared_arith = "off";

arriaii_lcell_comb \pipe~33 (
	.dataa(!pipefull_0),
	.datab(!pipefull_1),
	.datac(!pipe_22_1),
	.datad(!row_addr_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~33 .extended_lut = "off";
defparam \pipe~33 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~33 .shared_arith = "off";

arriaii_lcell_comb \pipe~34 (
	.dataa(!pipefull_6),
	.datab(!pipefull_5),
	.datac(!pipe_23_6),
	.datad(!row_addr_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~34 .extended_lut = "off";
defparam \pipe~34 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~34 .shared_arith = "off";

arriaii_lcell_comb \pipe~35 (
	.dataa(!pipefull_5),
	.datab(!pipefull_4),
	.datac(!pipe_23_5),
	.datad(!row_addr_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~35 .extended_lut = "off";
defparam \pipe~35 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~35 .shared_arith = "off";

arriaii_lcell_comb \pipe~36 (
	.dataa(!pipefull_0),
	.datab(!pipefull_1),
	.datac(!pipe_23_1),
	.datad(!row_addr_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~36 .extended_lut = "off";
defparam \pipe~36 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~36 .shared_arith = "off";

arriaii_lcell_comb \pipe~37 (
	.dataa(!pipefull_6),
	.datab(!pipefull_5),
	.datac(!pipe_21_6),
	.datad(!row_addr_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~37 .extended_lut = "off";
defparam \pipe~37 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~37 .shared_arith = "off";

arriaii_lcell_comb \pipe~38 (
	.dataa(!pipefull_5),
	.datab(!pipefull_4),
	.datac(!pipe_21_5),
	.datad(!row_addr_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~38 .extended_lut = "off";
defparam \pipe~38 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~38 .shared_arith = "off";

arriaii_lcell_comb \pipe~39 (
	.dataa(!pipefull_0),
	.datab(!pipefull_1),
	.datac(!pipe_21_1),
	.datad(!row_addr_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~39 .extended_lut = "off";
defparam \pipe~39 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~39 .shared_arith = "off";

arriaii_lcell_comb \pipe~40 (
	.dataa(!pipefull_6),
	.datab(!pipefull_5),
	.datac(!pipe_19_6),
	.datad(!row_addr_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~40 .extended_lut = "off";
defparam \pipe~40 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~40 .shared_arith = "off";

arriaii_lcell_comb \pipe~41 (
	.dataa(!pipefull_5),
	.datab(!pipefull_4),
	.datac(!pipe_19_5),
	.datad(!row_addr_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~41 .extended_lut = "off";
defparam \pipe~41 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~41 .shared_arith = "off";

arriaii_lcell_comb \pipe~42 (
	.dataa(!pipefull_0),
	.datab(!pipefull_1),
	.datac(!pipe_19_1),
	.datad(!row_addr_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~42 .extended_lut = "off";
defparam \pipe~42 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~42 .shared_arith = "off";

arriaii_lcell_comb \pipe~43 (
	.dataa(!pipefull_6),
	.datab(!pipefull_5),
	.datac(!pipe_20_6),
	.datad(!row_addr_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~43 .extended_lut = "off";
defparam \pipe~43 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~43 .shared_arith = "off";

arriaii_lcell_comb \pipe~44 (
	.dataa(!pipefull_5),
	.datab(!pipefull_4),
	.datac(!pipe_20_5),
	.datad(!row_addr_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~44 .extended_lut = "off";
defparam \pipe~44 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~44 .shared_arith = "off";

arriaii_lcell_comb \pipe~45 (
	.dataa(!pipefull_0),
	.datab(!pipefull_1),
	.datac(!pipe_20_1),
	.datad(!row_addr_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~45 .extended_lut = "off";
defparam \pipe~45 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~45 .shared_arith = "off";

arriaii_lcell_comb \pipe~46 (
	.dataa(!pipefull_6),
	.datab(!pipefull_5),
	.datac(!pipe_15_6),
	.datad(!row_addr_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~46 .extended_lut = "off";
defparam \pipe~46 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~46 .shared_arith = "off";

arriaii_lcell_comb \pipe~47 (
	.dataa(!pipefull_5),
	.datab(!pipefull_4),
	.datac(!pipe_15_5),
	.datad(!row_addr_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~47 .extended_lut = "off";
defparam \pipe~47 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~47 .shared_arith = "off";

arriaii_lcell_comb \pipe~48 (
	.dataa(!pipefull_0),
	.datab(!pipefull_1),
	.datac(!pipe_15_1),
	.datad(!row_addr_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~48 .extended_lut = "off";
defparam \pipe~48 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~48 .shared_arith = "off";

arriaii_lcell_comb \pipe~49 (
	.dataa(!pipefull_6),
	.datab(!pipefull_5),
	.datac(!pipe_13_6),
	.datad(!row_addr_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~49 .extended_lut = "off";
defparam \pipe~49 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~49 .shared_arith = "off";

arriaii_lcell_comb \pipe~50 (
	.dataa(!pipefull_5),
	.datab(!pipefull_4),
	.datac(!pipe_13_5),
	.datad(!row_addr_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~50_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~50 .extended_lut = "off";
defparam \pipe~50 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~50 .shared_arith = "off";

arriaii_lcell_comb \pipe~51 (
	.dataa(!pipefull_0),
	.datab(!pipefull_1),
	.datac(!pipe_13_1),
	.datad(!row_addr_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~51 .extended_lut = "off";
defparam \pipe~51 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~51 .shared_arith = "off";

arriaii_lcell_comb \pipe~52 (
	.dataa(!pipefull_6),
	.datab(!pipefull_5),
	.datac(!pipe_14_6),
	.datad(!row_addr_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~52 .extended_lut = "off";
defparam \pipe~52 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~52 .shared_arith = "off";

arriaii_lcell_comb \pipe~53 (
	.dataa(!pipefull_5),
	.datab(!pipefull_4),
	.datac(!pipe_14_5),
	.datad(!row_addr_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~53_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~53 .extended_lut = "off";
defparam \pipe~53 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~53 .shared_arith = "off";

arriaii_lcell_comb \pipe~54 (
	.dataa(!pipefull_0),
	.datab(!pipefull_1),
	.datac(!pipe_14_1),
	.datad(!row_addr_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~54_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~54 .extended_lut = "off";
defparam \pipe~54 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~54 .shared_arith = "off";

arriaii_lcell_comb \pipe~55 (
	.dataa(!pipefull_6),
	.datab(!pipefull_5),
	.datac(!pipe_18_6),
	.datad(!row_addr_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~55_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~55 .extended_lut = "off";
defparam \pipe~55 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~55 .shared_arith = "off";

arriaii_lcell_comb \pipe~56 (
	.dataa(!pipefull_5),
	.datab(!pipefull_4),
	.datac(!pipe_18_5),
	.datad(!row_addr_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~56_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~56 .extended_lut = "off";
defparam \pipe~56 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~56 .shared_arith = "off";

arriaii_lcell_comb \pipe~57 (
	.dataa(!pipefull_0),
	.datab(!pipefull_1),
	.datac(!pipe_18_1),
	.datad(!row_addr_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~57_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~57 .extended_lut = "off";
defparam \pipe~57 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~57 .shared_arith = "off";

arriaii_lcell_comb \pipe~58 (
	.dataa(!pipefull_6),
	.datab(!pipefull_5),
	.datac(!pipe_16_6),
	.datad(!row_addr_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~58_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~58 .extended_lut = "off";
defparam \pipe~58 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~58 .shared_arith = "off";

arriaii_lcell_comb \pipe~59 (
	.dataa(!pipefull_5),
	.datab(!pipefull_4),
	.datac(!pipe_16_5),
	.datad(!row_addr_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~59_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~59 .extended_lut = "off";
defparam \pipe~59 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~59 .shared_arith = "off";

arriaii_lcell_comb \pipe~60 (
	.dataa(!pipefull_0),
	.datab(!pipefull_1),
	.datac(!pipe_16_1),
	.datad(!row_addr_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~60_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~60 .extended_lut = "off";
defparam \pipe~60 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~60 .shared_arith = "off";

arriaii_lcell_comb \pipe~61 (
	.dataa(!pipefull_6),
	.datab(!pipefull_5),
	.datac(!pipe_17_6),
	.datad(!row_addr_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~61_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~61 .extended_lut = "off";
defparam \pipe~61 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~61 .shared_arith = "off";

arriaii_lcell_comb \pipe~62 (
	.dataa(!pipefull_5),
	.datab(!pipefull_4),
	.datac(!pipe_17_5),
	.datad(!row_addr_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~62_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~62 .extended_lut = "off";
defparam \pipe~62 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~62 .shared_arith = "off";

arriaii_lcell_comb \pipe~63 (
	.dataa(!pipefull_0),
	.datab(!pipefull_1),
	.datac(!pipe_17_1),
	.datad(!row_addr_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~63_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~63 .extended_lut = "off";
defparam \pipe~63 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~63 .shared_arith = "off";

arriaii_lcell_comb \pipe~64 (
	.dataa(!pipefull_6),
	.datab(!pipefull_5),
	.datac(!bank_addr_2),
	.datad(!pipe_12_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~64_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~64 .extended_lut = "off";
defparam \pipe~64 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~64 .shared_arith = "off";

arriaii_lcell_comb \pipe~65 (
	.dataa(!pipefull_6),
	.datab(!pipefull_5),
	.datac(!bank_addr_1),
	.datad(!pipe_11_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~65_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~65 .extended_lut = "off";
defparam \pipe~65 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~65 .shared_arith = "off";

arriaii_lcell_comb \pipe~66 (
	.dataa(!pipefull_6),
	.datab(!pipefull_5),
	.datac(!bank_addr_0),
	.datad(!pipe_10_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~66_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~66 .extended_lut = "off";
defparam \pipe~66 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~66 .shared_arith = "off";

arriaii_lcell_comb \pipe~67 (
	.dataa(!pipefull_4),
	.datab(!pipefull_3),
	.datac(!pipe_25_4),
	.datad(!row_addr_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~67_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~67 .extended_lut = "off";
defparam \pipe~67 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~67 .shared_arith = "off";

arriaii_lcell_comb \pipe~68 (
	.dataa(!pipefull_2),
	.datab(!pipefull_3),
	.datac(!pipe_25_3),
	.datad(!row_addr_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~68_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~68 .extended_lut = "off";
defparam \pipe~68 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~68 .shared_arith = "off";

arriaii_lcell_comb \pipe~69 (
	.dataa(!pipefull_4),
	.datab(!pipefull_3),
	.datac(!pipe_26_4),
	.datad(!row_addr_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~69_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~69 .extended_lut = "off";
defparam \pipe~69 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~69 .shared_arith = "off";

arriaii_lcell_comb \pipe~70 (
	.dataa(!pipefull_2),
	.datab(!pipefull_3),
	.datac(!pipe_26_3),
	.datad(!row_addr_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~70_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~70 .extended_lut = "off";
defparam \pipe~70 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~70 .shared_arith = "off";

arriaii_lcell_comb \pipe~71 (
	.dataa(!pipefull_4),
	.datab(!pipefull_3),
	.datac(!pipe_24_4),
	.datad(!row_addr_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~71_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~71 .extended_lut = "off";
defparam \pipe~71 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~71 .shared_arith = "off";

arriaii_lcell_comb \pipe~72 (
	.dataa(!pipefull_2),
	.datab(!pipefull_3),
	.datac(!pipe_24_3),
	.datad(!row_addr_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~72_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~72 .extended_lut = "off";
defparam \pipe~72 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~72 .shared_arith = "off";

arriaii_lcell_comb \pipe~73 (
	.dataa(!pipefull_4),
	.datab(!pipefull_3),
	.datac(!pipe_22_4),
	.datad(!row_addr_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~73_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~73 .extended_lut = "off";
defparam \pipe~73 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~73 .shared_arith = "off";

arriaii_lcell_comb \pipe~74 (
	.dataa(!pipefull_2),
	.datab(!pipefull_3),
	.datac(!pipe_22_3),
	.datad(!row_addr_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~74_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~74 .extended_lut = "off";
defparam \pipe~74 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~74 .shared_arith = "off";

arriaii_lcell_comb \pipe~75 (
	.dataa(!pipefull_4),
	.datab(!pipefull_3),
	.datac(!pipe_23_4),
	.datad(!row_addr_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~75_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~75 .extended_lut = "off";
defparam \pipe~75 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~75 .shared_arith = "off";

arriaii_lcell_comb \pipe~76 (
	.dataa(!pipefull_2),
	.datab(!pipefull_3),
	.datac(!pipe_23_3),
	.datad(!row_addr_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~76_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~76 .extended_lut = "off";
defparam \pipe~76 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~76 .shared_arith = "off";

arriaii_lcell_comb \pipe~77 (
	.dataa(!pipefull_4),
	.datab(!pipefull_3),
	.datac(!pipe_21_4),
	.datad(!row_addr_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~77_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~77 .extended_lut = "off";
defparam \pipe~77 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~77 .shared_arith = "off";

arriaii_lcell_comb \pipe~78 (
	.dataa(!pipefull_2),
	.datab(!pipefull_3),
	.datac(!pipe_21_3),
	.datad(!row_addr_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~78_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~78 .extended_lut = "off";
defparam \pipe~78 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~78 .shared_arith = "off";

arriaii_lcell_comb \pipe~79 (
	.dataa(!pipefull_4),
	.datab(!pipefull_3),
	.datac(!pipe_19_4),
	.datad(!row_addr_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~79_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~79 .extended_lut = "off";
defparam \pipe~79 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~79 .shared_arith = "off";

arriaii_lcell_comb \pipe~80 (
	.dataa(!pipefull_2),
	.datab(!pipefull_3),
	.datac(!pipe_19_3),
	.datad(!row_addr_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~80_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~80 .extended_lut = "off";
defparam \pipe~80 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~80 .shared_arith = "off";

arriaii_lcell_comb \pipe~81 (
	.dataa(!pipefull_4),
	.datab(!pipefull_3),
	.datac(!pipe_20_4),
	.datad(!row_addr_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~81_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~81 .extended_lut = "off";
defparam \pipe~81 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~81 .shared_arith = "off";

arriaii_lcell_comb \pipe~82 (
	.dataa(!pipefull_2),
	.datab(!pipefull_3),
	.datac(!pipe_20_3),
	.datad(!row_addr_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~82_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~82 .extended_lut = "off";
defparam \pipe~82 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~82 .shared_arith = "off";

arriaii_lcell_comb \pipe~83 (
	.dataa(!pipefull_4),
	.datab(!pipefull_3),
	.datac(!pipe_15_4),
	.datad(!row_addr_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~83_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~83 .extended_lut = "off";
defparam \pipe~83 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~83 .shared_arith = "off";

arriaii_lcell_comb \pipe~84 (
	.dataa(!pipefull_2),
	.datab(!pipefull_3),
	.datac(!pipe_15_3),
	.datad(!row_addr_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~84_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~84 .extended_lut = "off";
defparam \pipe~84 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~84 .shared_arith = "off";

arriaii_lcell_comb \pipe~85 (
	.dataa(!pipefull_4),
	.datab(!pipefull_3),
	.datac(!pipe_13_4),
	.datad(!row_addr_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~85_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~85 .extended_lut = "off";
defparam \pipe~85 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~85 .shared_arith = "off";

arriaii_lcell_comb \pipe~86 (
	.dataa(!pipefull_2),
	.datab(!pipefull_3),
	.datac(!pipe_13_3),
	.datad(!row_addr_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~86_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~86 .extended_lut = "off";
defparam \pipe~86 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~86 .shared_arith = "off";

arriaii_lcell_comb \pipe~87 (
	.dataa(!pipefull_4),
	.datab(!pipefull_3),
	.datac(!pipe_14_4),
	.datad(!row_addr_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~87_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~87 .extended_lut = "off";
defparam \pipe~87 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~87 .shared_arith = "off";

arriaii_lcell_comb \pipe~88 (
	.dataa(!pipefull_2),
	.datab(!pipefull_3),
	.datac(!pipe_14_3),
	.datad(!row_addr_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~88_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~88 .extended_lut = "off";
defparam \pipe~88 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~88 .shared_arith = "off";

arriaii_lcell_comb \pipe~89 (
	.dataa(!pipefull_4),
	.datab(!pipefull_3),
	.datac(!pipe_18_4),
	.datad(!row_addr_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~89_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~89 .extended_lut = "off";
defparam \pipe~89 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~89 .shared_arith = "off";

arriaii_lcell_comb \pipe~90 (
	.dataa(!pipefull_2),
	.datab(!pipefull_3),
	.datac(!pipe_18_3),
	.datad(!row_addr_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~90_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~90 .extended_lut = "off";
defparam \pipe~90 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~90 .shared_arith = "off";

arriaii_lcell_comb \pipe~91 (
	.dataa(!pipefull_4),
	.datab(!pipefull_3),
	.datac(!pipe_16_4),
	.datad(!row_addr_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~91_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~91 .extended_lut = "off";
defparam \pipe~91 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~91 .shared_arith = "off";

arriaii_lcell_comb \pipe~92 (
	.dataa(!pipefull_2),
	.datab(!pipefull_3),
	.datac(!pipe_16_3),
	.datad(!row_addr_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~92_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~92 .extended_lut = "off";
defparam \pipe~92 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~92 .shared_arith = "off";

arriaii_lcell_comb \pipe~93 (
	.dataa(!pipefull_4),
	.datab(!pipefull_3),
	.datac(!pipe_17_4),
	.datad(!row_addr_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~93_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~93 .extended_lut = "off";
defparam \pipe~93 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~93 .shared_arith = "off";

arriaii_lcell_comb \pipe~94 (
	.dataa(!pipefull_2),
	.datab(!pipefull_3),
	.datac(!pipe_17_3),
	.datad(!row_addr_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~94_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~94 .extended_lut = "off";
defparam \pipe~94 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~94 .shared_arith = "off";

arriaii_lcell_comb \pipe~95 (
	.dataa(!pipefull_7),
	.datab(!pipefull_6),
	.datac(!bank_addr_2),
	.datad(!pipe_12_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~95_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~95 .extended_lut = "off";
defparam \pipe~95 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~95 .shared_arith = "off";

arriaii_lcell_comb \pipe~96 (
	.dataa(!pipefull_7),
	.datab(!pipefull_6),
	.datac(!bank_addr_1),
	.datad(!pipe_11_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~96_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~96 .extended_lut = "off";
defparam \pipe~96 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~96 .shared_arith = "off";

arriaii_lcell_comb \pipe~97 (
	.dataa(!pipefull_7),
	.datab(!pipefull_6),
	.datac(!bank_addr_0),
	.datad(!pipe_10_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~97_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~97 .extended_lut = "off";
defparam \pipe~97 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~97 .shared_arith = "off";

arriaii_lcell_comb \pipe~98 (
	.dataa(!pipefull_7),
	.datab(!pipefull_6),
	.datac(!pipe_25_7),
	.datad(!row_addr_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~98_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~98 .extended_lut = "off";
defparam \pipe~98 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~98 .shared_arith = "off";

arriaii_lcell_comb \pipe~99 (
	.dataa(!pipefull_7),
	.datab(!pipefull_6),
	.datac(!pipe_26_7),
	.datad(!row_addr_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~99_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~99 .extended_lut = "off";
defparam \pipe~99 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~99 .shared_arith = "off";

arriaii_lcell_comb \pipe~100 (
	.dataa(!pipefull_7),
	.datab(!pipefull_6),
	.datac(!pipe_24_7),
	.datad(!row_addr_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~100_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~100 .extended_lut = "off";
defparam \pipe~100 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~100 .shared_arith = "off";

arriaii_lcell_comb \pipe~101 (
	.dataa(!pipefull_7),
	.datab(!pipefull_6),
	.datac(!pipe_22_7),
	.datad(!row_addr_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~101_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~101 .extended_lut = "off";
defparam \pipe~101 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~101 .shared_arith = "off";

arriaii_lcell_comb \pipe~102 (
	.dataa(!pipefull_7),
	.datab(!pipefull_6),
	.datac(!pipe_23_7),
	.datad(!row_addr_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~102_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~102 .extended_lut = "off";
defparam \pipe~102 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~102 .shared_arith = "off";

arriaii_lcell_comb \pipe~103 (
	.dataa(!pipefull_7),
	.datab(!pipefull_6),
	.datac(!pipe_21_7),
	.datad(!row_addr_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~103_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~103 .extended_lut = "off";
defparam \pipe~103 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~103 .shared_arith = "off";

arriaii_lcell_comb \pipe~104 (
	.dataa(!pipefull_7),
	.datab(!pipefull_6),
	.datac(!pipe_19_7),
	.datad(!row_addr_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~104_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~104 .extended_lut = "off";
defparam \pipe~104 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~104 .shared_arith = "off";

arriaii_lcell_comb \pipe~105 (
	.dataa(!pipefull_7),
	.datab(!pipefull_6),
	.datac(!pipe_20_7),
	.datad(!row_addr_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~105_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~105 .extended_lut = "off";
defparam \pipe~105 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~105 .shared_arith = "off";

arriaii_lcell_comb \pipe~106 (
	.dataa(!pipefull_7),
	.datab(!pipefull_6),
	.datac(!pipe_15_7),
	.datad(!row_addr_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~106_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~106 .extended_lut = "off";
defparam \pipe~106 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~106 .shared_arith = "off";

arriaii_lcell_comb \pipe~107 (
	.dataa(!pipefull_7),
	.datab(!pipefull_6),
	.datac(!pipe_13_7),
	.datad(!row_addr_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~107_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~107 .extended_lut = "off";
defparam \pipe~107 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~107 .shared_arith = "off";

arriaii_lcell_comb \pipe~108 (
	.dataa(!pipefull_7),
	.datab(!pipefull_6),
	.datac(!pipe_14_7),
	.datad(!row_addr_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~108_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~108 .extended_lut = "off";
defparam \pipe~108 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~108 .shared_arith = "off";

arriaii_lcell_comb \pipe~109 (
	.dataa(!pipefull_7),
	.datab(!pipefull_6),
	.datac(!pipe_18_7),
	.datad(!row_addr_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~109_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~109 .extended_lut = "off";
defparam \pipe~109 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~109 .shared_arith = "off";

arriaii_lcell_comb \pipe~110 (
	.dataa(!pipefull_7),
	.datab(!pipefull_6),
	.datac(!pipe_16_7),
	.datad(!row_addr_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~110_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~110 .extended_lut = "off";
defparam \pipe~110 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~110 .shared_arith = "off";

arriaii_lcell_comb \pipe~111 (
	.dataa(!pipefull_7),
	.datab(!pipefull_6),
	.datac(!pipe_17_7),
	.datad(!row_addr_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~111_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~111 .extended_lut = "off";
defparam \pipe~111 .lut_mask = 64'h0D2F0D2F0D2F0D2F;
defparam \pipe~111 .shared_arith = "off";

arriaii_lcell_comb \pipe~112 (
	.dataa(!generating),
	.datab(!pipe_26_7),
	.datac(!buf_row_addr_13),
	.datad(!local_address_24),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~112_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~112 .extended_lut = "off";
defparam \pipe~112 .lut_mask = 64'h0123012301230123;
defparam \pipe~112 .shared_arith = "off";

arriaii_lcell_comb \pipe~113 (
	.dataa(!generating),
	.datab(!pipe_24_7),
	.datac(!buf_row_addr_11),
	.datad(!local_address_22),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~113_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~113 .extended_lut = "off";
defparam \pipe~113 .lut_mask = 64'h0123012301230123;
defparam \pipe~113 .shared_arith = "off";

arriaii_lcell_comb \pipe~114 (
	.dataa(!generating),
	.datab(!pipe_25_7),
	.datac(!buf_row_addr_12),
	.datad(!local_address_23),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~114_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~114 .extended_lut = "off";
defparam \pipe~114 .lut_mask = 64'h0123012301230123;
defparam \pipe~114 .shared_arith = "off";

arriaii_lcell_comb \pipe~115 (
	.dataa(!generating),
	.datab(!pipe_23_7),
	.datac(!buf_row_addr_10),
	.datad(!local_address_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~115_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~115 .extended_lut = "off";
defparam \pipe~115 .lut_mask = 64'h0123012301230123;
defparam \pipe~115 .shared_arith = "off";

arriaii_lcell_comb \pipe~116 (
	.dataa(!generating),
	.datab(!pipe_21_7),
	.datac(!buf_row_addr_8),
	.datad(!local_address_19),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~116_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~116 .extended_lut = "off";
defparam \pipe~116 .lut_mask = 64'h0123012301230123;
defparam \pipe~116 .shared_arith = "off";

arriaii_lcell_comb \pipe~117 (
	.dataa(!generating),
	.datab(!pipe_22_7),
	.datac(!buf_row_addr_9),
	.datad(!local_address_20),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~117_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~117 .extended_lut = "off";
defparam \pipe~117 .lut_mask = 64'h0123012301230123;
defparam \pipe~117 .shared_arith = "off";

arriaii_lcell_comb \pipe~118 (
	.dataa(!generating),
	.datab(!pipe_20_7),
	.datac(!buf_row_addr_7),
	.datad(!local_address_18),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~118_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~118 .extended_lut = "off";
defparam \pipe~118 .lut_mask = 64'h0123012301230123;
defparam \pipe~118 .shared_arith = "off";

arriaii_lcell_comb \pipe~119 (
	.dataa(!generating),
	.datab(!pipe_18_7),
	.datac(!buf_row_addr_5),
	.datad(!local_address_16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~119_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~119 .extended_lut = "off";
defparam \pipe~119 .lut_mask = 64'h0123012301230123;
defparam \pipe~119 .shared_arith = "off";

arriaii_lcell_comb \pipe~120 (
	.dataa(!generating),
	.datab(!pipe_19_7),
	.datac(!buf_row_addr_6),
	.datad(!local_address_17),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~120_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~120 .extended_lut = "off";
defparam \pipe~120 .lut_mask = 64'h0123012301230123;
defparam \pipe~120 .shared_arith = "off";

arriaii_lcell_comb \pipe~121 (
	.dataa(!generating),
	.datab(!pipe_17_7),
	.datac(!buf_row_addr_4),
	.datad(!local_address_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~121_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~121 .extended_lut = "off";
defparam \pipe~121 .lut_mask = 64'h0123012301230123;
defparam \pipe~121 .shared_arith = "off";

arriaii_lcell_comb \pipe~122 (
	.dataa(!generating),
	.datab(!pipe_15_7),
	.datac(!buf_row_addr_2),
	.datad(!local_address_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~122_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~122 .extended_lut = "off";
defparam \pipe~122 .lut_mask = 64'h0123012301230123;
defparam \pipe~122 .shared_arith = "off";

arriaii_lcell_comb \pipe~123 (
	.dataa(!generating),
	.datab(!pipe_16_7),
	.datac(!buf_row_addr_3),
	.datad(!local_address_14),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~123_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~123 .extended_lut = "off";
defparam \pipe~123 .lut_mask = 64'h0123012301230123;
defparam \pipe~123 .shared_arith = "off";

arriaii_lcell_comb \pipe~124 (
	.dataa(!generating),
	.datab(!buf_bank_addr_1),
	.datac(!local_address_9),
	.datad(!pipe_11_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~124_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~124 .extended_lut = "off";
defparam \pipe~124 .lut_mask = 64'h001B001B001B001B;
defparam \pipe~124 .shared_arith = "off";

arriaii_lcell_comb \pipe~125 (
	.dataa(!generating),
	.datab(!buf_bank_addr_0),
	.datac(!local_address_8),
	.datad(!pipe_10_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~125_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~125 .extended_lut = "off";
defparam \pipe~125 .lut_mask = 64'h001B001B001B001B;
defparam \pipe~125 .shared_arith = "off";

arriaii_lcell_comb \pipe~126 (
	.dataa(!generating),
	.datab(!pipe_14_7),
	.datac(!buf_row_addr_1),
	.datad(!local_address_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~126_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~126 .extended_lut = "off";
defparam \pipe~126 .lut_mask = 64'h0123012301230123;
defparam \pipe~126 .shared_arith = "off";

arriaii_lcell_comb \pipe~127 (
	.dataa(!generating),
	.datab(!buf_bank_addr_2),
	.datac(!local_address_10),
	.datad(!pipe_12_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~127_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~127 .extended_lut = "off";
defparam \pipe~127 .lut_mask = 64'h001B001B001B001B;
defparam \pipe~127 .shared_arith = "off";

arriaii_lcell_comb \pipe~128 (
	.dataa(!generating),
	.datab(!pipe_13_7),
	.datac(!buf_row_addr_0),
	.datad(!local_address_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~128_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~128 .extended_lut = "off";
defparam \pipe~128 .lut_mask = 64'h0123012301230123;
defparam \pipe~128 .shared_arith = "off";

arriaii_lcell_comb \pipe~129 (
	.dataa(!pipefull_1),
	.datab(!pipefull_2),
	.datac(!pipe_25_2),
	.datad(!row_addr_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~129_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~129 .extended_lut = "off";
defparam \pipe~129 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~129 .shared_arith = "off";

arriaii_lcell_comb \pipe~130 (
	.dataa(!pipefull_1),
	.datab(!pipefull_2),
	.datac(!pipe_26_2),
	.datad(!row_addr_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~130_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~130 .extended_lut = "off";
defparam \pipe~130 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~130 .shared_arith = "off";

arriaii_lcell_comb \pipe~131 (
	.dataa(!pipefull_1),
	.datab(!pipefull_2),
	.datac(!pipe_24_2),
	.datad(!row_addr_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~131_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~131 .extended_lut = "off";
defparam \pipe~131 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~131 .shared_arith = "off";

arriaii_lcell_comb \pipe~132 (
	.dataa(!pipefull_1),
	.datab(!pipefull_2),
	.datac(!pipe_22_2),
	.datad(!row_addr_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~132_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~132 .extended_lut = "off";
defparam \pipe~132 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~132 .shared_arith = "off";

arriaii_lcell_comb \pipe~133 (
	.dataa(!pipefull_1),
	.datab(!pipefull_2),
	.datac(!pipe_23_2),
	.datad(!row_addr_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~133_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~133 .extended_lut = "off";
defparam \pipe~133 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~133 .shared_arith = "off";

arriaii_lcell_comb \pipe~134 (
	.dataa(!pipefull_1),
	.datab(!pipefull_2),
	.datac(!pipe_21_2),
	.datad(!row_addr_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~134_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~134 .extended_lut = "off";
defparam \pipe~134 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~134 .shared_arith = "off";

arriaii_lcell_comb \pipe~135 (
	.dataa(!pipefull_1),
	.datab(!pipefull_2),
	.datac(!pipe_19_2),
	.datad(!row_addr_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~135_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~135 .extended_lut = "off";
defparam \pipe~135 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~135 .shared_arith = "off";

arriaii_lcell_comb \pipe~136 (
	.dataa(!pipefull_1),
	.datab(!pipefull_2),
	.datac(!pipe_20_2),
	.datad(!row_addr_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~136_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~136 .extended_lut = "off";
defparam \pipe~136 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~136 .shared_arith = "off";

arriaii_lcell_comb \pipe~137 (
	.dataa(!pipefull_1),
	.datab(!pipefull_2),
	.datac(!pipe_15_2),
	.datad(!row_addr_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~137_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~137 .extended_lut = "off";
defparam \pipe~137 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~137 .shared_arith = "off";

arriaii_lcell_comb \pipe~138 (
	.dataa(!pipefull_1),
	.datab(!pipefull_2),
	.datac(!pipe_13_2),
	.datad(!row_addr_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~138_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~138 .extended_lut = "off";
defparam \pipe~138 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~138 .shared_arith = "off";

arriaii_lcell_comb \pipe~139 (
	.dataa(!pipefull_1),
	.datab(!pipefull_2),
	.datac(!pipe_14_2),
	.datad(!row_addr_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~139_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~139 .extended_lut = "off";
defparam \pipe~139 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~139 .shared_arith = "off";

arriaii_lcell_comb \pipe~140 (
	.dataa(!pipefull_1),
	.datab(!pipefull_2),
	.datac(!pipe_18_2),
	.datad(!row_addr_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~140_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~140 .extended_lut = "off";
defparam \pipe~140 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~140 .shared_arith = "off";

arriaii_lcell_comb \pipe~141 (
	.dataa(!pipefull_1),
	.datab(!pipefull_2),
	.datac(!pipe_16_2),
	.datad(!row_addr_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~141_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~141 .extended_lut = "off";
defparam \pipe~141 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~141 .shared_arith = "off";

arriaii_lcell_comb \pipe~142 (
	.dataa(!pipefull_1),
	.datab(!pipefull_2),
	.datac(!pipe_17_2),
	.datad(!row_addr_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~142_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~142 .extended_lut = "off";
defparam \pipe~142 .lut_mask = 64'h0B4F0B4F0B4F0B4F;
defparam \pipe~142 .shared_arith = "off";

arriaii_lcell_comb \pipe~212 (
	.dataa(!local_address_0),
	.datab(!generating),
	.datac(!\pipe[7][2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~212_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~212 .extended_lut = "off";
defparam \pipe~212 .lut_mask = 64'h0404040404040404;
defparam \pipe~212 .shared_arith = "off";

dffeas \pipe[7][2] (
	.clk(ctl_clk),
	.d(\pipe~212_combout ),
	.asdata(\pipe~204_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[7][2]~q ),
	.prn(vcc));
defparam \pipe[7][2] .is_wysiwyg = "true";
defparam \pipe[7][2] .power_up = "low";

arriaii_lcell_comb \pipe~204 (
	.dataa(!pipefull_7),
	.datab(!pipefull_6),
	.datac(!col_addr_2),
	.datad(!\pipe[7][2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~204_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~204 .extended_lut = "off";
defparam \pipe~204 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~204 .shared_arith = "off";

dffeas \pipe[6][2] (
	.clk(ctl_clk),
	.d(\pipe~204_combout ),
	.asdata(\pipe~193_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[6][2]~q ),
	.prn(vcc));
defparam \pipe[6][2] .is_wysiwyg = "true";
defparam \pipe[6][2] .power_up = "low";

arriaii_lcell_comb \pipe~193 (
	.dataa(!pipefull_6),
	.datab(!pipefull_5),
	.datac(!col_addr_2),
	.datad(!\pipe[6][2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~193_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~193 .extended_lut = "off";
defparam \pipe~193 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~193 .shared_arith = "off";

dffeas \pipe[5][2] (
	.clk(ctl_clk),
	.d(\pipe~193_combout ),
	.asdata(\pipe~181_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[5][2]~q ),
	.prn(vcc));
defparam \pipe[5][2] .is_wysiwyg = "true";
defparam \pipe[5][2] .power_up = "low";

arriaii_lcell_comb \pipe~181 (
	.dataa(!pipefull_5),
	.datab(!pipefull_4),
	.datac(!col_addr_2),
	.datad(!\pipe[5][2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~181_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~181 .extended_lut = "off";
defparam \pipe~181 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~181 .shared_arith = "off";

dffeas \pipe[4][2] (
	.clk(ctl_clk),
	.d(\pipe~181_combout ),
	.asdata(\pipe~169_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[4][2]~q ),
	.prn(vcc));
defparam \pipe[4][2] .is_wysiwyg = "true";
defparam \pipe[4][2] .power_up = "low";

arriaii_lcell_comb \pipe~169 (
	.dataa(!pipefull_4),
	.datab(!pipefull_3),
	.datac(!col_addr_2),
	.datad(!\pipe[4][2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~169_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~169 .extended_lut = "off";
defparam \pipe~169 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~169 .shared_arith = "off";

dffeas \pipe[3][2] (
	.clk(ctl_clk),
	.d(\pipe~169_combout ),
	.asdata(\pipe~157_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[3][2]~q ),
	.prn(vcc));
defparam \pipe[3][2] .is_wysiwyg = "true";
defparam \pipe[3][2] .power_up = "low";

arriaii_lcell_comb \pipe~157 (
	.dataa(!pipefull_2),
	.datab(!pipefull_3),
	.datac(!col_addr_2),
	.datad(!\pipe[3][2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~157_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~157 .extended_lut = "off";
defparam \pipe~157 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \pipe~157 .shared_arith = "off";

dffeas \pipe[2][2] (
	.clk(ctl_clk),
	.d(\pipe~157_combout ),
	.asdata(\pipe~152_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[2][2]~q ),
	.prn(vcc));
defparam \pipe[2][2] .is_wysiwyg = "true";
defparam \pipe[2][2] .power_up = "low";

arriaii_lcell_comb \pipe~152 (
	.dataa(!pipefull_1),
	.datab(!pipefull_2),
	.datac(!col_addr_2),
	.datad(!\pipe[2][2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~152_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~152 .extended_lut = "off";
defparam \pipe~152 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \pipe~152 .shared_arith = "off";

dffeas \pipe[1][2] (
	.clk(ctl_clk),
	.d(\pipe~152_combout ),
	.asdata(\pipe~147_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[1][2]~q ),
	.prn(vcc));
defparam \pipe[1][2] .is_wysiwyg = "true";
defparam \pipe[1][2] .power_up = "low";

arriaii_lcell_comb \pipe~147 (
	.dataa(!pipefull_0),
	.datab(!pipefull_1),
	.datac(!col_addr_2),
	.datad(!\pipe[1][2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~147_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~147 .extended_lut = "off";
defparam \pipe~147 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \pipe~147 .shared_arith = "off";

arriaii_lcell_comb \pipe~227 (
	.dataa(!generating),
	.datab(!buf_col_addr_3),
	.datac(!local_address_1),
	.datad(!\pipe[7][3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~227_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~227 .extended_lut = "off";
defparam \pipe~227 .lut_mask = 64'h001B001B001B001B;
defparam \pipe~227 .shared_arith = "off";

dffeas \pipe[7][3] (
	.clk(ctl_clk),
	.d(\pipe~227_combout ),
	.asdata(\pipe~220_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[7][3]~q ),
	.prn(vcc));
defparam \pipe[7][3] .is_wysiwyg = "true";
defparam \pipe[7][3] .power_up = "low";

arriaii_lcell_comb \pipe~220 (
	.dataa(!pipefull_7),
	.datab(!pipefull_6),
	.datac(!col_addr_3),
	.datad(!\pipe[7][3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~220_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~220 .extended_lut = "off";
defparam \pipe~220 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~220 .shared_arith = "off";

dffeas \pipe[6][3] (
	.clk(ctl_clk),
	.d(\pipe~220_combout ),
	.asdata(\pipe~213_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[6][3]~q ),
	.prn(vcc));
defparam \pipe[6][3] .is_wysiwyg = "true";
defparam \pipe[6][3] .power_up = "low";

arriaii_lcell_comb \pipe~213 (
	.dataa(!pipefull_6),
	.datab(!pipefull_5),
	.datac(!col_addr_3),
	.datad(!\pipe[6][3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~213_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~213 .extended_lut = "off";
defparam \pipe~213 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~213 .shared_arith = "off";

dffeas \pipe[5][3] (
	.clk(ctl_clk),
	.d(\pipe~213_combout ),
	.asdata(\pipe~205_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[5][3]~q ),
	.prn(vcc));
defparam \pipe[5][3] .is_wysiwyg = "true";
defparam \pipe[5][3] .power_up = "low";

arriaii_lcell_comb \pipe~205 (
	.dataa(!pipefull_5),
	.datab(!pipefull_4),
	.datac(!col_addr_3),
	.datad(!\pipe[5][3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~205_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~205 .extended_lut = "off";
defparam \pipe~205 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~205 .shared_arith = "off";

dffeas \pipe[4][3] (
	.clk(ctl_clk),
	.d(\pipe~205_combout ),
	.asdata(\pipe~197_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[4][3]~q ),
	.prn(vcc));
defparam \pipe[4][3] .is_wysiwyg = "true";
defparam \pipe[4][3] .power_up = "low";

arriaii_lcell_comb \pipe~197 (
	.dataa(!pipefull_4),
	.datab(!pipefull_3),
	.datac(!col_addr_3),
	.datad(!\pipe[4][3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~197_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~197 .extended_lut = "off";
defparam \pipe~197 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~197 .shared_arith = "off";

dffeas \pipe[3][3] (
	.clk(ctl_clk),
	.d(\pipe~197_combout ),
	.asdata(\pipe~185_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[3][3]~q ),
	.prn(vcc));
defparam \pipe[3][3] .is_wysiwyg = "true";
defparam \pipe[3][3] .power_up = "low";

arriaii_lcell_comb \pipe~185 (
	.dataa(!pipefull_2),
	.datab(!pipefull_3),
	.datac(!col_addr_3),
	.datad(!\pipe[3][3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~185_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~185 .extended_lut = "off";
defparam \pipe~185 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \pipe~185 .shared_arith = "off";

dffeas \pipe[2][3] (
	.clk(ctl_clk),
	.d(\pipe~185_combout ),
	.asdata(\pipe~173_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[2][3]~q ),
	.prn(vcc));
defparam \pipe[2][3] .is_wysiwyg = "true";
defparam \pipe[2][3] .power_up = "low";

arriaii_lcell_comb \pipe~173 (
	.dataa(!pipefull_1),
	.datab(!pipefull_2),
	.datac(!col_addr_3),
	.datad(!\pipe[2][3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~173_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~173 .extended_lut = "off";
defparam \pipe~173 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \pipe~173 .shared_arith = "off";

dffeas \pipe[1][3] (
	.clk(ctl_clk),
	.d(\pipe~173_combout ),
	.asdata(\pipe~161_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[1][3]~q ),
	.prn(vcc));
defparam \pipe[1][3] .is_wysiwyg = "true";
defparam \pipe[1][3] .power_up = "low";

arriaii_lcell_comb \pipe~161 (
	.dataa(!pipefull_0),
	.datab(!pipefull_1),
	.datac(!col_addr_3),
	.datad(!\pipe[1][3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~161_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~161 .extended_lut = "off";
defparam \pipe~161 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \pipe~161 .shared_arith = "off";

arriaii_lcell_comb \pipe~228 (
	.dataa(!generating),
	.datab(!buf_col_addr_4),
	.datac(!local_address_2),
	.datad(!\pipe[7][4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~228_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~228 .extended_lut = "off";
defparam \pipe~228 .lut_mask = 64'h001B001B001B001B;
defparam \pipe~228 .shared_arith = "off";

dffeas \pipe[7][4] (
	.clk(ctl_clk),
	.d(\pipe~228_combout ),
	.asdata(\pipe~221_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[7][4]~q ),
	.prn(vcc));
defparam \pipe[7][4] .is_wysiwyg = "true";
defparam \pipe[7][4] .power_up = "low";

arriaii_lcell_comb \pipe~221 (
	.dataa(!pipefull_7),
	.datab(!pipefull_6),
	.datac(!col_addr_4),
	.datad(!\pipe[7][4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~221_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~221 .extended_lut = "off";
defparam \pipe~221 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~221 .shared_arith = "off";

dffeas \pipe[6][4] (
	.clk(ctl_clk),
	.d(\pipe~221_combout ),
	.asdata(\pipe~214_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[6][4]~q ),
	.prn(vcc));
defparam \pipe[6][4] .is_wysiwyg = "true";
defparam \pipe[6][4] .power_up = "low";

arriaii_lcell_comb \pipe~214 (
	.dataa(!pipefull_6),
	.datab(!pipefull_5),
	.datac(!col_addr_4),
	.datad(!\pipe[6][4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~214_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~214 .extended_lut = "off";
defparam \pipe~214 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~214 .shared_arith = "off";

dffeas \pipe[5][4] (
	.clk(ctl_clk),
	.d(\pipe~214_combout ),
	.asdata(\pipe~206_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[5][4]~q ),
	.prn(vcc));
defparam \pipe[5][4] .is_wysiwyg = "true";
defparam \pipe[5][4] .power_up = "low";

arriaii_lcell_comb \pipe~206 (
	.dataa(!pipefull_5),
	.datab(!pipefull_4),
	.datac(!col_addr_4),
	.datad(!\pipe[5][4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~206_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~206 .extended_lut = "off";
defparam \pipe~206 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~206 .shared_arith = "off";

dffeas \pipe[4][4] (
	.clk(ctl_clk),
	.d(\pipe~206_combout ),
	.asdata(\pipe~198_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[4][4]~q ),
	.prn(vcc));
defparam \pipe[4][4] .is_wysiwyg = "true";
defparam \pipe[4][4] .power_up = "low";

arriaii_lcell_comb \pipe~198 (
	.dataa(!pipefull_4),
	.datab(!pipefull_3),
	.datac(!col_addr_4),
	.datad(!\pipe[4][4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~198_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~198 .extended_lut = "off";
defparam \pipe~198 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~198 .shared_arith = "off";

dffeas \pipe[3][4] (
	.clk(ctl_clk),
	.d(\pipe~198_combout ),
	.asdata(\pipe~186_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[3][4]~q ),
	.prn(vcc));
defparam \pipe[3][4] .is_wysiwyg = "true";
defparam \pipe[3][4] .power_up = "low";

arriaii_lcell_comb \pipe~186 (
	.dataa(!pipefull_2),
	.datab(!pipefull_3),
	.datac(!col_addr_4),
	.datad(!\pipe[3][4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~186_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~186 .extended_lut = "off";
defparam \pipe~186 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \pipe~186 .shared_arith = "off";

dffeas \pipe[2][4] (
	.clk(ctl_clk),
	.d(\pipe~186_combout ),
	.asdata(\pipe~174_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[2][4]~q ),
	.prn(vcc));
defparam \pipe[2][4] .is_wysiwyg = "true";
defparam \pipe[2][4] .power_up = "low";

arriaii_lcell_comb \pipe~174 (
	.dataa(!pipefull_1),
	.datab(!pipefull_2),
	.datac(!col_addr_4),
	.datad(!\pipe[2][4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~174_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~174 .extended_lut = "off";
defparam \pipe~174 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \pipe~174 .shared_arith = "off";

dffeas \pipe[1][4] (
	.clk(ctl_clk),
	.d(\pipe~174_combout ),
	.asdata(\pipe~162_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[1][4]~q ),
	.prn(vcc));
defparam \pipe[1][4] .is_wysiwyg = "true";
defparam \pipe[1][4] .power_up = "low";

arriaii_lcell_comb \pipe~162 (
	.dataa(!pipefull_0),
	.datab(!pipefull_1),
	.datac(!col_addr_4),
	.datad(!\pipe[1][4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~162_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~162 .extended_lut = "off";
defparam \pipe~162 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \pipe~162 .shared_arith = "off";

arriaii_lcell_comb \pipe~229 (
	.dataa(!generating),
	.datab(!buf_col_addr_5),
	.datac(!local_address_3),
	.datad(!\pipe[7][5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~229_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~229 .extended_lut = "off";
defparam \pipe~229 .lut_mask = 64'h001B001B001B001B;
defparam \pipe~229 .shared_arith = "off";

dffeas \pipe[7][5] (
	.clk(ctl_clk),
	.d(\pipe~229_combout ),
	.asdata(\pipe~222_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[7][5]~q ),
	.prn(vcc));
defparam \pipe[7][5] .is_wysiwyg = "true";
defparam \pipe[7][5] .power_up = "low";

arriaii_lcell_comb \pipe~222 (
	.dataa(!pipefull_7),
	.datab(!pipefull_6),
	.datac(!col_addr_5),
	.datad(!\pipe[7][5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~222_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~222 .extended_lut = "off";
defparam \pipe~222 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~222 .shared_arith = "off";

dffeas \pipe[6][5] (
	.clk(ctl_clk),
	.d(\pipe~222_combout ),
	.asdata(\pipe~215_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[6][5]~q ),
	.prn(vcc));
defparam \pipe[6][5] .is_wysiwyg = "true";
defparam \pipe[6][5] .power_up = "low";

arriaii_lcell_comb \pipe~215 (
	.dataa(!pipefull_6),
	.datab(!pipefull_5),
	.datac(!col_addr_5),
	.datad(!\pipe[6][5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~215_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~215 .extended_lut = "off";
defparam \pipe~215 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~215 .shared_arith = "off";

dffeas \pipe[5][5] (
	.clk(ctl_clk),
	.d(\pipe~215_combout ),
	.asdata(\pipe~207_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[5][5]~q ),
	.prn(vcc));
defparam \pipe[5][5] .is_wysiwyg = "true";
defparam \pipe[5][5] .power_up = "low";

arriaii_lcell_comb \pipe~207 (
	.dataa(!pipefull_5),
	.datab(!pipefull_4),
	.datac(!col_addr_5),
	.datad(!\pipe[5][5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~207_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~207 .extended_lut = "off";
defparam \pipe~207 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~207 .shared_arith = "off";

dffeas \pipe[4][5] (
	.clk(ctl_clk),
	.d(\pipe~207_combout ),
	.asdata(\pipe~199_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[4][5]~q ),
	.prn(vcc));
defparam \pipe[4][5] .is_wysiwyg = "true";
defparam \pipe[4][5] .power_up = "low";

arriaii_lcell_comb \pipe~199 (
	.dataa(!pipefull_4),
	.datab(!pipefull_3),
	.datac(!col_addr_5),
	.datad(!\pipe[4][5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~199_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~199 .extended_lut = "off";
defparam \pipe~199 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~199 .shared_arith = "off";

dffeas \pipe[3][5] (
	.clk(ctl_clk),
	.d(\pipe~199_combout ),
	.asdata(\pipe~187_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[3][5]~q ),
	.prn(vcc));
defparam \pipe[3][5] .is_wysiwyg = "true";
defparam \pipe[3][5] .power_up = "low";

arriaii_lcell_comb \pipe~187 (
	.dataa(!pipefull_2),
	.datab(!pipefull_3),
	.datac(!col_addr_5),
	.datad(!\pipe[3][5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~187_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~187 .extended_lut = "off";
defparam \pipe~187 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \pipe~187 .shared_arith = "off";

dffeas \pipe[2][5] (
	.clk(ctl_clk),
	.d(\pipe~187_combout ),
	.asdata(\pipe~175_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[2][5]~q ),
	.prn(vcc));
defparam \pipe[2][5] .is_wysiwyg = "true";
defparam \pipe[2][5] .power_up = "low";

arriaii_lcell_comb \pipe~175 (
	.dataa(!pipefull_1),
	.datab(!pipefull_2),
	.datac(!col_addr_5),
	.datad(!\pipe[2][5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~175_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~175 .extended_lut = "off";
defparam \pipe~175 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \pipe~175 .shared_arith = "off";

dffeas \pipe[1][5] (
	.clk(ctl_clk),
	.d(\pipe~175_combout ),
	.asdata(\pipe~163_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[1][5]~q ),
	.prn(vcc));
defparam \pipe[1][5] .is_wysiwyg = "true";
defparam \pipe[1][5] .power_up = "low";

arriaii_lcell_comb \pipe~163 (
	.dataa(!pipefull_0),
	.datab(!pipefull_1),
	.datac(!col_addr_5),
	.datad(!\pipe[1][5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~163_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~163 .extended_lut = "off";
defparam \pipe~163 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \pipe~163 .shared_arith = "off";

arriaii_lcell_comb \pipe~230 (
	.dataa(!generating),
	.datab(!buf_col_addr_6),
	.datac(!local_address_4),
	.datad(!\pipe[7][6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~230_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~230 .extended_lut = "off";
defparam \pipe~230 .lut_mask = 64'h001B001B001B001B;
defparam \pipe~230 .shared_arith = "off";

dffeas \pipe[7][6] (
	.clk(ctl_clk),
	.d(\pipe~230_combout ),
	.asdata(\pipe~223_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[7][6]~q ),
	.prn(vcc));
defparam \pipe[7][6] .is_wysiwyg = "true";
defparam \pipe[7][6] .power_up = "low";

arriaii_lcell_comb \pipe~223 (
	.dataa(!pipefull_7),
	.datab(!pipefull_6),
	.datac(!col_addr_6),
	.datad(!\pipe[7][6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~223_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~223 .extended_lut = "off";
defparam \pipe~223 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~223 .shared_arith = "off";

dffeas \pipe[6][6] (
	.clk(ctl_clk),
	.d(\pipe~223_combout ),
	.asdata(\pipe~216_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[6][6]~q ),
	.prn(vcc));
defparam \pipe[6][6] .is_wysiwyg = "true";
defparam \pipe[6][6] .power_up = "low";

arriaii_lcell_comb \pipe~216 (
	.dataa(!pipefull_6),
	.datab(!pipefull_5),
	.datac(!col_addr_6),
	.datad(!\pipe[6][6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~216_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~216 .extended_lut = "off";
defparam \pipe~216 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~216 .shared_arith = "off";

dffeas \pipe[5][6] (
	.clk(ctl_clk),
	.d(\pipe~216_combout ),
	.asdata(\pipe~208_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[5][6]~q ),
	.prn(vcc));
defparam \pipe[5][6] .is_wysiwyg = "true";
defparam \pipe[5][6] .power_up = "low";

arriaii_lcell_comb \pipe~208 (
	.dataa(!pipefull_5),
	.datab(!pipefull_4),
	.datac(!col_addr_6),
	.datad(!\pipe[5][6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~208_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~208 .extended_lut = "off";
defparam \pipe~208 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~208 .shared_arith = "off";

dffeas \pipe[4][6] (
	.clk(ctl_clk),
	.d(\pipe~208_combout ),
	.asdata(\pipe~200_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[4][6]~q ),
	.prn(vcc));
defparam \pipe[4][6] .is_wysiwyg = "true";
defparam \pipe[4][6] .power_up = "low";

arriaii_lcell_comb \pipe~200 (
	.dataa(!pipefull_4),
	.datab(!pipefull_3),
	.datac(!col_addr_6),
	.datad(!\pipe[4][6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~200_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~200 .extended_lut = "off";
defparam \pipe~200 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~200 .shared_arith = "off";

dffeas \pipe[3][6] (
	.clk(ctl_clk),
	.d(\pipe~200_combout ),
	.asdata(\pipe~188_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[3][6]~q ),
	.prn(vcc));
defparam \pipe[3][6] .is_wysiwyg = "true";
defparam \pipe[3][6] .power_up = "low";

arriaii_lcell_comb \pipe~188 (
	.dataa(!pipefull_2),
	.datab(!pipefull_3),
	.datac(!col_addr_6),
	.datad(!\pipe[3][6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~188_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~188 .extended_lut = "off";
defparam \pipe~188 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \pipe~188 .shared_arith = "off";

dffeas \pipe[2][6] (
	.clk(ctl_clk),
	.d(\pipe~188_combout ),
	.asdata(\pipe~176_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[2][6]~q ),
	.prn(vcc));
defparam \pipe[2][6] .is_wysiwyg = "true";
defparam \pipe[2][6] .power_up = "low";

arriaii_lcell_comb \pipe~176 (
	.dataa(!pipefull_1),
	.datab(!pipefull_2),
	.datac(!col_addr_6),
	.datad(!\pipe[2][6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~176_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~176 .extended_lut = "off";
defparam \pipe~176 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \pipe~176 .shared_arith = "off";

dffeas \pipe[1][6] (
	.clk(ctl_clk),
	.d(\pipe~176_combout ),
	.asdata(\pipe~164_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[1][6]~q ),
	.prn(vcc));
defparam \pipe[1][6] .is_wysiwyg = "true";
defparam \pipe[1][6] .power_up = "low";

arriaii_lcell_comb \pipe~164 (
	.dataa(!pipefull_0),
	.datab(!pipefull_1),
	.datac(!col_addr_6),
	.datad(!\pipe[1][6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~164_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~164 .extended_lut = "off";
defparam \pipe~164 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \pipe~164 .shared_arith = "off";

arriaii_lcell_comb \pipe~231 (
	.dataa(!generating),
	.datab(!buf_col_addr_7),
	.datac(!local_address_5),
	.datad(!\pipe[7][7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~231_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~231 .extended_lut = "off";
defparam \pipe~231 .lut_mask = 64'h001B001B001B001B;
defparam \pipe~231 .shared_arith = "off";

dffeas \pipe[7][7] (
	.clk(ctl_clk),
	.d(\pipe~231_combout ),
	.asdata(\pipe~224_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[7][7]~q ),
	.prn(vcc));
defparam \pipe[7][7] .is_wysiwyg = "true";
defparam \pipe[7][7] .power_up = "low";

arriaii_lcell_comb \pipe~224 (
	.dataa(!pipefull_7),
	.datab(!pipefull_6),
	.datac(!col_addr_7),
	.datad(!\pipe[7][7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~224_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~224 .extended_lut = "off";
defparam \pipe~224 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~224 .shared_arith = "off";

dffeas \pipe[6][7] (
	.clk(ctl_clk),
	.d(\pipe~224_combout ),
	.asdata(\pipe~217_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[6][7]~q ),
	.prn(vcc));
defparam \pipe[6][7] .is_wysiwyg = "true";
defparam \pipe[6][7] .power_up = "low";

arriaii_lcell_comb \pipe~217 (
	.dataa(!pipefull_6),
	.datab(!pipefull_5),
	.datac(!col_addr_7),
	.datad(!\pipe[6][7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~217_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~217 .extended_lut = "off";
defparam \pipe~217 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~217 .shared_arith = "off";

dffeas \pipe[5][7] (
	.clk(ctl_clk),
	.d(\pipe~217_combout ),
	.asdata(\pipe~209_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[5][7]~q ),
	.prn(vcc));
defparam \pipe[5][7] .is_wysiwyg = "true";
defparam \pipe[5][7] .power_up = "low";

arriaii_lcell_comb \pipe~209 (
	.dataa(!pipefull_5),
	.datab(!pipefull_4),
	.datac(!col_addr_7),
	.datad(!\pipe[5][7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~209_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~209 .extended_lut = "off";
defparam \pipe~209 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~209 .shared_arith = "off";

dffeas \pipe[4][7] (
	.clk(ctl_clk),
	.d(\pipe~209_combout ),
	.asdata(\pipe~201_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[4][7]~q ),
	.prn(vcc));
defparam \pipe[4][7] .is_wysiwyg = "true";
defparam \pipe[4][7] .power_up = "low";

arriaii_lcell_comb \pipe~201 (
	.dataa(!pipefull_4),
	.datab(!pipefull_3),
	.datac(!col_addr_7),
	.datad(!\pipe[4][7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~201_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~201 .extended_lut = "off";
defparam \pipe~201 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~201 .shared_arith = "off";

dffeas \pipe[3][7] (
	.clk(ctl_clk),
	.d(\pipe~201_combout ),
	.asdata(\pipe~189_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[3][7]~q ),
	.prn(vcc));
defparam \pipe[3][7] .is_wysiwyg = "true";
defparam \pipe[3][7] .power_up = "low";

arriaii_lcell_comb \pipe~189 (
	.dataa(!pipefull_2),
	.datab(!pipefull_3),
	.datac(!col_addr_7),
	.datad(!\pipe[3][7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~189_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~189 .extended_lut = "off";
defparam \pipe~189 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \pipe~189 .shared_arith = "off";

dffeas \pipe[2][7] (
	.clk(ctl_clk),
	.d(\pipe~189_combout ),
	.asdata(\pipe~177_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[2][7]~q ),
	.prn(vcc));
defparam \pipe[2][7] .is_wysiwyg = "true";
defparam \pipe[2][7] .power_up = "low";

arriaii_lcell_comb \pipe~177 (
	.dataa(!pipefull_1),
	.datab(!pipefull_2),
	.datac(!col_addr_7),
	.datad(!\pipe[2][7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~177_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~177 .extended_lut = "off";
defparam \pipe~177 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \pipe~177 .shared_arith = "off";

dffeas \pipe[1][7] (
	.clk(ctl_clk),
	.d(\pipe~177_combout ),
	.asdata(\pipe~165_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[1][7]~q ),
	.prn(vcc));
defparam \pipe[1][7] .is_wysiwyg = "true";
defparam \pipe[1][7] .power_up = "low";

arriaii_lcell_comb \pipe~165 (
	.dataa(!pipefull_0),
	.datab(!pipefull_1),
	.datac(!col_addr_7),
	.datad(!\pipe[1][7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~165_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~165 .extended_lut = "off";
defparam \pipe~165 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \pipe~165 .shared_arith = "off";

arriaii_lcell_comb \pipe~232 (
	.dataa(!generating),
	.datab(!buf_col_addr_8),
	.datac(!local_address_6),
	.datad(!\pipe[7][8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~232_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~232 .extended_lut = "off";
defparam \pipe~232 .lut_mask = 64'h001B001B001B001B;
defparam \pipe~232 .shared_arith = "off";

dffeas \pipe[7][8] (
	.clk(ctl_clk),
	.d(\pipe~232_combout ),
	.asdata(\pipe~225_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[7][8]~q ),
	.prn(vcc));
defparam \pipe[7][8] .is_wysiwyg = "true";
defparam \pipe[7][8] .power_up = "low";

arriaii_lcell_comb \pipe~225 (
	.dataa(!pipefull_7),
	.datab(!pipefull_6),
	.datac(!col_addr_8),
	.datad(!\pipe[7][8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~225_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~225 .extended_lut = "off";
defparam \pipe~225 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~225 .shared_arith = "off";

dffeas \pipe[6][8] (
	.clk(ctl_clk),
	.d(\pipe~225_combout ),
	.asdata(\pipe~218_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[6][8]~q ),
	.prn(vcc));
defparam \pipe[6][8] .is_wysiwyg = "true";
defparam \pipe[6][8] .power_up = "low";

arriaii_lcell_comb \pipe~218 (
	.dataa(!pipefull_6),
	.datab(!pipefull_5),
	.datac(!col_addr_8),
	.datad(!\pipe[6][8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~218_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~218 .extended_lut = "off";
defparam \pipe~218 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~218 .shared_arith = "off";

dffeas \pipe[5][8] (
	.clk(ctl_clk),
	.d(\pipe~218_combout ),
	.asdata(\pipe~210_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[5][8]~q ),
	.prn(vcc));
defparam \pipe[5][8] .is_wysiwyg = "true";
defparam \pipe[5][8] .power_up = "low";

arriaii_lcell_comb \pipe~210 (
	.dataa(!pipefull_5),
	.datab(!pipefull_4),
	.datac(!col_addr_8),
	.datad(!\pipe[5][8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~210_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~210 .extended_lut = "off";
defparam \pipe~210 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~210 .shared_arith = "off";

dffeas \pipe[4][8] (
	.clk(ctl_clk),
	.d(\pipe~210_combout ),
	.asdata(\pipe~202_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[4][8]~q ),
	.prn(vcc));
defparam \pipe[4][8] .is_wysiwyg = "true";
defparam \pipe[4][8] .power_up = "low";

arriaii_lcell_comb \pipe~202 (
	.dataa(!pipefull_4),
	.datab(!pipefull_3),
	.datac(!col_addr_8),
	.datad(!\pipe[4][8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~202_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~202 .extended_lut = "off";
defparam \pipe~202 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~202 .shared_arith = "off";

dffeas \pipe[3][8] (
	.clk(ctl_clk),
	.d(\pipe~202_combout ),
	.asdata(\pipe~190_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[3][8]~q ),
	.prn(vcc));
defparam \pipe[3][8] .is_wysiwyg = "true";
defparam \pipe[3][8] .power_up = "low";

arriaii_lcell_comb \pipe~190 (
	.dataa(!pipefull_2),
	.datab(!pipefull_3),
	.datac(!col_addr_8),
	.datad(!\pipe[3][8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~190_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~190 .extended_lut = "off";
defparam \pipe~190 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \pipe~190 .shared_arith = "off";

dffeas \pipe[2][8] (
	.clk(ctl_clk),
	.d(\pipe~190_combout ),
	.asdata(\pipe~178_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[2][8]~q ),
	.prn(vcc));
defparam \pipe[2][8] .is_wysiwyg = "true";
defparam \pipe[2][8] .power_up = "low";

arriaii_lcell_comb \pipe~178 (
	.dataa(!pipefull_1),
	.datab(!pipefull_2),
	.datac(!col_addr_8),
	.datad(!\pipe[2][8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~178_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~178 .extended_lut = "off";
defparam \pipe~178 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \pipe~178 .shared_arith = "off";

dffeas \pipe[1][8] (
	.clk(ctl_clk),
	.d(\pipe~178_combout ),
	.asdata(\pipe~166_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[1][8]~q ),
	.prn(vcc));
defparam \pipe[1][8] .is_wysiwyg = "true";
defparam \pipe[1][8] .power_up = "low";

arriaii_lcell_comb \pipe~166 (
	.dataa(!pipefull_0),
	.datab(!pipefull_1),
	.datac(!col_addr_8),
	.datad(!\pipe[1][8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~166_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~166 .extended_lut = "off";
defparam \pipe~166 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \pipe~166 .shared_arith = "off";

arriaii_lcell_comb \pipe~233 (
	.dataa(!generating),
	.datab(!buf_col_addr_9),
	.datac(!local_address_7),
	.datad(!\pipe[7][9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~233_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~233 .extended_lut = "off";
defparam \pipe~233 .lut_mask = 64'h001B001B001B001B;
defparam \pipe~233 .shared_arith = "off";

dffeas \pipe[7][9] (
	.clk(ctl_clk),
	.d(\pipe~233_combout ),
	.asdata(\pipe~226_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[7][9]~q ),
	.prn(vcc));
defparam \pipe[7][9] .is_wysiwyg = "true";
defparam \pipe[7][9] .power_up = "low";

arriaii_lcell_comb \pipe~226 (
	.dataa(!pipefull_7),
	.datab(!pipefull_6),
	.datac(!col_addr_9),
	.datad(!\pipe[7][9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~226_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~226 .extended_lut = "off";
defparam \pipe~226 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~226 .shared_arith = "off";

dffeas \pipe[6][9] (
	.clk(ctl_clk),
	.d(\pipe~226_combout ),
	.asdata(\pipe~219_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[6][9]~q ),
	.prn(vcc));
defparam \pipe[6][9] .is_wysiwyg = "true";
defparam \pipe[6][9] .power_up = "low";

arriaii_lcell_comb \pipe~219 (
	.dataa(!pipefull_6),
	.datab(!pipefull_5),
	.datac(!col_addr_9),
	.datad(!\pipe[6][9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~219_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~219 .extended_lut = "off";
defparam \pipe~219 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~219 .shared_arith = "off";

dffeas \pipe[5][9] (
	.clk(ctl_clk),
	.d(\pipe~219_combout ),
	.asdata(\pipe~211_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[5][9]~q ),
	.prn(vcc));
defparam \pipe[5][9] .is_wysiwyg = "true";
defparam \pipe[5][9] .power_up = "low";

arriaii_lcell_comb \pipe~211 (
	.dataa(!pipefull_5),
	.datab(!pipefull_4),
	.datac(!col_addr_9),
	.datad(!\pipe[5][9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~211_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~211 .extended_lut = "off";
defparam \pipe~211 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~211 .shared_arith = "off";

dffeas \pipe[4][9] (
	.clk(ctl_clk),
	.d(\pipe~211_combout ),
	.asdata(\pipe~203_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[4][9]~q ),
	.prn(vcc));
defparam \pipe[4][9] .is_wysiwyg = "true";
defparam \pipe[4][9] .power_up = "low";

arriaii_lcell_comb \pipe~203 (
	.dataa(!pipefull_4),
	.datab(!pipefull_3),
	.datac(!col_addr_9),
	.datad(!\pipe[4][9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~203_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~203 .extended_lut = "off";
defparam \pipe~203 .lut_mask = 64'h02DF02DF02DF02DF;
defparam \pipe~203 .shared_arith = "off";

dffeas \pipe[3][9] (
	.clk(ctl_clk),
	.d(\pipe~203_combout ),
	.asdata(\pipe~191_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[3][9]~q ),
	.prn(vcc));
defparam \pipe[3][9] .is_wysiwyg = "true";
defparam \pipe[3][9] .power_up = "low";

arriaii_lcell_comb \pipe~191 (
	.dataa(!pipefull_2),
	.datab(!pipefull_3),
	.datac(!col_addr_9),
	.datad(!\pipe[3][9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~191_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~191 .extended_lut = "off";
defparam \pipe~191 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \pipe~191 .shared_arith = "off";

dffeas \pipe[2][9] (
	.clk(ctl_clk),
	.d(\pipe~191_combout ),
	.asdata(\pipe~179_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[2][9]~q ),
	.prn(vcc));
defparam \pipe[2][9] .is_wysiwyg = "true";
defparam \pipe[2][9] .power_up = "low";

arriaii_lcell_comb \pipe~179 (
	.dataa(!pipefull_1),
	.datab(!pipefull_2),
	.datac(!col_addr_9),
	.datad(!\pipe[2][9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~179_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~179 .extended_lut = "off";
defparam \pipe~179 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \pipe~179 .shared_arith = "off";

dffeas \pipe[1][9] (
	.clk(ctl_clk),
	.d(\pipe~179_combout ),
	.asdata(\pipe~167_combout ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!fetch),
	.ena(\pipe[1][11]~7_combout ),
	.q(\pipe[1][9]~q ),
	.prn(vcc));
defparam \pipe[1][9] .is_wysiwyg = "true";
defparam \pipe[1][9] .power_up = "low";

arriaii_lcell_comb \pipe~167 (
	.dataa(!pipefull_0),
	.datab(!pipefull_1),
	.datac(!col_addr_9),
	.datad(!\pipe[1][9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipe~167_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipe~167 .extended_lut = "off";
defparam \pipe~167 .lut_mask = 64'h04BF04BF04BF04BF;
defparam \pipe~167 .shared_arith = "off";

arriaii_lcell_comb \pipefull~0 (
	.dataa(!pipefull_7),
	.datab(!fetch),
	.datac(!read_req),
	.datad(!write_req),
	.datae(!pipefull_6),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipefull~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipefull~0 .extended_lut = "off";
defparam \pipefull~0 .lut_mask = 64'h44444CCC44444CCC;
defparam \pipefull~0 .shared_arith = "off";

arriaii_lcell_comb \pipefull~1 (
	.dataa(!pipefull_7),
	.datab(!fetch),
	.datac(!always38),
	.datad(!pipefull_6),
	.datae(!pipefull_5),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipefull~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipefull~1 .extended_lut = "off";
defparam \pipefull~1 .lut_mask = 64'h11FDD1FD11FDD1FD;
defparam \pipefull~1 .shared_arith = "off";

arriaii_lcell_comb \pipefull~2 (
	.dataa(!fetch),
	.datab(!read_req),
	.datac(!write_req),
	.datad(!pipefull_0),
	.datae(!pipefull_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipefull~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipefull~2 .extended_lut = "off";
defparam \pipefull~2 .lut_mask = 64'h2ABF7FFF2ABF7FFF;
defparam \pipefull~2 .shared_arith = "off";

arriaii_lcell_comb \pipefull~3 (
	.dataa(!fetch),
	.datab(!always38),
	.datac(!pipefull_6),
	.datad(!pipefull_5),
	.datae(!pipefull_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipefull~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipefull~3 .extended_lut = "off";
defparam \pipefull~3 .lut_mask = 64'h05EF8DEF05EF8DEF;
defparam \pipefull~3 .shared_arith = "off";

arriaii_lcell_comb \pipefull~4 (
	.dataa(!fetch),
	.datab(!always38),
	.datac(!pipefull_0),
	.datad(!pipefull_1),
	.datae(!pipefull_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipefull~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipefull~4 .extended_lut = "off";
defparam \pipefull~4 .lut_mask = 64'h08EE5DFF08EE5DFF;
defparam \pipefull~4 .shared_arith = "off";

arriaii_lcell_comb \pipefull~5 (
	.dataa(!fetch),
	.datab(!always38),
	.datac(!pipefull_5),
	.datad(!pipefull_4),
	.datae(!pipefull_3),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipefull~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipefull~5 .extended_lut = "off";
defparam \pipefull~5 .lut_mask = 64'h05EF8DEF05EF8DEF;
defparam \pipefull~5 .shared_arith = "off";

arriaii_lcell_comb \pipefull~6 (
	.dataa(!fetch),
	.datab(!always38),
	.datac(!pipefull_1),
	.datad(!pipefull_2),
	.datae(!pipefull_3),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipefull~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipefull~6 .extended_lut = "off";
defparam \pipefull~6 .lut_mask = 64'h08EE5DFF08EE5DFF;
defparam \pipefull~6 .shared_arith = "off";

arriaii_lcell_comb \pipefull~7 (
	.dataa(!fetch),
	.datab(!always38),
	.datac(!pipefull_4),
	.datad(!pipefull_2),
	.datae(!pipefull_3),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pipefull~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pipefull~7 .extended_lut = "off";
defparam \pipefull~7 .lut_mask = 64'h058DEFEF058DEFEF;
defparam \pipefull~7 .shared_arith = "off";

endmodule

module ddr3_int_alt_ddrx_wdata_fifo (
	clk_0,
	q_b_132,
	q_b_140,
	q_b_128,
	q_b_136,
	q_b_133,
	q_b_141,
	q_b_129,
	q_b_137,
	q_b_134,
	q_b_142,
	q_b_130,
	q_b_138,
	q_b_135,
	q_b_143,
	q_b_131,
	q_b_139,
	q_b_96,
	q_b_32,
	q_b_64,
	q_b_0,
	q_b_97,
	q_b_33,
	q_b_65,
	q_b_1,
	q_b_98,
	q_b_34,
	q_b_66,
	q_b_2,
	q_b_99,
	q_b_35,
	q_b_67,
	q_b_3,
	q_b_100,
	q_b_36,
	q_b_68,
	q_b_4,
	q_b_101,
	q_b_37,
	q_b_69,
	q_b_5,
	q_b_102,
	q_b_38,
	q_b_70,
	q_b_6,
	q_b_103,
	q_b_39,
	q_b_71,
	q_b_7,
	q_b_104,
	q_b_40,
	q_b_72,
	q_b_8,
	q_b_105,
	q_b_41,
	q_b_73,
	q_b_9,
	q_b_106,
	q_b_42,
	q_b_74,
	q_b_10,
	q_b_107,
	q_b_43,
	q_b_75,
	q_b_11,
	q_b_108,
	q_b_44,
	q_b_76,
	q_b_12,
	q_b_109,
	q_b_45,
	q_b_77,
	q_b_13,
	q_b_110,
	q_b_46,
	q_b_78,
	q_b_14,
	q_b_111,
	q_b_47,
	q_b_79,
	q_b_15,
	q_b_112,
	q_b_48,
	q_b_80,
	q_b_16,
	q_b_113,
	q_b_49,
	q_b_81,
	q_b_17,
	q_b_114,
	q_b_50,
	q_b_82,
	q_b_18,
	q_b_115,
	q_b_51,
	q_b_83,
	q_b_19,
	q_b_116,
	q_b_52,
	q_b_84,
	q_b_20,
	q_b_117,
	q_b_53,
	q_b_85,
	q_b_21,
	q_b_118,
	q_b_54,
	q_b_86,
	q_b_22,
	q_b_119,
	q_b_55,
	q_b_87,
	q_b_23,
	q_b_120,
	q_b_56,
	q_b_88,
	q_b_24,
	q_b_121,
	q_b_57,
	q_b_89,
	q_b_25,
	q_b_122,
	q_b_58,
	q_b_90,
	q_b_26,
	q_b_123,
	q_b_59,
	q_b_91,
	q_b_27,
	q_b_124,
	q_b_60,
	q_b_92,
	q_b_28,
	q_b_125,
	q_b_61,
	q_b_93,
	q_b_29,
	q_b_126,
	q_b_62,
	q_b_94,
	q_b_30,
	q_b_127,
	q_b_63,
	q_b_95,
	q_b_31,
	dffe_af,
	ready_out,
	avalon_write_req,
	ecc_wdata_fifo_read,
	reset_reg_3,
	local_write_req,
	local_be_4,
	local_be_12,
	local_be_0,
	local_be_8,
	local_be_5,
	local_be_13,
	local_be_1,
	local_be_9,
	local_be_6,
	local_be_14,
	local_be_2,
	local_be_10,
	local_be_7,
	local_be_15,
	local_be_3,
	local_be_11,
	local_wdata_96,
	local_wdata_32,
	local_wdata_64,
	local_wdata_0,
	local_wdata_97,
	local_wdata_33,
	local_wdata_65,
	local_wdata_1,
	local_wdata_98,
	local_wdata_34,
	local_wdata_66,
	local_wdata_2,
	local_wdata_99,
	local_wdata_35,
	local_wdata_67,
	local_wdata_3,
	local_wdata_100,
	local_wdata_36,
	local_wdata_68,
	local_wdata_4,
	local_wdata_101,
	local_wdata_37,
	local_wdata_69,
	local_wdata_5,
	local_wdata_102,
	local_wdata_38,
	local_wdata_70,
	local_wdata_6,
	local_wdata_103,
	local_wdata_39,
	local_wdata_71,
	local_wdata_7,
	local_wdata_104,
	local_wdata_40,
	local_wdata_72,
	local_wdata_8,
	local_wdata_105,
	local_wdata_41,
	local_wdata_73,
	local_wdata_9,
	local_wdata_106,
	local_wdata_42,
	local_wdata_74,
	local_wdata_10,
	local_wdata_107,
	local_wdata_43,
	local_wdata_75,
	local_wdata_11,
	local_wdata_108,
	local_wdata_44,
	local_wdata_76,
	local_wdata_12,
	local_wdata_109,
	local_wdata_45,
	local_wdata_77,
	local_wdata_13,
	local_wdata_110,
	local_wdata_46,
	local_wdata_78,
	local_wdata_14,
	local_wdata_111,
	local_wdata_47,
	local_wdata_79,
	local_wdata_15,
	local_wdata_112,
	local_wdata_48,
	local_wdata_80,
	local_wdata_16,
	local_wdata_113,
	local_wdata_49,
	local_wdata_81,
	local_wdata_17,
	local_wdata_114,
	local_wdata_50,
	local_wdata_82,
	local_wdata_18,
	local_wdata_115,
	local_wdata_51,
	local_wdata_83,
	local_wdata_19,
	local_wdata_116,
	local_wdata_52,
	local_wdata_84,
	local_wdata_20,
	local_wdata_117,
	local_wdata_53,
	local_wdata_85,
	local_wdata_21,
	local_wdata_118,
	local_wdata_54,
	local_wdata_86,
	local_wdata_22,
	local_wdata_119,
	local_wdata_55,
	local_wdata_87,
	local_wdata_23,
	local_wdata_120,
	local_wdata_56,
	local_wdata_88,
	local_wdata_24,
	local_wdata_121,
	local_wdata_57,
	local_wdata_89,
	local_wdata_25,
	local_wdata_122,
	local_wdata_58,
	local_wdata_90,
	local_wdata_26,
	local_wdata_123,
	local_wdata_59,
	local_wdata_91,
	local_wdata_27,
	local_wdata_124,
	local_wdata_60,
	local_wdata_92,
	local_wdata_28,
	local_wdata_125,
	local_wdata_61,
	local_wdata_93,
	local_wdata_29,
	local_wdata_126,
	local_wdata_62,
	local_wdata_94,
	local_wdata_30,
	local_wdata_127,
	local_wdata_63,
	local_wdata_95,
	local_wdata_31)/* synthesis synthesis_greybox=0 */;
input 	clk_0;
output 	q_b_132;
output 	q_b_140;
output 	q_b_128;
output 	q_b_136;
output 	q_b_133;
output 	q_b_141;
output 	q_b_129;
output 	q_b_137;
output 	q_b_134;
output 	q_b_142;
output 	q_b_130;
output 	q_b_138;
output 	q_b_135;
output 	q_b_143;
output 	q_b_131;
output 	q_b_139;
output 	q_b_96;
output 	q_b_32;
output 	q_b_64;
output 	q_b_0;
output 	q_b_97;
output 	q_b_33;
output 	q_b_65;
output 	q_b_1;
output 	q_b_98;
output 	q_b_34;
output 	q_b_66;
output 	q_b_2;
output 	q_b_99;
output 	q_b_35;
output 	q_b_67;
output 	q_b_3;
output 	q_b_100;
output 	q_b_36;
output 	q_b_68;
output 	q_b_4;
output 	q_b_101;
output 	q_b_37;
output 	q_b_69;
output 	q_b_5;
output 	q_b_102;
output 	q_b_38;
output 	q_b_70;
output 	q_b_6;
output 	q_b_103;
output 	q_b_39;
output 	q_b_71;
output 	q_b_7;
output 	q_b_104;
output 	q_b_40;
output 	q_b_72;
output 	q_b_8;
output 	q_b_105;
output 	q_b_41;
output 	q_b_73;
output 	q_b_9;
output 	q_b_106;
output 	q_b_42;
output 	q_b_74;
output 	q_b_10;
output 	q_b_107;
output 	q_b_43;
output 	q_b_75;
output 	q_b_11;
output 	q_b_108;
output 	q_b_44;
output 	q_b_76;
output 	q_b_12;
output 	q_b_109;
output 	q_b_45;
output 	q_b_77;
output 	q_b_13;
output 	q_b_110;
output 	q_b_46;
output 	q_b_78;
output 	q_b_14;
output 	q_b_111;
output 	q_b_47;
output 	q_b_79;
output 	q_b_15;
output 	q_b_112;
output 	q_b_48;
output 	q_b_80;
output 	q_b_16;
output 	q_b_113;
output 	q_b_49;
output 	q_b_81;
output 	q_b_17;
output 	q_b_114;
output 	q_b_50;
output 	q_b_82;
output 	q_b_18;
output 	q_b_115;
output 	q_b_51;
output 	q_b_83;
output 	q_b_19;
output 	q_b_116;
output 	q_b_52;
output 	q_b_84;
output 	q_b_20;
output 	q_b_117;
output 	q_b_53;
output 	q_b_85;
output 	q_b_21;
output 	q_b_118;
output 	q_b_54;
output 	q_b_86;
output 	q_b_22;
output 	q_b_119;
output 	q_b_55;
output 	q_b_87;
output 	q_b_23;
output 	q_b_120;
output 	q_b_56;
output 	q_b_88;
output 	q_b_24;
output 	q_b_121;
output 	q_b_57;
output 	q_b_89;
output 	q_b_25;
output 	q_b_122;
output 	q_b_58;
output 	q_b_90;
output 	q_b_26;
output 	q_b_123;
output 	q_b_59;
output 	q_b_91;
output 	q_b_27;
output 	q_b_124;
output 	q_b_60;
output 	q_b_92;
output 	q_b_28;
output 	q_b_125;
output 	q_b_61;
output 	q_b_93;
output 	q_b_29;
output 	q_b_126;
output 	q_b_62;
output 	q_b_94;
output 	q_b_30;
output 	q_b_127;
output 	q_b_63;
output 	q_b_95;
output 	q_b_31;
output 	dffe_af;
input 	ready_out;
input 	avalon_write_req;
input 	ecc_wdata_fifo_read;
input 	reset_reg_3;
input 	local_write_req;
input 	local_be_4;
input 	local_be_12;
input 	local_be_0;
input 	local_be_8;
input 	local_be_5;
input 	local_be_13;
input 	local_be_1;
input 	local_be_9;
input 	local_be_6;
input 	local_be_14;
input 	local_be_2;
input 	local_be_10;
input 	local_be_7;
input 	local_be_15;
input 	local_be_3;
input 	local_be_11;
input 	local_wdata_96;
input 	local_wdata_32;
input 	local_wdata_64;
input 	local_wdata_0;
input 	local_wdata_97;
input 	local_wdata_33;
input 	local_wdata_65;
input 	local_wdata_1;
input 	local_wdata_98;
input 	local_wdata_34;
input 	local_wdata_66;
input 	local_wdata_2;
input 	local_wdata_99;
input 	local_wdata_35;
input 	local_wdata_67;
input 	local_wdata_3;
input 	local_wdata_100;
input 	local_wdata_36;
input 	local_wdata_68;
input 	local_wdata_4;
input 	local_wdata_101;
input 	local_wdata_37;
input 	local_wdata_69;
input 	local_wdata_5;
input 	local_wdata_102;
input 	local_wdata_38;
input 	local_wdata_70;
input 	local_wdata_6;
input 	local_wdata_103;
input 	local_wdata_39;
input 	local_wdata_71;
input 	local_wdata_7;
input 	local_wdata_104;
input 	local_wdata_40;
input 	local_wdata_72;
input 	local_wdata_8;
input 	local_wdata_105;
input 	local_wdata_41;
input 	local_wdata_73;
input 	local_wdata_9;
input 	local_wdata_106;
input 	local_wdata_42;
input 	local_wdata_74;
input 	local_wdata_10;
input 	local_wdata_107;
input 	local_wdata_43;
input 	local_wdata_75;
input 	local_wdata_11;
input 	local_wdata_108;
input 	local_wdata_44;
input 	local_wdata_76;
input 	local_wdata_12;
input 	local_wdata_109;
input 	local_wdata_45;
input 	local_wdata_77;
input 	local_wdata_13;
input 	local_wdata_110;
input 	local_wdata_46;
input 	local_wdata_78;
input 	local_wdata_14;
input 	local_wdata_111;
input 	local_wdata_47;
input 	local_wdata_79;
input 	local_wdata_15;
input 	local_wdata_112;
input 	local_wdata_48;
input 	local_wdata_80;
input 	local_wdata_16;
input 	local_wdata_113;
input 	local_wdata_49;
input 	local_wdata_81;
input 	local_wdata_17;
input 	local_wdata_114;
input 	local_wdata_50;
input 	local_wdata_82;
input 	local_wdata_18;
input 	local_wdata_115;
input 	local_wdata_51;
input 	local_wdata_83;
input 	local_wdata_19;
input 	local_wdata_116;
input 	local_wdata_52;
input 	local_wdata_84;
input 	local_wdata_20;
input 	local_wdata_117;
input 	local_wdata_53;
input 	local_wdata_85;
input 	local_wdata_21;
input 	local_wdata_118;
input 	local_wdata_54;
input 	local_wdata_86;
input 	local_wdata_22;
input 	local_wdata_119;
input 	local_wdata_55;
input 	local_wdata_87;
input 	local_wdata_23;
input 	local_wdata_120;
input 	local_wdata_56;
input 	local_wdata_88;
input 	local_wdata_24;
input 	local_wdata_121;
input 	local_wdata_57;
input 	local_wdata_89;
input 	local_wdata_25;
input 	local_wdata_122;
input 	local_wdata_58;
input 	local_wdata_90;
input 	local_wdata_26;
input 	local_wdata_123;
input 	local_wdata_59;
input 	local_wdata_91;
input 	local_wdata_27;
input 	local_wdata_124;
input 	local_wdata_60;
input 	local_wdata_92;
input 	local_wdata_28;
input 	local_wdata_125;
input 	local_wdata_61;
input 	local_wdata_93;
input 	local_wdata_29;
input 	local_wdata_126;
input 	local_wdata_62;
input 	local_wdata_94;
input 	local_wdata_30;
input 	local_wdata_127;
input 	local_wdata_63;
input 	local_wdata_95;
input 	local_wdata_31;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_scfifo_1 wdata_fifo(
	.clock(clk_0),
	.q({q_b_143,q_b_142,q_b_141,q_b_140,q_b_139,q_b_138,q_b_137,q_b_136,q_b_135,q_b_134,q_b_133,q_b_132,q_b_131,q_b_130,q_b_129,q_b_128,q_b_127,q_b_126,q_b_125,q_b_124,q_b_123,q_b_122,q_b_121,q_b_120,q_b_119,q_b_118,q_b_117,q_b_116,q_b_115,q_b_114,q_b_113,q_b_112,q_b_111,q_b_110,q_b_109,q_b_108,
q_b_107,q_b_106,q_b_105,q_b_104,q_b_103,q_b_102,q_b_101,q_b_100,q_b_99,q_b_98,q_b_97,q_b_96,q_b_95,q_b_94,q_b_93,q_b_92,q_b_91,q_b_90,q_b_89,q_b_88,q_b_87,q_b_86,q_b_85,q_b_84,q_b_83,q_b_82,q_b_81,q_b_80,q_b_79,q_b_78,q_b_77,q_b_76,q_b_75,q_b_74,q_b_73,q_b_72,q_b_71,q_b_70,q_b_69,q_b_68,q_b_67,
q_b_66,q_b_65,q_b_64,q_b_63,q_b_62,q_b_61,q_b_60,q_b_59,q_b_58,q_b_57,q_b_56,q_b_55,q_b_54,q_b_53,q_b_52,q_b_51,q_b_50,q_b_49,q_b_48,q_b_47,q_b_46,q_b_45,q_b_44,q_b_43,q_b_42,q_b_41,q_b_40,q_b_39,q_b_38,q_b_37,q_b_36,q_b_35,q_b_34,q_b_33,q_b_32,q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,
q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.dffe_af(dffe_af),
	.ready_out(ready_out),
	.wrreq(avalon_write_req),
	.rdreq(ecc_wdata_fifo_read),
	.reset_reg_3(reset_reg_3),
	.local_write_req(local_write_req),
	.data({local_be_15,local_be_14,local_be_13,local_be_12,local_be_11,local_be_10,local_be_9,local_be_8,local_be_7,local_be_6,local_be_5,local_be_4,local_be_3,local_be_2,local_be_1,local_be_0,local_wdata_127,local_wdata_126,local_wdata_125,local_wdata_124,local_wdata_123,local_wdata_122,
local_wdata_121,local_wdata_120,local_wdata_119,local_wdata_118,local_wdata_117,local_wdata_116,local_wdata_115,local_wdata_114,local_wdata_113,local_wdata_112,local_wdata_111,local_wdata_110,local_wdata_109,local_wdata_108,local_wdata_107,local_wdata_106,local_wdata_105,
local_wdata_104,local_wdata_103,local_wdata_102,local_wdata_101,local_wdata_100,local_wdata_99,local_wdata_98,local_wdata_97,local_wdata_96,local_wdata_95,local_wdata_94,local_wdata_93,local_wdata_92,local_wdata_91,local_wdata_90,local_wdata_89,local_wdata_88,
local_wdata_87,local_wdata_86,local_wdata_85,local_wdata_84,local_wdata_83,local_wdata_82,local_wdata_81,local_wdata_80,local_wdata_79,local_wdata_78,local_wdata_77,local_wdata_76,local_wdata_75,local_wdata_74,local_wdata_73,local_wdata_72,local_wdata_71,local_wdata_70,
local_wdata_69,local_wdata_68,local_wdata_67,local_wdata_66,local_wdata_65,local_wdata_64,local_wdata_63,local_wdata_62,local_wdata_61,local_wdata_60,local_wdata_59,local_wdata_58,local_wdata_57,local_wdata_56,local_wdata_55,local_wdata_54,local_wdata_53,local_wdata_52,
local_wdata_51,local_wdata_50,local_wdata_49,local_wdata_48,local_wdata_47,local_wdata_46,local_wdata_45,local_wdata_44,local_wdata_43,local_wdata_42,local_wdata_41,local_wdata_40,local_wdata_39,local_wdata_38,local_wdata_37,local_wdata_36,local_wdata_35,local_wdata_34,
local_wdata_33,local_wdata_32,local_wdata_31,local_wdata_30,local_wdata_29,local_wdata_28,local_wdata_27,local_wdata_26,local_wdata_25,local_wdata_24,local_wdata_23,local_wdata_22,local_wdata_21,local_wdata_20,local_wdata_19,local_wdata_18,local_wdata_17,local_wdata_16,
local_wdata_15,local_wdata_14,local_wdata_13,local_wdata_12,local_wdata_11,local_wdata_10,local_wdata_9,local_wdata_8,local_wdata_7,local_wdata_6,local_wdata_5,local_wdata_4,local_wdata_3,local_wdata_2,local_wdata_1,local_wdata_0}));

endmodule

module ddr3_int_scfifo_1 (
	clock,
	q,
	dffe_af,
	ready_out,
	wrreq,
	rdreq,
	reset_reg_3,
	local_write_req,
	data)/* synthesis synthesis_greybox=0 */;
input 	clock;
output 	[143:0] q;
output 	dffe_af;
input 	ready_out;
input 	wrreq;
input 	rdreq;
input 	reset_reg_3;
input 	local_write_req;
input 	[143:0] data;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_scfifo_2a61 auto_generated(
	.clock(clock),
	.q({q[143],q[142],q[141],q[140],q[139],q[138],q[137],q[136],q[135],q[134],q[133],q[132],q[131],q[130],q[129],q[128],q[127],q[126],q[125],q[124],q[123],q[122],q[121],q[120],q[119],q[118],q[117],q[116],q[115],q[114],q[113],q[112],q[111],q[110],q[109],q[108],q[107],q[106],q[105],q[104],q[103],q[102],q[101],q[100],q[99],q[98],q[97],q[96],q[95],q[94],q[93],q[92],q[91],q[90],q[89],q[88],q[87],q[86],q[85],q[84],q[83],q[82],q[81],q[80],q[79],q[78],q[77],q[76],q[75],q[74],q[73],q[72],q[71],q[70],q[69],q[68],q[67],q[66],q[65],q[64],q[63],q[62],q[61],q[60],q[59],q[58],q[57],q[56],q[55],q[54],q[53],q[52],q[51],q[50],q[49],q[48],q[47],q[46],q[45],q[44],q[43],q[42],q[41],q[40],q[39],q[38],q[37],q[36],q[35],q[34],q[33],q[32],q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.dffe_af1(dffe_af),
	.ready_out(ready_out),
	.wrreq(wrreq),
	.rdreq(rdreq),
	.reset_reg_3(reset_reg_3),
	.local_write_req(local_write_req),
	.data({data[143],data[142],data[141],data[140],data[139],data[138],data[137],data[136],data[135],data[134],data[133],data[132],data[131],data[130],data[129],data[128],data[127],data[126],data[125],data[124],data[123],data[122],data[121],data[120],data[119],data[118],data[117],data[116],data[115],data[114],data[113],data[112],data[111],data[110],data[109],data[108],data[107],data[106],data[105],data[104],data[103],data[102],data[101],data[100],data[99],data[98],data[97],data[96],data[95],data[94],data[93],data[92],data[91],data[90],data[89],data[88],data[87],data[86],data[85],data[84],data[83],data[82],data[81],data[80],
data[79],data[78],data[77],data[76],data[75],data[74],data[73],data[72],data[71],data[70],data[69],data[68],data[67],data[66],data[65],data[64],data[63],data[62],data[61],data[60],data[59],data[58],data[57],data[56],data[55],data[54],data[53],data[52],data[51],data[50],data[49],data[48],data[47],data[46],data[45],data[44],data[43],data[42],data[41],data[40],data[39],data[38],data[37],data[36],data[35],data[34],data[33],data[32],data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],
data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}));

endmodule

module ddr3_int_scfifo_2a61 (
	clock,
	q,
	dffe_af1,
	ready_out,
	wrreq,
	rdreq,
	reset_reg_3,
	local_write_req,
	data)/* synthesis synthesis_greybox=0 */;
input 	clock;
output 	[143:0] q;
output 	dffe_af1;
input 	ready_out;
input 	wrreq;
input 	rdreq;
input 	reset_reg_3;
input 	local_write_req;
input 	[143:0] data;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \dpfifo|usedw_counter|counter_reg_bit[5]~q ;
wire \dpfifo|usedw_counter|counter_reg_bit[7]~q ;
wire \dpfifo|usedw_counter|counter_reg_bit[6]~q ;
wire \dpfifo|usedw_counter|counter_reg_bit[0]~q ;
wire \dpfifo|usedw_counter|counter_reg_bit[1]~q ;
wire \dpfifo|usedw_counter|counter_reg_bit[2]~q ;
wire \dpfifo|usedw_counter|counter_reg_bit[4]~q ;
wire \dpfifo|usedw_counter|counter_reg_bit[3]~q ;
wire \dffe_af~0_combout ;
wire \dffe_af~1_combout ;
wire \dffe_af~2_combout ;
wire \dffe_af~3_combout ;


ddr3_int_a_dpfifo_0131 dpfifo(
	.clock(clock),
	.q({q[143],q[142],q[141],q[140],q[139],q[138],q[137],q[136],q[135],q[134],q[133],q[132],q[131],q[130],q[129],q[128],q[127],q[126],q[125],q[124],q[123],q[122],q[121],q[120],q[119],q[118],q[117],q[116],q[115],q[114],q[113],q[112],q[111],q[110],q[109],q[108],q[107],q[106],q[105],q[104],q[103],q[102],q[101],q[100],q[99],q[98],q[97],q[96],q[95],q[94],q[93],q[92],q[91],q[90],q[89],q[88],q[87],q[86],q[85],q[84],q[83],q[82],q[81],q[80],q[79],q[78],q[77],q[76],q[75],q[74],q[73],q[72],q[71],q[70],q[69],q[68],q[67],q[66],q[65],q[64],q[63],q[62],q[61],q[60],q[59],q[58],q[57],q[56],q[55],q[54],q[53],q[52],q[51],q[50],q[49],q[48],q[47],q[46],q[45],q[44],q[43],q[42],q[41],q[40],q[39],q[38],q[37],q[36],q[35],q[34],q[33],q[32],q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.ready_out(ready_out),
	.wreq(wrreq),
	.counter_reg_bit_5(\dpfifo|usedw_counter|counter_reg_bit[5]~q ),
	.counter_reg_bit_7(\dpfifo|usedw_counter|counter_reg_bit[7]~q ),
	.counter_reg_bit_6(\dpfifo|usedw_counter|counter_reg_bit[6]~q ),
	.rreq(rdreq),
	.counter_reg_bit_0(\dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.counter_reg_bit_4(\dpfifo|usedw_counter|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\dpfifo|usedw_counter|counter_reg_bit[3]~q ),
	.reset_reg_3(reset_reg_3),
	.local_write_req(local_write_req),
	.data({data[143],data[142],data[141],data[140],data[139],data[138],data[137],data[136],data[135],data[134],data[133],data[132],data[131],data[130],data[129],data[128],data[127],data[126],data[125],data[124],data[123],data[122],data[121],data[120],data[119],data[118],data[117],data[116],data[115],data[114],data[113],data[112],data[111],data[110],data[109],data[108],data[107],data[106],data[105],data[104],data[103],data[102],data[101],data[100],data[99],data[98],data[97],data[96],data[95],data[94],data[93],data[92],data[91],data[90],data[89],data[88],data[87],data[86],data[85],data[84],data[83],data[82],data[81],data[80],
data[79],data[78],data[77],data[76],data[75],data[74],data[73],data[72],data[71],data[70],data[69],data[68],data[67],data[66],data[65],data[64],data[63],data[62],data[61],data[60],data[59],data[58],data[57],data[56],data[55],data[54],data[53],data[52],data[51],data[50],data[49],data[48],data[47],data[46],data[45],data[44],data[43],data[42],data[41],data[40],data[39],data[38],data[37],data[36],data[35],data[34],data[33],data[32],data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],
data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}));

dffeas dffe_af(
	.clk(clock),
	.d(\dffe_af~3_combout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dffe_af1),
	.prn(vcc));
defparam dffe_af.is_wysiwyg = "true";
defparam dffe_af.power_up = "low";

arriaii_lcell_comb \dffe_af~0 (
	.dataa(!\dpfifo|usedw_counter|counter_reg_bit[5]~q ),
	.datab(!\dpfifo|usedw_counter|counter_reg_bit[7]~q ),
	.datac(!\dpfifo|usedw_counter|counter_reg_bit[6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffe_af~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffe_af~0 .extended_lut = "off";
defparam \dffe_af~0 .lut_mask = 64'h0101010101010101;
defparam \dffe_af~0 .shared_arith = "off";

arriaii_lcell_comb \dffe_af~1 (
	.dataa(!\dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.datab(!\dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.datac(!\dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.datad(!\dpfifo|usedw_counter|counter_reg_bit[4]~q ),
	.datae(!\dpfifo|usedw_counter|counter_reg_bit[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffe_af~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffe_af~1 .extended_lut = "off";
defparam \dffe_af~1 .lut_mask = 64'h0080000000800000;
defparam \dffe_af~1 .shared_arith = "off";

arriaii_lcell_comb \dffe_af~2 (
	.dataa(!\dpfifo|usedw_counter|counter_reg_bit[0]~q ),
	.datab(!\dpfifo|usedw_counter|counter_reg_bit[1]~q ),
	.datac(!\dpfifo|usedw_counter|counter_reg_bit[2]~q ),
	.datad(!\dpfifo|usedw_counter|counter_reg_bit[4]~q ),
	.datae(!\dpfifo|usedw_counter|counter_reg_bit[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffe_af~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffe_af~2 .extended_lut = "off";
defparam \dffe_af~2 .lut_mask = 64'h0000010000000100;
defparam \dffe_af~2 .shared_arith = "off";

arriaii_lcell_comb \dffe_af~3 (
	.dataa(!dffe_af1),
	.datab(!wrreq),
	.datac(!\dffe_af~0_combout ),
	.datad(!rdreq),
	.datae(!\dffe_af~1_combout ),
	.dataf(!\dffe_af~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dffe_af~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffe_af~3 .extended_lut = "off";
defparam \dffe_af~3 .lut_mask = 64'h5555555057555750;
defparam \dffe_af~3 .shared_arith = "off";

endmodule

module ddr3_int_a_dpfifo_0131 (
	clock,
	q,
	ready_out,
	wreq,
	counter_reg_bit_5,
	counter_reg_bit_7,
	counter_reg_bit_6,
	rreq,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_4,
	counter_reg_bit_3,
	reset_reg_3,
	local_write_req,
	data)/* synthesis synthesis_greybox=0 */;
input 	clock;
output 	[143:0] q;
input 	ready_out;
input 	wreq;
output 	counter_reg_bit_5;
output 	counter_reg_bit_7;
output 	counter_reg_bit_6;
input 	rreq;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
input 	reset_reg_3;
input 	local_write_req;
input 	[143:0] data;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \_~0_combout ;
wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \wr_ptr|counter_reg_bit[5]~q ;
wire \wr_ptr|counter_reg_bit[6]~q ;
wire \wr_ptr|counter_reg_bit[7]~q ;
wire \rd_ptr_lsb~q ;
wire \low_addressa[0]~q ;
wire \ram_read_address[0]~0_combout ;
wire \rd_ptr_msb|counter_reg_bit[0]~q ;
wire \low_addressa[1]~q ;
wire \ram_read_address[1]~1_combout ;
wire \rd_ptr_msb|counter_reg_bit[1]~q ;
wire \low_addressa[2]~q ;
wire \ram_read_address[2]~2_combout ;
wire \rd_ptr_msb|counter_reg_bit[2]~q ;
wire \low_addressa[3]~q ;
wire \ram_read_address[3]~3_combout ;
wire \rd_ptr_msb|counter_reg_bit[3]~q ;
wire \low_addressa[4]~q ;
wire \ram_read_address[4]~4_combout ;
wire \rd_ptr_msb|counter_reg_bit[4]~q ;
wire \low_addressa[5]~q ;
wire \ram_read_address[5]~5_combout ;
wire \rd_ptr_msb|counter_reg_bit[5]~q ;
wire \low_addressa[6]~q ;
wire \ram_read_address[6]~6_combout ;
wire \rd_ptr_msb|counter_reg_bit[6]~q ;
wire \low_addressa[7]~q ;
wire \ram_read_address[7]~7_combout ;
wire \_~1_combout ;
wire \rd_ptr_lsb~0_combout ;


ddr3_int_cntr_hkb rd_ptr_msb(
	.clock(clock),
	.reset_reg_3(reset_reg_3),
	.counter_reg_bit_0(\rd_ptr_msb|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_msb|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_msb|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_msb|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\rd_ptr_msb|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\rd_ptr_msb|counter_reg_bit[5]~q ),
	.counter_reg_bit_6(\rd_ptr_msb|counter_reg_bit[6]~q ),
	._(\_~1_combout ));

ddr3_int_cntr_uk7 usedw_counter(
	.clock(clock),
	.avalon_write_req(wreq),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_7(counter_reg_bit_7),
	.counter_reg_bit_6(counter_reg_bit_6),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.reset_reg_3(reset_reg_3),
	._(\_~0_combout ));

ddr3_int_cntr_ikb wr_ptr(
	.clock(clock),
	.avalon_write_req(wreq),
	.reset_reg_3(reset_reg_3),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\wr_ptr|counter_reg_bit[5]~q ),
	.counter_reg_bit_6(\wr_ptr|counter_reg_bit[6]~q ),
	.counter_reg_bit_7(\wr_ptr|counter_reg_bit[7]~q ));

ddr3_int_altsyncram_u1e1 FIFOram(
	.clock0(clock),
	.clock1(clock),
	.q_b({q[143],q[142],q[141],q[140],q[139],q[138],q[137],q[136],q[135],q[134],q[133],q[132],q[131],q[130],q[129],q[128],q[127],q[126],q[125],q[124],q[123],q[122],q[121],q[120],q[119],q[118],q[117],q[116],q[115],q[114],q[113],q[112],q[111],q[110],q[109],q[108],q[107],q[106],q[105],q[104],q[103],q[102],q[101],q[100],q[99],q[98],q[97],q[96],q[95],q[94],q[93],q[92],q[91],q[90],q[89],q[88],q[87],q[86],q[85],q[84],q[83],q[82],q[81],q[80],q[79],q[78],q[77],q[76],q[75],q[74],q[73],q[72],q[71],q[70],q[69],q[68],q[67],q[66],q[65],q[64],q[63],q[62],q[61],q[60],q[59],q[58],q[57],q[56],q[55],q[54],q[53],q[52],q[51],q[50],q[49],q[48],q[47],q[46],q[45],q[44],q[43],q[42],q[41],q[40],q[39],q[38],q[37],q[36],q[35],q[34],q[33],q[32],q[31],q[30],q[29],q[28],q[27],q[26],q[25],q[24],q[23],q[22],q[21],q[20],q[19],q[18],q[17],q[16],q[15],q[14],q[13],q[12],q[11],q[10],q[9],q[8],q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.wren_a(wreq),
	.clocken1(rreq),
	.address_a({\wr_ptr|counter_reg_bit[7]~q ,\wr_ptr|counter_reg_bit[6]~q ,\wr_ptr|counter_reg_bit[5]~q ,\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.address_b({\ram_read_address[7]~7_combout ,\ram_read_address[6]~6_combout ,\ram_read_address[5]~5_combout ,\ram_read_address[4]~4_combout ,\ram_read_address[3]~3_combout ,\ram_read_address[2]~2_combout ,\ram_read_address[1]~1_combout ,\ram_read_address[0]~0_combout }),
	.data_a({data[143],data[142],data[141],data[140],data[139],data[138],data[137],data[136],data[135],data[134],data[133],data[132],data[131],data[130],data[129],data[128],data[127],data[126],data[125],data[124],data[123],data[122],data[121],data[120],data[119],data[118],data[117],data[116],data[115],data[114],data[113],data[112],data[111],data[110],data[109],data[108],data[107],data[106],data[105],data[104],data[103],data[102],data[101],data[100],data[99],data[98],data[97],data[96],data[95],data[94],data[93],data[92],data[91],data[90],data[89],data[88],data[87],data[86],data[85],data[84],data[83],data[82],data[81],data[80],
data[79],data[78],data[77],data[76],data[75],data[74],data[73],data[72],data[71],data[70],data[69],data[68],data[67],data[66],data[65],data[64],data[63],data[62],data[61],data[60],data[59],data[58],data[57],data[56],data[55],data[54],data[53],data[52],data[51],data[50],data[49],data[48],data[47],data[46],data[45],data[44],data[43],data[42],data[41],data[40],data[39],data[38],data[37],data[36],data[35],data[34],data[33],data[32],data[31],data[30],data[29],data[28],data[27],data[26],data[25],data[24],data[23],data[22],data[21],data[20],data[19],data[18],data[17],data[16],
data[15],data[14],data[13],data[12],data[11],data[10],data[9],data[8],data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}));

arriaii_lcell_comb \_~0 (
	.dataa(!ready_out),
	.datab(!local_write_req),
	.datac(!rreq),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~0 .extended_lut = "off";
defparam \_~0 .lut_mask = 64'h1E1E1E1E1E1E1E1E;
defparam \_~0 .shared_arith = "off";

dffeas rd_ptr_lsb(
	.clk(clock),
	.d(\rd_ptr_lsb~0_combout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rreq),
	.q(\rd_ptr_lsb~q ),
	.prn(vcc));
defparam rd_ptr_lsb.is_wysiwyg = "true";
defparam rd_ptr_lsb.power_up = "low";

dffeas \low_addressa[0] (
	.clk(clock),
	.d(\ram_read_address[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[0]~q ),
	.prn(vcc));
defparam \low_addressa[0] .is_wysiwyg = "true";
defparam \low_addressa[0] .power_up = "low";

arriaii_lcell_comb \ram_read_address[0]~0 (
	.dataa(!rreq),
	.datab(!\rd_ptr_lsb~q ),
	.datac(!\low_addressa[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_read_address[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_read_address[0]~0 .extended_lut = "off";
defparam \ram_read_address[0]~0 .lut_mask = 64'h4E4E4E4E4E4E4E4E;
defparam \ram_read_address[0]~0 .shared_arith = "off";

dffeas \low_addressa[1] (
	.clk(clock),
	.d(\ram_read_address[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[1]~q ),
	.prn(vcc));
defparam \low_addressa[1] .is_wysiwyg = "true";
defparam \low_addressa[1] .power_up = "low";

arriaii_lcell_comb \ram_read_address[1]~1 (
	.dataa(!rreq),
	.datab(!\rd_ptr_msb|counter_reg_bit[0]~q ),
	.datac(!\low_addressa[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_read_address[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_read_address[1]~1 .extended_lut = "off";
defparam \ram_read_address[1]~1 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \ram_read_address[1]~1 .shared_arith = "off";

dffeas \low_addressa[2] (
	.clk(clock),
	.d(\ram_read_address[2]~2_combout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[2]~q ),
	.prn(vcc));
defparam \low_addressa[2] .is_wysiwyg = "true";
defparam \low_addressa[2] .power_up = "low";

arriaii_lcell_comb \ram_read_address[2]~2 (
	.dataa(!rreq),
	.datab(!\rd_ptr_msb|counter_reg_bit[1]~q ),
	.datac(!\low_addressa[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_read_address[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_read_address[2]~2 .extended_lut = "off";
defparam \ram_read_address[2]~2 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \ram_read_address[2]~2 .shared_arith = "off";

dffeas \low_addressa[3] (
	.clk(clock),
	.d(\ram_read_address[3]~3_combout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[3]~q ),
	.prn(vcc));
defparam \low_addressa[3] .is_wysiwyg = "true";
defparam \low_addressa[3] .power_up = "low";

arriaii_lcell_comb \ram_read_address[3]~3 (
	.dataa(!rreq),
	.datab(!\rd_ptr_msb|counter_reg_bit[2]~q ),
	.datac(!\low_addressa[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_read_address[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_read_address[3]~3 .extended_lut = "off";
defparam \ram_read_address[3]~3 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \ram_read_address[3]~3 .shared_arith = "off";

dffeas \low_addressa[4] (
	.clk(clock),
	.d(\ram_read_address[4]~4_combout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[4]~q ),
	.prn(vcc));
defparam \low_addressa[4] .is_wysiwyg = "true";
defparam \low_addressa[4] .power_up = "low";

arriaii_lcell_comb \ram_read_address[4]~4 (
	.dataa(!rreq),
	.datab(!\rd_ptr_msb|counter_reg_bit[3]~q ),
	.datac(!\low_addressa[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_read_address[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_read_address[4]~4 .extended_lut = "off";
defparam \ram_read_address[4]~4 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \ram_read_address[4]~4 .shared_arith = "off";

dffeas \low_addressa[5] (
	.clk(clock),
	.d(\ram_read_address[5]~5_combout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[5]~q ),
	.prn(vcc));
defparam \low_addressa[5] .is_wysiwyg = "true";
defparam \low_addressa[5] .power_up = "low";

arriaii_lcell_comb \ram_read_address[5]~5 (
	.dataa(!rreq),
	.datab(!\rd_ptr_msb|counter_reg_bit[4]~q ),
	.datac(!\low_addressa[5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_read_address[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_read_address[5]~5 .extended_lut = "off";
defparam \ram_read_address[5]~5 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \ram_read_address[5]~5 .shared_arith = "off";

dffeas \low_addressa[6] (
	.clk(clock),
	.d(\ram_read_address[6]~6_combout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[6]~q ),
	.prn(vcc));
defparam \low_addressa[6] .is_wysiwyg = "true";
defparam \low_addressa[6] .power_up = "low";

arriaii_lcell_comb \ram_read_address[6]~6 (
	.dataa(!rreq),
	.datab(!\rd_ptr_msb|counter_reg_bit[5]~q ),
	.datac(!\low_addressa[6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_read_address[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_read_address[6]~6 .extended_lut = "off";
defparam \ram_read_address[6]~6 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \ram_read_address[6]~6 .shared_arith = "off";

dffeas \low_addressa[7] (
	.clk(clock),
	.d(\ram_read_address[7]~7_combout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\low_addressa[7]~q ),
	.prn(vcc));
defparam \low_addressa[7] .is_wysiwyg = "true";
defparam \low_addressa[7] .power_up = "low";

arriaii_lcell_comb \ram_read_address[7]~7 (
	.dataa(!rreq),
	.datab(!\rd_ptr_msb|counter_reg_bit[6]~q ),
	.datac(!\low_addressa[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ram_read_address[7]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ram_read_address[7]~7 .extended_lut = "off";
defparam \ram_read_address[7]~7 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \ram_read_address[7]~7 .shared_arith = "off";

arriaii_lcell_comb \_~1 (
	.dataa(!rreq),
	.datab(!\rd_ptr_lsb~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~1 .extended_lut = "off";
defparam \_~1 .lut_mask = 64'h4444444444444444;
defparam \_~1 .shared_arith = "off";

arriaii_lcell_comb \rd_ptr_lsb~0 (
	.dataa(!\rd_ptr_lsb~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rd_ptr_lsb~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_ptr_lsb~0 .extended_lut = "off";
defparam \rd_ptr_lsb~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rd_ptr_lsb~0 .shared_arith = "off";

endmodule

module ddr3_int_altsyncram_u1e1 (
	clock0,
	clock1,
	q_b,
	wren_a,
	clocken1,
	address_a,
	address_b,
	data_a)/* synthesis synthesis_greybox=0 */;
input 	clock0;
input 	clock1;
output 	[143:0] q_b;
input 	wren_a;
input 	clocken1;
input 	[7:0] address_a;
input 	[7:0] address_b;
input 	[143:0] data_a;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a132_PORTBDATAOUT_bus;
wire [143:0] ram_block1a140_PORTBDATAOUT_bus;
wire [143:0] ram_block1a128_PORTBDATAOUT_bus;
wire [143:0] ram_block1a136_PORTBDATAOUT_bus;
wire [143:0] ram_block1a133_PORTBDATAOUT_bus;
wire [143:0] ram_block1a141_PORTBDATAOUT_bus;
wire [143:0] ram_block1a129_PORTBDATAOUT_bus;
wire [143:0] ram_block1a137_PORTBDATAOUT_bus;
wire [143:0] ram_block1a134_PORTBDATAOUT_bus;
wire [143:0] ram_block1a142_PORTBDATAOUT_bus;
wire [143:0] ram_block1a130_PORTBDATAOUT_bus;
wire [143:0] ram_block1a138_PORTBDATAOUT_bus;
wire [143:0] ram_block1a135_PORTBDATAOUT_bus;
wire [143:0] ram_block1a143_PORTBDATAOUT_bus;
wire [143:0] ram_block1a131_PORTBDATAOUT_bus;
wire [143:0] ram_block1a139_PORTBDATAOUT_bus;
wire [143:0] ram_block1a96_PORTBDATAOUT_bus;
wire [143:0] ram_block1a32_PORTBDATAOUT_bus;
wire [143:0] ram_block1a64_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a97_PORTBDATAOUT_bus;
wire [143:0] ram_block1a33_PORTBDATAOUT_bus;
wire [143:0] ram_block1a65_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a98_PORTBDATAOUT_bus;
wire [143:0] ram_block1a34_PORTBDATAOUT_bus;
wire [143:0] ram_block1a66_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a99_PORTBDATAOUT_bus;
wire [143:0] ram_block1a35_PORTBDATAOUT_bus;
wire [143:0] ram_block1a67_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a100_PORTBDATAOUT_bus;
wire [143:0] ram_block1a36_PORTBDATAOUT_bus;
wire [143:0] ram_block1a68_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a101_PORTBDATAOUT_bus;
wire [143:0] ram_block1a37_PORTBDATAOUT_bus;
wire [143:0] ram_block1a69_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a102_PORTBDATAOUT_bus;
wire [143:0] ram_block1a38_PORTBDATAOUT_bus;
wire [143:0] ram_block1a70_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a103_PORTBDATAOUT_bus;
wire [143:0] ram_block1a39_PORTBDATAOUT_bus;
wire [143:0] ram_block1a71_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a104_PORTBDATAOUT_bus;
wire [143:0] ram_block1a40_PORTBDATAOUT_bus;
wire [143:0] ram_block1a72_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a105_PORTBDATAOUT_bus;
wire [143:0] ram_block1a41_PORTBDATAOUT_bus;
wire [143:0] ram_block1a73_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a106_PORTBDATAOUT_bus;
wire [143:0] ram_block1a42_PORTBDATAOUT_bus;
wire [143:0] ram_block1a74_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a107_PORTBDATAOUT_bus;
wire [143:0] ram_block1a43_PORTBDATAOUT_bus;
wire [143:0] ram_block1a75_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a108_PORTBDATAOUT_bus;
wire [143:0] ram_block1a44_PORTBDATAOUT_bus;
wire [143:0] ram_block1a76_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a109_PORTBDATAOUT_bus;
wire [143:0] ram_block1a45_PORTBDATAOUT_bus;
wire [143:0] ram_block1a77_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a110_PORTBDATAOUT_bus;
wire [143:0] ram_block1a46_PORTBDATAOUT_bus;
wire [143:0] ram_block1a78_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a111_PORTBDATAOUT_bus;
wire [143:0] ram_block1a47_PORTBDATAOUT_bus;
wire [143:0] ram_block1a79_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a112_PORTBDATAOUT_bus;
wire [143:0] ram_block1a48_PORTBDATAOUT_bus;
wire [143:0] ram_block1a80_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a113_PORTBDATAOUT_bus;
wire [143:0] ram_block1a49_PORTBDATAOUT_bus;
wire [143:0] ram_block1a81_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a114_PORTBDATAOUT_bus;
wire [143:0] ram_block1a50_PORTBDATAOUT_bus;
wire [143:0] ram_block1a82_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a115_PORTBDATAOUT_bus;
wire [143:0] ram_block1a51_PORTBDATAOUT_bus;
wire [143:0] ram_block1a83_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a116_PORTBDATAOUT_bus;
wire [143:0] ram_block1a52_PORTBDATAOUT_bus;
wire [143:0] ram_block1a84_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a117_PORTBDATAOUT_bus;
wire [143:0] ram_block1a53_PORTBDATAOUT_bus;
wire [143:0] ram_block1a85_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a118_PORTBDATAOUT_bus;
wire [143:0] ram_block1a54_PORTBDATAOUT_bus;
wire [143:0] ram_block1a86_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a119_PORTBDATAOUT_bus;
wire [143:0] ram_block1a55_PORTBDATAOUT_bus;
wire [143:0] ram_block1a87_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a120_PORTBDATAOUT_bus;
wire [143:0] ram_block1a56_PORTBDATAOUT_bus;
wire [143:0] ram_block1a88_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a121_PORTBDATAOUT_bus;
wire [143:0] ram_block1a57_PORTBDATAOUT_bus;
wire [143:0] ram_block1a89_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a122_PORTBDATAOUT_bus;
wire [143:0] ram_block1a58_PORTBDATAOUT_bus;
wire [143:0] ram_block1a90_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a123_PORTBDATAOUT_bus;
wire [143:0] ram_block1a59_PORTBDATAOUT_bus;
wire [143:0] ram_block1a91_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a124_PORTBDATAOUT_bus;
wire [143:0] ram_block1a60_PORTBDATAOUT_bus;
wire [143:0] ram_block1a92_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a125_PORTBDATAOUT_bus;
wire [143:0] ram_block1a61_PORTBDATAOUT_bus;
wire [143:0] ram_block1a93_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a126_PORTBDATAOUT_bus;
wire [143:0] ram_block1a62_PORTBDATAOUT_bus;
wire [143:0] ram_block1a94_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a127_PORTBDATAOUT_bus;
wire [143:0] ram_block1a63_PORTBDATAOUT_bus;
wire [143:0] ram_block1a95_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;

assign q_b[132] = ram_block1a132_PORTBDATAOUT_bus[0];

assign q_b[140] = ram_block1a140_PORTBDATAOUT_bus[0];

assign q_b[128] = ram_block1a128_PORTBDATAOUT_bus[0];

assign q_b[136] = ram_block1a136_PORTBDATAOUT_bus[0];

assign q_b[133] = ram_block1a133_PORTBDATAOUT_bus[0];

assign q_b[141] = ram_block1a141_PORTBDATAOUT_bus[0];

assign q_b[129] = ram_block1a129_PORTBDATAOUT_bus[0];

assign q_b[137] = ram_block1a137_PORTBDATAOUT_bus[0];

assign q_b[134] = ram_block1a134_PORTBDATAOUT_bus[0];

assign q_b[142] = ram_block1a142_PORTBDATAOUT_bus[0];

assign q_b[130] = ram_block1a130_PORTBDATAOUT_bus[0];

assign q_b[138] = ram_block1a138_PORTBDATAOUT_bus[0];

assign q_b[135] = ram_block1a135_PORTBDATAOUT_bus[0];

assign q_b[143] = ram_block1a143_PORTBDATAOUT_bus[0];

assign q_b[131] = ram_block1a131_PORTBDATAOUT_bus[0];

assign q_b[139] = ram_block1a139_PORTBDATAOUT_bus[0];

assign q_b[96] = ram_block1a96_PORTBDATAOUT_bus[0];

assign q_b[32] = ram_block1a32_PORTBDATAOUT_bus[0];

assign q_b[64] = ram_block1a64_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[97] = ram_block1a97_PORTBDATAOUT_bus[0];

assign q_b[33] = ram_block1a33_PORTBDATAOUT_bus[0];

assign q_b[65] = ram_block1a65_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[98] = ram_block1a98_PORTBDATAOUT_bus[0];

assign q_b[34] = ram_block1a34_PORTBDATAOUT_bus[0];

assign q_b[66] = ram_block1a66_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[99] = ram_block1a99_PORTBDATAOUT_bus[0];

assign q_b[35] = ram_block1a35_PORTBDATAOUT_bus[0];

assign q_b[67] = ram_block1a67_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[100] = ram_block1a100_PORTBDATAOUT_bus[0];

assign q_b[36] = ram_block1a36_PORTBDATAOUT_bus[0];

assign q_b[68] = ram_block1a68_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[101] = ram_block1a101_PORTBDATAOUT_bus[0];

assign q_b[37] = ram_block1a37_PORTBDATAOUT_bus[0];

assign q_b[69] = ram_block1a69_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[102] = ram_block1a102_PORTBDATAOUT_bus[0];

assign q_b[38] = ram_block1a38_PORTBDATAOUT_bus[0];

assign q_b[70] = ram_block1a70_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[103] = ram_block1a103_PORTBDATAOUT_bus[0];

assign q_b[39] = ram_block1a39_PORTBDATAOUT_bus[0];

assign q_b[71] = ram_block1a71_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[104] = ram_block1a104_PORTBDATAOUT_bus[0];

assign q_b[40] = ram_block1a40_PORTBDATAOUT_bus[0];

assign q_b[72] = ram_block1a72_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[105] = ram_block1a105_PORTBDATAOUT_bus[0];

assign q_b[41] = ram_block1a41_PORTBDATAOUT_bus[0];

assign q_b[73] = ram_block1a73_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[106] = ram_block1a106_PORTBDATAOUT_bus[0];

assign q_b[42] = ram_block1a42_PORTBDATAOUT_bus[0];

assign q_b[74] = ram_block1a74_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[107] = ram_block1a107_PORTBDATAOUT_bus[0];

assign q_b[43] = ram_block1a43_PORTBDATAOUT_bus[0];

assign q_b[75] = ram_block1a75_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[108] = ram_block1a108_PORTBDATAOUT_bus[0];

assign q_b[44] = ram_block1a44_PORTBDATAOUT_bus[0];

assign q_b[76] = ram_block1a76_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[109] = ram_block1a109_PORTBDATAOUT_bus[0];

assign q_b[45] = ram_block1a45_PORTBDATAOUT_bus[0];

assign q_b[77] = ram_block1a77_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[110] = ram_block1a110_PORTBDATAOUT_bus[0];

assign q_b[46] = ram_block1a46_PORTBDATAOUT_bus[0];

assign q_b[78] = ram_block1a78_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[111] = ram_block1a111_PORTBDATAOUT_bus[0];

assign q_b[47] = ram_block1a47_PORTBDATAOUT_bus[0];

assign q_b[79] = ram_block1a79_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[112] = ram_block1a112_PORTBDATAOUT_bus[0];

assign q_b[48] = ram_block1a48_PORTBDATAOUT_bus[0];

assign q_b[80] = ram_block1a80_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[113] = ram_block1a113_PORTBDATAOUT_bus[0];

assign q_b[49] = ram_block1a49_PORTBDATAOUT_bus[0];

assign q_b[81] = ram_block1a81_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[114] = ram_block1a114_PORTBDATAOUT_bus[0];

assign q_b[50] = ram_block1a50_PORTBDATAOUT_bus[0];

assign q_b[82] = ram_block1a82_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[115] = ram_block1a115_PORTBDATAOUT_bus[0];

assign q_b[51] = ram_block1a51_PORTBDATAOUT_bus[0];

assign q_b[83] = ram_block1a83_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[116] = ram_block1a116_PORTBDATAOUT_bus[0];

assign q_b[52] = ram_block1a52_PORTBDATAOUT_bus[0];

assign q_b[84] = ram_block1a84_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[117] = ram_block1a117_PORTBDATAOUT_bus[0];

assign q_b[53] = ram_block1a53_PORTBDATAOUT_bus[0];

assign q_b[85] = ram_block1a85_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[118] = ram_block1a118_PORTBDATAOUT_bus[0];

assign q_b[54] = ram_block1a54_PORTBDATAOUT_bus[0];

assign q_b[86] = ram_block1a86_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[119] = ram_block1a119_PORTBDATAOUT_bus[0];

assign q_b[55] = ram_block1a55_PORTBDATAOUT_bus[0];

assign q_b[87] = ram_block1a87_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[120] = ram_block1a120_PORTBDATAOUT_bus[0];

assign q_b[56] = ram_block1a56_PORTBDATAOUT_bus[0];

assign q_b[88] = ram_block1a88_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[121] = ram_block1a121_PORTBDATAOUT_bus[0];

assign q_b[57] = ram_block1a57_PORTBDATAOUT_bus[0];

assign q_b[89] = ram_block1a89_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[122] = ram_block1a122_PORTBDATAOUT_bus[0];

assign q_b[58] = ram_block1a58_PORTBDATAOUT_bus[0];

assign q_b[90] = ram_block1a90_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[123] = ram_block1a123_PORTBDATAOUT_bus[0];

assign q_b[59] = ram_block1a59_PORTBDATAOUT_bus[0];

assign q_b[91] = ram_block1a91_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[124] = ram_block1a124_PORTBDATAOUT_bus[0];

assign q_b[60] = ram_block1a60_PORTBDATAOUT_bus[0];

assign q_b[92] = ram_block1a92_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[125] = ram_block1a125_PORTBDATAOUT_bus[0];

assign q_b[61] = ram_block1a61_PORTBDATAOUT_bus[0];

assign q_b[93] = ram_block1a93_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[126] = ram_block1a126_PORTBDATAOUT_bus[0];

assign q_b[62] = ram_block1a62_PORTBDATAOUT_bus[0];

assign q_b[94] = ram_block1a94_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[127] = ram_block1a127_PORTBDATAOUT_bus[0];

assign q_b[63] = ram_block1a63_PORTBDATAOUT_bus[0];

assign q_b[95] = ram_block1a95_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

arriaii_ram_block ram_block1a132(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[132]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a132_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a132.clk0_core_clock_enable = "ena0";
defparam ram_block1a132.clk0_input_clock_enable = "ena2";
defparam ram_block1a132.clk1_core_clock_enable = "ena3";
defparam ram_block1a132.clk1_input_clock_enable = "ena3";
defparam ram_block1a132.clk1_output_clock_enable = "ena1";
defparam ram_block1a132.clock_duty_cycle_dependence = "on";
defparam ram_block1a132.data_interleave_offset_in_bits = 1;
defparam ram_block1a132.data_interleave_width_in_bits = 1;
defparam ram_block1a132.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a132.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a132.operation_mode = "dual_port";
defparam ram_block1a132.port_a_address_clear = "none";
defparam ram_block1a132.port_a_address_width = 8;
defparam ram_block1a132.port_a_data_out_clear = "none";
defparam ram_block1a132.port_a_data_out_clock = "none";
defparam ram_block1a132.port_a_data_width = 1;
defparam ram_block1a132.port_a_first_address = 0;
defparam ram_block1a132.port_a_first_bit_number = 132;
defparam ram_block1a132.port_a_last_address = 255;
defparam ram_block1a132.port_a_logical_ram_depth = 256;
defparam ram_block1a132.port_a_logical_ram_width = 144;
defparam ram_block1a132.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a132.port_b_address_clear = "none";
defparam ram_block1a132.port_b_address_clock = "clock1";
defparam ram_block1a132.port_b_address_width = 8;
defparam ram_block1a132.port_b_data_out_clear = "none";
defparam ram_block1a132.port_b_data_out_clock = "clock1";
defparam ram_block1a132.port_b_data_width = 1;
defparam ram_block1a132.port_b_first_address = 0;
defparam ram_block1a132.port_b_first_bit_number = 132;
defparam ram_block1a132.port_b_last_address = 255;
defparam ram_block1a132.port_b_logical_ram_depth = 256;
defparam ram_block1a132.port_b_logical_ram_width = 144;
defparam ram_block1a132.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a132.port_b_read_enable_clock = "clock1";
defparam ram_block1a132.ram_block_type = "auto";

arriaii_ram_block ram_block1a140(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[140]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a140_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a140.clk0_core_clock_enable = "ena0";
defparam ram_block1a140.clk0_input_clock_enable = "ena2";
defparam ram_block1a140.clk1_core_clock_enable = "ena3";
defparam ram_block1a140.clk1_input_clock_enable = "ena3";
defparam ram_block1a140.clk1_output_clock_enable = "ena1";
defparam ram_block1a140.clock_duty_cycle_dependence = "on";
defparam ram_block1a140.data_interleave_offset_in_bits = 1;
defparam ram_block1a140.data_interleave_width_in_bits = 1;
defparam ram_block1a140.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a140.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a140.operation_mode = "dual_port";
defparam ram_block1a140.port_a_address_clear = "none";
defparam ram_block1a140.port_a_address_width = 8;
defparam ram_block1a140.port_a_data_out_clear = "none";
defparam ram_block1a140.port_a_data_out_clock = "none";
defparam ram_block1a140.port_a_data_width = 1;
defparam ram_block1a140.port_a_first_address = 0;
defparam ram_block1a140.port_a_first_bit_number = 140;
defparam ram_block1a140.port_a_last_address = 255;
defparam ram_block1a140.port_a_logical_ram_depth = 256;
defparam ram_block1a140.port_a_logical_ram_width = 144;
defparam ram_block1a140.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a140.port_b_address_clear = "none";
defparam ram_block1a140.port_b_address_clock = "clock1";
defparam ram_block1a140.port_b_address_width = 8;
defparam ram_block1a140.port_b_data_out_clear = "none";
defparam ram_block1a140.port_b_data_out_clock = "clock1";
defparam ram_block1a140.port_b_data_width = 1;
defparam ram_block1a140.port_b_first_address = 0;
defparam ram_block1a140.port_b_first_bit_number = 140;
defparam ram_block1a140.port_b_last_address = 255;
defparam ram_block1a140.port_b_logical_ram_depth = 256;
defparam ram_block1a140.port_b_logical_ram_width = 144;
defparam ram_block1a140.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a140.port_b_read_enable_clock = "clock1";
defparam ram_block1a140.ram_block_type = "auto";

arriaii_ram_block ram_block1a128(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[128]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a128_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a128.clk0_core_clock_enable = "ena0";
defparam ram_block1a128.clk0_input_clock_enable = "ena2";
defparam ram_block1a128.clk1_core_clock_enable = "ena3";
defparam ram_block1a128.clk1_input_clock_enable = "ena3";
defparam ram_block1a128.clk1_output_clock_enable = "ena1";
defparam ram_block1a128.clock_duty_cycle_dependence = "on";
defparam ram_block1a128.data_interleave_offset_in_bits = 1;
defparam ram_block1a128.data_interleave_width_in_bits = 1;
defparam ram_block1a128.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a128.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a128.operation_mode = "dual_port";
defparam ram_block1a128.port_a_address_clear = "none";
defparam ram_block1a128.port_a_address_width = 8;
defparam ram_block1a128.port_a_data_out_clear = "none";
defparam ram_block1a128.port_a_data_out_clock = "none";
defparam ram_block1a128.port_a_data_width = 1;
defparam ram_block1a128.port_a_first_address = 0;
defparam ram_block1a128.port_a_first_bit_number = 128;
defparam ram_block1a128.port_a_last_address = 255;
defparam ram_block1a128.port_a_logical_ram_depth = 256;
defparam ram_block1a128.port_a_logical_ram_width = 144;
defparam ram_block1a128.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a128.port_b_address_clear = "none";
defparam ram_block1a128.port_b_address_clock = "clock1";
defparam ram_block1a128.port_b_address_width = 8;
defparam ram_block1a128.port_b_data_out_clear = "none";
defparam ram_block1a128.port_b_data_out_clock = "clock1";
defparam ram_block1a128.port_b_data_width = 1;
defparam ram_block1a128.port_b_first_address = 0;
defparam ram_block1a128.port_b_first_bit_number = 128;
defparam ram_block1a128.port_b_last_address = 255;
defparam ram_block1a128.port_b_logical_ram_depth = 256;
defparam ram_block1a128.port_b_logical_ram_width = 144;
defparam ram_block1a128.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a128.port_b_read_enable_clock = "clock1";
defparam ram_block1a128.ram_block_type = "auto";

arriaii_ram_block ram_block1a136(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[136]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a136_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a136.clk0_core_clock_enable = "ena0";
defparam ram_block1a136.clk0_input_clock_enable = "ena2";
defparam ram_block1a136.clk1_core_clock_enable = "ena3";
defparam ram_block1a136.clk1_input_clock_enable = "ena3";
defparam ram_block1a136.clk1_output_clock_enable = "ena1";
defparam ram_block1a136.clock_duty_cycle_dependence = "on";
defparam ram_block1a136.data_interleave_offset_in_bits = 1;
defparam ram_block1a136.data_interleave_width_in_bits = 1;
defparam ram_block1a136.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a136.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a136.operation_mode = "dual_port";
defparam ram_block1a136.port_a_address_clear = "none";
defparam ram_block1a136.port_a_address_width = 8;
defparam ram_block1a136.port_a_data_out_clear = "none";
defparam ram_block1a136.port_a_data_out_clock = "none";
defparam ram_block1a136.port_a_data_width = 1;
defparam ram_block1a136.port_a_first_address = 0;
defparam ram_block1a136.port_a_first_bit_number = 136;
defparam ram_block1a136.port_a_last_address = 255;
defparam ram_block1a136.port_a_logical_ram_depth = 256;
defparam ram_block1a136.port_a_logical_ram_width = 144;
defparam ram_block1a136.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a136.port_b_address_clear = "none";
defparam ram_block1a136.port_b_address_clock = "clock1";
defparam ram_block1a136.port_b_address_width = 8;
defparam ram_block1a136.port_b_data_out_clear = "none";
defparam ram_block1a136.port_b_data_out_clock = "clock1";
defparam ram_block1a136.port_b_data_width = 1;
defparam ram_block1a136.port_b_first_address = 0;
defparam ram_block1a136.port_b_first_bit_number = 136;
defparam ram_block1a136.port_b_last_address = 255;
defparam ram_block1a136.port_b_logical_ram_depth = 256;
defparam ram_block1a136.port_b_logical_ram_width = 144;
defparam ram_block1a136.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a136.port_b_read_enable_clock = "clock1";
defparam ram_block1a136.ram_block_type = "auto";

arriaii_ram_block ram_block1a133(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[133]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a133_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a133.clk0_core_clock_enable = "ena0";
defparam ram_block1a133.clk0_input_clock_enable = "ena2";
defparam ram_block1a133.clk1_core_clock_enable = "ena3";
defparam ram_block1a133.clk1_input_clock_enable = "ena3";
defparam ram_block1a133.clk1_output_clock_enable = "ena1";
defparam ram_block1a133.clock_duty_cycle_dependence = "on";
defparam ram_block1a133.data_interleave_offset_in_bits = 1;
defparam ram_block1a133.data_interleave_width_in_bits = 1;
defparam ram_block1a133.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a133.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a133.operation_mode = "dual_port";
defparam ram_block1a133.port_a_address_clear = "none";
defparam ram_block1a133.port_a_address_width = 8;
defparam ram_block1a133.port_a_data_out_clear = "none";
defparam ram_block1a133.port_a_data_out_clock = "none";
defparam ram_block1a133.port_a_data_width = 1;
defparam ram_block1a133.port_a_first_address = 0;
defparam ram_block1a133.port_a_first_bit_number = 133;
defparam ram_block1a133.port_a_last_address = 255;
defparam ram_block1a133.port_a_logical_ram_depth = 256;
defparam ram_block1a133.port_a_logical_ram_width = 144;
defparam ram_block1a133.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a133.port_b_address_clear = "none";
defparam ram_block1a133.port_b_address_clock = "clock1";
defparam ram_block1a133.port_b_address_width = 8;
defparam ram_block1a133.port_b_data_out_clear = "none";
defparam ram_block1a133.port_b_data_out_clock = "clock1";
defparam ram_block1a133.port_b_data_width = 1;
defparam ram_block1a133.port_b_first_address = 0;
defparam ram_block1a133.port_b_first_bit_number = 133;
defparam ram_block1a133.port_b_last_address = 255;
defparam ram_block1a133.port_b_logical_ram_depth = 256;
defparam ram_block1a133.port_b_logical_ram_width = 144;
defparam ram_block1a133.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a133.port_b_read_enable_clock = "clock1";
defparam ram_block1a133.ram_block_type = "auto";

arriaii_ram_block ram_block1a141(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[141]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a141_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a141.clk0_core_clock_enable = "ena0";
defparam ram_block1a141.clk0_input_clock_enable = "ena2";
defparam ram_block1a141.clk1_core_clock_enable = "ena3";
defparam ram_block1a141.clk1_input_clock_enable = "ena3";
defparam ram_block1a141.clk1_output_clock_enable = "ena1";
defparam ram_block1a141.clock_duty_cycle_dependence = "on";
defparam ram_block1a141.data_interleave_offset_in_bits = 1;
defparam ram_block1a141.data_interleave_width_in_bits = 1;
defparam ram_block1a141.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a141.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a141.operation_mode = "dual_port";
defparam ram_block1a141.port_a_address_clear = "none";
defparam ram_block1a141.port_a_address_width = 8;
defparam ram_block1a141.port_a_data_out_clear = "none";
defparam ram_block1a141.port_a_data_out_clock = "none";
defparam ram_block1a141.port_a_data_width = 1;
defparam ram_block1a141.port_a_first_address = 0;
defparam ram_block1a141.port_a_first_bit_number = 141;
defparam ram_block1a141.port_a_last_address = 255;
defparam ram_block1a141.port_a_logical_ram_depth = 256;
defparam ram_block1a141.port_a_logical_ram_width = 144;
defparam ram_block1a141.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a141.port_b_address_clear = "none";
defparam ram_block1a141.port_b_address_clock = "clock1";
defparam ram_block1a141.port_b_address_width = 8;
defparam ram_block1a141.port_b_data_out_clear = "none";
defparam ram_block1a141.port_b_data_out_clock = "clock1";
defparam ram_block1a141.port_b_data_width = 1;
defparam ram_block1a141.port_b_first_address = 0;
defparam ram_block1a141.port_b_first_bit_number = 141;
defparam ram_block1a141.port_b_last_address = 255;
defparam ram_block1a141.port_b_logical_ram_depth = 256;
defparam ram_block1a141.port_b_logical_ram_width = 144;
defparam ram_block1a141.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a141.port_b_read_enable_clock = "clock1";
defparam ram_block1a141.ram_block_type = "auto";

arriaii_ram_block ram_block1a129(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[129]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a129_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a129.clk0_core_clock_enable = "ena0";
defparam ram_block1a129.clk0_input_clock_enable = "ena2";
defparam ram_block1a129.clk1_core_clock_enable = "ena3";
defparam ram_block1a129.clk1_input_clock_enable = "ena3";
defparam ram_block1a129.clk1_output_clock_enable = "ena1";
defparam ram_block1a129.clock_duty_cycle_dependence = "on";
defparam ram_block1a129.data_interleave_offset_in_bits = 1;
defparam ram_block1a129.data_interleave_width_in_bits = 1;
defparam ram_block1a129.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a129.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a129.operation_mode = "dual_port";
defparam ram_block1a129.port_a_address_clear = "none";
defparam ram_block1a129.port_a_address_width = 8;
defparam ram_block1a129.port_a_data_out_clear = "none";
defparam ram_block1a129.port_a_data_out_clock = "none";
defparam ram_block1a129.port_a_data_width = 1;
defparam ram_block1a129.port_a_first_address = 0;
defparam ram_block1a129.port_a_first_bit_number = 129;
defparam ram_block1a129.port_a_last_address = 255;
defparam ram_block1a129.port_a_logical_ram_depth = 256;
defparam ram_block1a129.port_a_logical_ram_width = 144;
defparam ram_block1a129.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a129.port_b_address_clear = "none";
defparam ram_block1a129.port_b_address_clock = "clock1";
defparam ram_block1a129.port_b_address_width = 8;
defparam ram_block1a129.port_b_data_out_clear = "none";
defparam ram_block1a129.port_b_data_out_clock = "clock1";
defparam ram_block1a129.port_b_data_width = 1;
defparam ram_block1a129.port_b_first_address = 0;
defparam ram_block1a129.port_b_first_bit_number = 129;
defparam ram_block1a129.port_b_last_address = 255;
defparam ram_block1a129.port_b_logical_ram_depth = 256;
defparam ram_block1a129.port_b_logical_ram_width = 144;
defparam ram_block1a129.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a129.port_b_read_enable_clock = "clock1";
defparam ram_block1a129.ram_block_type = "auto";

arriaii_ram_block ram_block1a137(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[137]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a137_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a137.clk0_core_clock_enable = "ena0";
defparam ram_block1a137.clk0_input_clock_enable = "ena2";
defparam ram_block1a137.clk1_core_clock_enable = "ena3";
defparam ram_block1a137.clk1_input_clock_enable = "ena3";
defparam ram_block1a137.clk1_output_clock_enable = "ena1";
defparam ram_block1a137.clock_duty_cycle_dependence = "on";
defparam ram_block1a137.data_interleave_offset_in_bits = 1;
defparam ram_block1a137.data_interleave_width_in_bits = 1;
defparam ram_block1a137.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a137.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a137.operation_mode = "dual_port";
defparam ram_block1a137.port_a_address_clear = "none";
defparam ram_block1a137.port_a_address_width = 8;
defparam ram_block1a137.port_a_data_out_clear = "none";
defparam ram_block1a137.port_a_data_out_clock = "none";
defparam ram_block1a137.port_a_data_width = 1;
defparam ram_block1a137.port_a_first_address = 0;
defparam ram_block1a137.port_a_first_bit_number = 137;
defparam ram_block1a137.port_a_last_address = 255;
defparam ram_block1a137.port_a_logical_ram_depth = 256;
defparam ram_block1a137.port_a_logical_ram_width = 144;
defparam ram_block1a137.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a137.port_b_address_clear = "none";
defparam ram_block1a137.port_b_address_clock = "clock1";
defparam ram_block1a137.port_b_address_width = 8;
defparam ram_block1a137.port_b_data_out_clear = "none";
defparam ram_block1a137.port_b_data_out_clock = "clock1";
defparam ram_block1a137.port_b_data_width = 1;
defparam ram_block1a137.port_b_first_address = 0;
defparam ram_block1a137.port_b_first_bit_number = 137;
defparam ram_block1a137.port_b_last_address = 255;
defparam ram_block1a137.port_b_logical_ram_depth = 256;
defparam ram_block1a137.port_b_logical_ram_width = 144;
defparam ram_block1a137.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a137.port_b_read_enable_clock = "clock1";
defparam ram_block1a137.ram_block_type = "auto";

arriaii_ram_block ram_block1a134(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[134]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a134_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a134.clk0_core_clock_enable = "ena0";
defparam ram_block1a134.clk0_input_clock_enable = "ena2";
defparam ram_block1a134.clk1_core_clock_enable = "ena3";
defparam ram_block1a134.clk1_input_clock_enable = "ena3";
defparam ram_block1a134.clk1_output_clock_enable = "ena1";
defparam ram_block1a134.clock_duty_cycle_dependence = "on";
defparam ram_block1a134.data_interleave_offset_in_bits = 1;
defparam ram_block1a134.data_interleave_width_in_bits = 1;
defparam ram_block1a134.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a134.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a134.operation_mode = "dual_port";
defparam ram_block1a134.port_a_address_clear = "none";
defparam ram_block1a134.port_a_address_width = 8;
defparam ram_block1a134.port_a_data_out_clear = "none";
defparam ram_block1a134.port_a_data_out_clock = "none";
defparam ram_block1a134.port_a_data_width = 1;
defparam ram_block1a134.port_a_first_address = 0;
defparam ram_block1a134.port_a_first_bit_number = 134;
defparam ram_block1a134.port_a_last_address = 255;
defparam ram_block1a134.port_a_logical_ram_depth = 256;
defparam ram_block1a134.port_a_logical_ram_width = 144;
defparam ram_block1a134.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a134.port_b_address_clear = "none";
defparam ram_block1a134.port_b_address_clock = "clock1";
defparam ram_block1a134.port_b_address_width = 8;
defparam ram_block1a134.port_b_data_out_clear = "none";
defparam ram_block1a134.port_b_data_out_clock = "clock1";
defparam ram_block1a134.port_b_data_width = 1;
defparam ram_block1a134.port_b_first_address = 0;
defparam ram_block1a134.port_b_first_bit_number = 134;
defparam ram_block1a134.port_b_last_address = 255;
defparam ram_block1a134.port_b_logical_ram_depth = 256;
defparam ram_block1a134.port_b_logical_ram_width = 144;
defparam ram_block1a134.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a134.port_b_read_enable_clock = "clock1";
defparam ram_block1a134.ram_block_type = "auto";

arriaii_ram_block ram_block1a142(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[142]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a142_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a142.clk0_core_clock_enable = "ena0";
defparam ram_block1a142.clk0_input_clock_enable = "ena2";
defparam ram_block1a142.clk1_core_clock_enable = "ena3";
defparam ram_block1a142.clk1_input_clock_enable = "ena3";
defparam ram_block1a142.clk1_output_clock_enable = "ena1";
defparam ram_block1a142.clock_duty_cycle_dependence = "on";
defparam ram_block1a142.data_interleave_offset_in_bits = 1;
defparam ram_block1a142.data_interleave_width_in_bits = 1;
defparam ram_block1a142.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a142.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a142.operation_mode = "dual_port";
defparam ram_block1a142.port_a_address_clear = "none";
defparam ram_block1a142.port_a_address_width = 8;
defparam ram_block1a142.port_a_data_out_clear = "none";
defparam ram_block1a142.port_a_data_out_clock = "none";
defparam ram_block1a142.port_a_data_width = 1;
defparam ram_block1a142.port_a_first_address = 0;
defparam ram_block1a142.port_a_first_bit_number = 142;
defparam ram_block1a142.port_a_last_address = 255;
defparam ram_block1a142.port_a_logical_ram_depth = 256;
defparam ram_block1a142.port_a_logical_ram_width = 144;
defparam ram_block1a142.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a142.port_b_address_clear = "none";
defparam ram_block1a142.port_b_address_clock = "clock1";
defparam ram_block1a142.port_b_address_width = 8;
defparam ram_block1a142.port_b_data_out_clear = "none";
defparam ram_block1a142.port_b_data_out_clock = "clock1";
defparam ram_block1a142.port_b_data_width = 1;
defparam ram_block1a142.port_b_first_address = 0;
defparam ram_block1a142.port_b_first_bit_number = 142;
defparam ram_block1a142.port_b_last_address = 255;
defparam ram_block1a142.port_b_logical_ram_depth = 256;
defparam ram_block1a142.port_b_logical_ram_width = 144;
defparam ram_block1a142.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a142.port_b_read_enable_clock = "clock1";
defparam ram_block1a142.ram_block_type = "auto";

arriaii_ram_block ram_block1a130(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[130]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a130_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a130.clk0_core_clock_enable = "ena0";
defparam ram_block1a130.clk0_input_clock_enable = "ena2";
defparam ram_block1a130.clk1_core_clock_enable = "ena3";
defparam ram_block1a130.clk1_input_clock_enable = "ena3";
defparam ram_block1a130.clk1_output_clock_enable = "ena1";
defparam ram_block1a130.clock_duty_cycle_dependence = "on";
defparam ram_block1a130.data_interleave_offset_in_bits = 1;
defparam ram_block1a130.data_interleave_width_in_bits = 1;
defparam ram_block1a130.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a130.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a130.operation_mode = "dual_port";
defparam ram_block1a130.port_a_address_clear = "none";
defparam ram_block1a130.port_a_address_width = 8;
defparam ram_block1a130.port_a_data_out_clear = "none";
defparam ram_block1a130.port_a_data_out_clock = "none";
defparam ram_block1a130.port_a_data_width = 1;
defparam ram_block1a130.port_a_first_address = 0;
defparam ram_block1a130.port_a_first_bit_number = 130;
defparam ram_block1a130.port_a_last_address = 255;
defparam ram_block1a130.port_a_logical_ram_depth = 256;
defparam ram_block1a130.port_a_logical_ram_width = 144;
defparam ram_block1a130.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a130.port_b_address_clear = "none";
defparam ram_block1a130.port_b_address_clock = "clock1";
defparam ram_block1a130.port_b_address_width = 8;
defparam ram_block1a130.port_b_data_out_clear = "none";
defparam ram_block1a130.port_b_data_out_clock = "clock1";
defparam ram_block1a130.port_b_data_width = 1;
defparam ram_block1a130.port_b_first_address = 0;
defparam ram_block1a130.port_b_first_bit_number = 130;
defparam ram_block1a130.port_b_last_address = 255;
defparam ram_block1a130.port_b_logical_ram_depth = 256;
defparam ram_block1a130.port_b_logical_ram_width = 144;
defparam ram_block1a130.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a130.port_b_read_enable_clock = "clock1";
defparam ram_block1a130.ram_block_type = "auto";

arriaii_ram_block ram_block1a138(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[138]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a138_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a138.clk0_core_clock_enable = "ena0";
defparam ram_block1a138.clk0_input_clock_enable = "ena2";
defparam ram_block1a138.clk1_core_clock_enable = "ena3";
defparam ram_block1a138.clk1_input_clock_enable = "ena3";
defparam ram_block1a138.clk1_output_clock_enable = "ena1";
defparam ram_block1a138.clock_duty_cycle_dependence = "on";
defparam ram_block1a138.data_interleave_offset_in_bits = 1;
defparam ram_block1a138.data_interleave_width_in_bits = 1;
defparam ram_block1a138.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a138.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a138.operation_mode = "dual_port";
defparam ram_block1a138.port_a_address_clear = "none";
defparam ram_block1a138.port_a_address_width = 8;
defparam ram_block1a138.port_a_data_out_clear = "none";
defparam ram_block1a138.port_a_data_out_clock = "none";
defparam ram_block1a138.port_a_data_width = 1;
defparam ram_block1a138.port_a_first_address = 0;
defparam ram_block1a138.port_a_first_bit_number = 138;
defparam ram_block1a138.port_a_last_address = 255;
defparam ram_block1a138.port_a_logical_ram_depth = 256;
defparam ram_block1a138.port_a_logical_ram_width = 144;
defparam ram_block1a138.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a138.port_b_address_clear = "none";
defparam ram_block1a138.port_b_address_clock = "clock1";
defparam ram_block1a138.port_b_address_width = 8;
defparam ram_block1a138.port_b_data_out_clear = "none";
defparam ram_block1a138.port_b_data_out_clock = "clock1";
defparam ram_block1a138.port_b_data_width = 1;
defparam ram_block1a138.port_b_first_address = 0;
defparam ram_block1a138.port_b_first_bit_number = 138;
defparam ram_block1a138.port_b_last_address = 255;
defparam ram_block1a138.port_b_logical_ram_depth = 256;
defparam ram_block1a138.port_b_logical_ram_width = 144;
defparam ram_block1a138.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a138.port_b_read_enable_clock = "clock1";
defparam ram_block1a138.ram_block_type = "auto";

arriaii_ram_block ram_block1a135(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[135]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a135_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a135.clk0_core_clock_enable = "ena0";
defparam ram_block1a135.clk0_input_clock_enable = "ena2";
defparam ram_block1a135.clk1_core_clock_enable = "ena3";
defparam ram_block1a135.clk1_input_clock_enable = "ena3";
defparam ram_block1a135.clk1_output_clock_enable = "ena1";
defparam ram_block1a135.clock_duty_cycle_dependence = "on";
defparam ram_block1a135.data_interleave_offset_in_bits = 1;
defparam ram_block1a135.data_interleave_width_in_bits = 1;
defparam ram_block1a135.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a135.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a135.operation_mode = "dual_port";
defparam ram_block1a135.port_a_address_clear = "none";
defparam ram_block1a135.port_a_address_width = 8;
defparam ram_block1a135.port_a_data_out_clear = "none";
defparam ram_block1a135.port_a_data_out_clock = "none";
defparam ram_block1a135.port_a_data_width = 1;
defparam ram_block1a135.port_a_first_address = 0;
defparam ram_block1a135.port_a_first_bit_number = 135;
defparam ram_block1a135.port_a_last_address = 255;
defparam ram_block1a135.port_a_logical_ram_depth = 256;
defparam ram_block1a135.port_a_logical_ram_width = 144;
defparam ram_block1a135.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a135.port_b_address_clear = "none";
defparam ram_block1a135.port_b_address_clock = "clock1";
defparam ram_block1a135.port_b_address_width = 8;
defparam ram_block1a135.port_b_data_out_clear = "none";
defparam ram_block1a135.port_b_data_out_clock = "clock1";
defparam ram_block1a135.port_b_data_width = 1;
defparam ram_block1a135.port_b_first_address = 0;
defparam ram_block1a135.port_b_first_bit_number = 135;
defparam ram_block1a135.port_b_last_address = 255;
defparam ram_block1a135.port_b_logical_ram_depth = 256;
defparam ram_block1a135.port_b_logical_ram_width = 144;
defparam ram_block1a135.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a135.port_b_read_enable_clock = "clock1";
defparam ram_block1a135.ram_block_type = "auto";

arriaii_ram_block ram_block1a143(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[143]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a143_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a143.clk0_core_clock_enable = "ena0";
defparam ram_block1a143.clk0_input_clock_enable = "ena2";
defparam ram_block1a143.clk1_core_clock_enable = "ena3";
defparam ram_block1a143.clk1_input_clock_enable = "ena3";
defparam ram_block1a143.clk1_output_clock_enable = "ena1";
defparam ram_block1a143.clock_duty_cycle_dependence = "on";
defparam ram_block1a143.data_interleave_offset_in_bits = 1;
defparam ram_block1a143.data_interleave_width_in_bits = 1;
defparam ram_block1a143.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a143.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a143.operation_mode = "dual_port";
defparam ram_block1a143.port_a_address_clear = "none";
defparam ram_block1a143.port_a_address_width = 8;
defparam ram_block1a143.port_a_data_out_clear = "none";
defparam ram_block1a143.port_a_data_out_clock = "none";
defparam ram_block1a143.port_a_data_width = 1;
defparam ram_block1a143.port_a_first_address = 0;
defparam ram_block1a143.port_a_first_bit_number = 143;
defparam ram_block1a143.port_a_last_address = 255;
defparam ram_block1a143.port_a_logical_ram_depth = 256;
defparam ram_block1a143.port_a_logical_ram_width = 144;
defparam ram_block1a143.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a143.port_b_address_clear = "none";
defparam ram_block1a143.port_b_address_clock = "clock1";
defparam ram_block1a143.port_b_address_width = 8;
defparam ram_block1a143.port_b_data_out_clear = "none";
defparam ram_block1a143.port_b_data_out_clock = "clock1";
defparam ram_block1a143.port_b_data_width = 1;
defparam ram_block1a143.port_b_first_address = 0;
defparam ram_block1a143.port_b_first_bit_number = 143;
defparam ram_block1a143.port_b_last_address = 255;
defparam ram_block1a143.port_b_logical_ram_depth = 256;
defparam ram_block1a143.port_b_logical_ram_width = 144;
defparam ram_block1a143.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a143.port_b_read_enable_clock = "clock1";
defparam ram_block1a143.ram_block_type = "auto";

arriaii_ram_block ram_block1a131(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[131]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a131_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a131.clk0_core_clock_enable = "ena0";
defparam ram_block1a131.clk0_input_clock_enable = "ena2";
defparam ram_block1a131.clk1_core_clock_enable = "ena3";
defparam ram_block1a131.clk1_input_clock_enable = "ena3";
defparam ram_block1a131.clk1_output_clock_enable = "ena1";
defparam ram_block1a131.clock_duty_cycle_dependence = "on";
defparam ram_block1a131.data_interleave_offset_in_bits = 1;
defparam ram_block1a131.data_interleave_width_in_bits = 1;
defparam ram_block1a131.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a131.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a131.operation_mode = "dual_port";
defparam ram_block1a131.port_a_address_clear = "none";
defparam ram_block1a131.port_a_address_width = 8;
defparam ram_block1a131.port_a_data_out_clear = "none";
defparam ram_block1a131.port_a_data_out_clock = "none";
defparam ram_block1a131.port_a_data_width = 1;
defparam ram_block1a131.port_a_first_address = 0;
defparam ram_block1a131.port_a_first_bit_number = 131;
defparam ram_block1a131.port_a_last_address = 255;
defparam ram_block1a131.port_a_logical_ram_depth = 256;
defparam ram_block1a131.port_a_logical_ram_width = 144;
defparam ram_block1a131.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a131.port_b_address_clear = "none";
defparam ram_block1a131.port_b_address_clock = "clock1";
defparam ram_block1a131.port_b_address_width = 8;
defparam ram_block1a131.port_b_data_out_clear = "none";
defparam ram_block1a131.port_b_data_out_clock = "clock1";
defparam ram_block1a131.port_b_data_width = 1;
defparam ram_block1a131.port_b_first_address = 0;
defparam ram_block1a131.port_b_first_bit_number = 131;
defparam ram_block1a131.port_b_last_address = 255;
defparam ram_block1a131.port_b_logical_ram_depth = 256;
defparam ram_block1a131.port_b_logical_ram_width = 144;
defparam ram_block1a131.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a131.port_b_read_enable_clock = "clock1";
defparam ram_block1a131.ram_block_type = "auto";

arriaii_ram_block ram_block1a139(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[139]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a139_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a139.clk0_core_clock_enable = "ena0";
defparam ram_block1a139.clk0_input_clock_enable = "ena2";
defparam ram_block1a139.clk1_core_clock_enable = "ena3";
defparam ram_block1a139.clk1_input_clock_enable = "ena3";
defparam ram_block1a139.clk1_output_clock_enable = "ena1";
defparam ram_block1a139.clock_duty_cycle_dependence = "on";
defparam ram_block1a139.data_interleave_offset_in_bits = 1;
defparam ram_block1a139.data_interleave_width_in_bits = 1;
defparam ram_block1a139.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a139.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a139.operation_mode = "dual_port";
defparam ram_block1a139.port_a_address_clear = "none";
defparam ram_block1a139.port_a_address_width = 8;
defparam ram_block1a139.port_a_data_out_clear = "none";
defparam ram_block1a139.port_a_data_out_clock = "none";
defparam ram_block1a139.port_a_data_width = 1;
defparam ram_block1a139.port_a_first_address = 0;
defparam ram_block1a139.port_a_first_bit_number = 139;
defparam ram_block1a139.port_a_last_address = 255;
defparam ram_block1a139.port_a_logical_ram_depth = 256;
defparam ram_block1a139.port_a_logical_ram_width = 144;
defparam ram_block1a139.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a139.port_b_address_clear = "none";
defparam ram_block1a139.port_b_address_clock = "clock1";
defparam ram_block1a139.port_b_address_width = 8;
defparam ram_block1a139.port_b_data_out_clear = "none";
defparam ram_block1a139.port_b_data_out_clock = "clock1";
defparam ram_block1a139.port_b_data_width = 1;
defparam ram_block1a139.port_b_first_address = 0;
defparam ram_block1a139.port_b_first_bit_number = 139;
defparam ram_block1a139.port_b_last_address = 255;
defparam ram_block1a139.port_b_logical_ram_depth = 256;
defparam ram_block1a139.port_b_logical_ram_width = 144;
defparam ram_block1a139.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a139.port_b_read_enable_clock = "clock1";
defparam ram_block1a139.ram_block_type = "auto";

arriaii_ram_block ram_block1a96(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[96]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a96_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a96.clk0_core_clock_enable = "ena0";
defparam ram_block1a96.clk0_input_clock_enable = "ena2";
defparam ram_block1a96.clk1_core_clock_enable = "ena3";
defparam ram_block1a96.clk1_input_clock_enable = "ena3";
defparam ram_block1a96.clk1_output_clock_enable = "ena1";
defparam ram_block1a96.clock_duty_cycle_dependence = "on";
defparam ram_block1a96.data_interleave_offset_in_bits = 1;
defparam ram_block1a96.data_interleave_width_in_bits = 1;
defparam ram_block1a96.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a96.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a96.operation_mode = "dual_port";
defparam ram_block1a96.port_a_address_clear = "none";
defparam ram_block1a96.port_a_address_width = 8;
defparam ram_block1a96.port_a_data_out_clear = "none";
defparam ram_block1a96.port_a_data_out_clock = "none";
defparam ram_block1a96.port_a_data_width = 1;
defparam ram_block1a96.port_a_first_address = 0;
defparam ram_block1a96.port_a_first_bit_number = 96;
defparam ram_block1a96.port_a_last_address = 255;
defparam ram_block1a96.port_a_logical_ram_depth = 256;
defparam ram_block1a96.port_a_logical_ram_width = 144;
defparam ram_block1a96.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a96.port_b_address_clear = "none";
defparam ram_block1a96.port_b_address_clock = "clock1";
defparam ram_block1a96.port_b_address_width = 8;
defparam ram_block1a96.port_b_data_out_clear = "none";
defparam ram_block1a96.port_b_data_out_clock = "clock1";
defparam ram_block1a96.port_b_data_width = 1;
defparam ram_block1a96.port_b_first_address = 0;
defparam ram_block1a96.port_b_first_bit_number = 96;
defparam ram_block1a96.port_b_last_address = 255;
defparam ram_block1a96.port_b_logical_ram_depth = 256;
defparam ram_block1a96.port_b_logical_ram_width = 144;
defparam ram_block1a96.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a96.port_b_read_enable_clock = "clock1";
defparam ram_block1a96.ram_block_type = "auto";

arriaii_ram_block ram_block1a32(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[32]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a32_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a32.clk0_core_clock_enable = "ena0";
defparam ram_block1a32.clk0_input_clock_enable = "ena2";
defparam ram_block1a32.clk1_core_clock_enable = "ena3";
defparam ram_block1a32.clk1_input_clock_enable = "ena3";
defparam ram_block1a32.clk1_output_clock_enable = "ena1";
defparam ram_block1a32.clock_duty_cycle_dependence = "on";
defparam ram_block1a32.data_interleave_offset_in_bits = 1;
defparam ram_block1a32.data_interleave_width_in_bits = 1;
defparam ram_block1a32.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a32.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a32.operation_mode = "dual_port";
defparam ram_block1a32.port_a_address_clear = "none";
defparam ram_block1a32.port_a_address_width = 8;
defparam ram_block1a32.port_a_data_out_clear = "none";
defparam ram_block1a32.port_a_data_out_clock = "none";
defparam ram_block1a32.port_a_data_width = 1;
defparam ram_block1a32.port_a_first_address = 0;
defparam ram_block1a32.port_a_first_bit_number = 32;
defparam ram_block1a32.port_a_last_address = 255;
defparam ram_block1a32.port_a_logical_ram_depth = 256;
defparam ram_block1a32.port_a_logical_ram_width = 144;
defparam ram_block1a32.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a32.port_b_address_clear = "none";
defparam ram_block1a32.port_b_address_clock = "clock1";
defparam ram_block1a32.port_b_address_width = 8;
defparam ram_block1a32.port_b_data_out_clear = "none";
defparam ram_block1a32.port_b_data_out_clock = "clock1";
defparam ram_block1a32.port_b_data_width = 1;
defparam ram_block1a32.port_b_first_address = 0;
defparam ram_block1a32.port_b_first_bit_number = 32;
defparam ram_block1a32.port_b_last_address = 255;
defparam ram_block1a32.port_b_logical_ram_depth = 256;
defparam ram_block1a32.port_b_logical_ram_width = 144;
defparam ram_block1a32.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a32.port_b_read_enable_clock = "clock1";
defparam ram_block1a32.ram_block_type = "auto";

arriaii_ram_block ram_block1a64(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[64]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a64_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a64.clk0_core_clock_enable = "ena0";
defparam ram_block1a64.clk0_input_clock_enable = "ena2";
defparam ram_block1a64.clk1_core_clock_enable = "ena3";
defparam ram_block1a64.clk1_input_clock_enable = "ena3";
defparam ram_block1a64.clk1_output_clock_enable = "ena1";
defparam ram_block1a64.clock_duty_cycle_dependence = "on";
defparam ram_block1a64.data_interleave_offset_in_bits = 1;
defparam ram_block1a64.data_interleave_width_in_bits = 1;
defparam ram_block1a64.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a64.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a64.operation_mode = "dual_port";
defparam ram_block1a64.port_a_address_clear = "none";
defparam ram_block1a64.port_a_address_width = 8;
defparam ram_block1a64.port_a_data_out_clear = "none";
defparam ram_block1a64.port_a_data_out_clock = "none";
defparam ram_block1a64.port_a_data_width = 1;
defparam ram_block1a64.port_a_first_address = 0;
defparam ram_block1a64.port_a_first_bit_number = 64;
defparam ram_block1a64.port_a_last_address = 255;
defparam ram_block1a64.port_a_logical_ram_depth = 256;
defparam ram_block1a64.port_a_logical_ram_width = 144;
defparam ram_block1a64.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a64.port_b_address_clear = "none";
defparam ram_block1a64.port_b_address_clock = "clock1";
defparam ram_block1a64.port_b_address_width = 8;
defparam ram_block1a64.port_b_data_out_clear = "none";
defparam ram_block1a64.port_b_data_out_clock = "clock1";
defparam ram_block1a64.port_b_data_width = 1;
defparam ram_block1a64.port_b_first_address = 0;
defparam ram_block1a64.port_b_first_bit_number = 64;
defparam ram_block1a64.port_b_last_address = 255;
defparam ram_block1a64.port_b_logical_ram_depth = 256;
defparam ram_block1a64.port_b_logical_ram_width = 144;
defparam ram_block1a64.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a64.port_b_read_enable_clock = "clock1";
defparam ram_block1a64.ram_block_type = "auto";

arriaii_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena2";
defparam ram_block1a0.clk1_core_clock_enable = "ena3";
defparam ram_block1a0.clk1_input_clock_enable = "ena3";
defparam ram_block1a0.clk1_output_clock_enable = "ena1";
defparam ram_block1a0.clock_duty_cycle_dependence = "on";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 8;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 255;
defparam ram_block1a0.port_a_logical_ram_depth = 256;
defparam ram_block1a0.port_a_logical_ram_width = 144;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 8;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock1";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 255;
defparam ram_block1a0.port_b_logical_ram_depth = 256;
defparam ram_block1a0.port_b_logical_ram_width = 144;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

arriaii_ram_block ram_block1a97(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[97]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a97_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a97.clk0_core_clock_enable = "ena0";
defparam ram_block1a97.clk0_input_clock_enable = "ena2";
defparam ram_block1a97.clk1_core_clock_enable = "ena3";
defparam ram_block1a97.clk1_input_clock_enable = "ena3";
defparam ram_block1a97.clk1_output_clock_enable = "ena1";
defparam ram_block1a97.clock_duty_cycle_dependence = "on";
defparam ram_block1a97.data_interleave_offset_in_bits = 1;
defparam ram_block1a97.data_interleave_width_in_bits = 1;
defparam ram_block1a97.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a97.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a97.operation_mode = "dual_port";
defparam ram_block1a97.port_a_address_clear = "none";
defparam ram_block1a97.port_a_address_width = 8;
defparam ram_block1a97.port_a_data_out_clear = "none";
defparam ram_block1a97.port_a_data_out_clock = "none";
defparam ram_block1a97.port_a_data_width = 1;
defparam ram_block1a97.port_a_first_address = 0;
defparam ram_block1a97.port_a_first_bit_number = 97;
defparam ram_block1a97.port_a_last_address = 255;
defparam ram_block1a97.port_a_logical_ram_depth = 256;
defparam ram_block1a97.port_a_logical_ram_width = 144;
defparam ram_block1a97.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a97.port_b_address_clear = "none";
defparam ram_block1a97.port_b_address_clock = "clock1";
defparam ram_block1a97.port_b_address_width = 8;
defparam ram_block1a97.port_b_data_out_clear = "none";
defparam ram_block1a97.port_b_data_out_clock = "clock1";
defparam ram_block1a97.port_b_data_width = 1;
defparam ram_block1a97.port_b_first_address = 0;
defparam ram_block1a97.port_b_first_bit_number = 97;
defparam ram_block1a97.port_b_last_address = 255;
defparam ram_block1a97.port_b_logical_ram_depth = 256;
defparam ram_block1a97.port_b_logical_ram_width = 144;
defparam ram_block1a97.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a97.port_b_read_enable_clock = "clock1";
defparam ram_block1a97.ram_block_type = "auto";

arriaii_ram_block ram_block1a33(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[33]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a33_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a33.clk0_core_clock_enable = "ena0";
defparam ram_block1a33.clk0_input_clock_enable = "ena2";
defparam ram_block1a33.clk1_core_clock_enable = "ena3";
defparam ram_block1a33.clk1_input_clock_enable = "ena3";
defparam ram_block1a33.clk1_output_clock_enable = "ena1";
defparam ram_block1a33.clock_duty_cycle_dependence = "on";
defparam ram_block1a33.data_interleave_offset_in_bits = 1;
defparam ram_block1a33.data_interleave_width_in_bits = 1;
defparam ram_block1a33.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a33.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a33.operation_mode = "dual_port";
defparam ram_block1a33.port_a_address_clear = "none";
defparam ram_block1a33.port_a_address_width = 8;
defparam ram_block1a33.port_a_data_out_clear = "none";
defparam ram_block1a33.port_a_data_out_clock = "none";
defparam ram_block1a33.port_a_data_width = 1;
defparam ram_block1a33.port_a_first_address = 0;
defparam ram_block1a33.port_a_first_bit_number = 33;
defparam ram_block1a33.port_a_last_address = 255;
defparam ram_block1a33.port_a_logical_ram_depth = 256;
defparam ram_block1a33.port_a_logical_ram_width = 144;
defparam ram_block1a33.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a33.port_b_address_clear = "none";
defparam ram_block1a33.port_b_address_clock = "clock1";
defparam ram_block1a33.port_b_address_width = 8;
defparam ram_block1a33.port_b_data_out_clear = "none";
defparam ram_block1a33.port_b_data_out_clock = "clock1";
defparam ram_block1a33.port_b_data_width = 1;
defparam ram_block1a33.port_b_first_address = 0;
defparam ram_block1a33.port_b_first_bit_number = 33;
defparam ram_block1a33.port_b_last_address = 255;
defparam ram_block1a33.port_b_logical_ram_depth = 256;
defparam ram_block1a33.port_b_logical_ram_width = 144;
defparam ram_block1a33.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a33.port_b_read_enable_clock = "clock1";
defparam ram_block1a33.ram_block_type = "auto";

arriaii_ram_block ram_block1a65(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[65]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a65_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a65.clk0_core_clock_enable = "ena0";
defparam ram_block1a65.clk0_input_clock_enable = "ena2";
defparam ram_block1a65.clk1_core_clock_enable = "ena3";
defparam ram_block1a65.clk1_input_clock_enable = "ena3";
defparam ram_block1a65.clk1_output_clock_enable = "ena1";
defparam ram_block1a65.clock_duty_cycle_dependence = "on";
defparam ram_block1a65.data_interleave_offset_in_bits = 1;
defparam ram_block1a65.data_interleave_width_in_bits = 1;
defparam ram_block1a65.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a65.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a65.operation_mode = "dual_port";
defparam ram_block1a65.port_a_address_clear = "none";
defparam ram_block1a65.port_a_address_width = 8;
defparam ram_block1a65.port_a_data_out_clear = "none";
defparam ram_block1a65.port_a_data_out_clock = "none";
defparam ram_block1a65.port_a_data_width = 1;
defparam ram_block1a65.port_a_first_address = 0;
defparam ram_block1a65.port_a_first_bit_number = 65;
defparam ram_block1a65.port_a_last_address = 255;
defparam ram_block1a65.port_a_logical_ram_depth = 256;
defparam ram_block1a65.port_a_logical_ram_width = 144;
defparam ram_block1a65.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a65.port_b_address_clear = "none";
defparam ram_block1a65.port_b_address_clock = "clock1";
defparam ram_block1a65.port_b_address_width = 8;
defparam ram_block1a65.port_b_data_out_clear = "none";
defparam ram_block1a65.port_b_data_out_clock = "clock1";
defparam ram_block1a65.port_b_data_width = 1;
defparam ram_block1a65.port_b_first_address = 0;
defparam ram_block1a65.port_b_first_bit_number = 65;
defparam ram_block1a65.port_b_last_address = 255;
defparam ram_block1a65.port_b_logical_ram_depth = 256;
defparam ram_block1a65.port_b_logical_ram_width = 144;
defparam ram_block1a65.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a65.port_b_read_enable_clock = "clock1";
defparam ram_block1a65.ram_block_type = "auto";

arriaii_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena2";
defparam ram_block1a1.clk1_core_clock_enable = "ena3";
defparam ram_block1a1.clk1_input_clock_enable = "ena3";
defparam ram_block1a1.clk1_output_clock_enable = "ena1";
defparam ram_block1a1.clock_duty_cycle_dependence = "on";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 8;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 255;
defparam ram_block1a1.port_a_logical_ram_depth = 256;
defparam ram_block1a1.port_a_logical_ram_width = 144;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 8;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock1";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 255;
defparam ram_block1a1.port_b_logical_ram_depth = 256;
defparam ram_block1a1.port_b_logical_ram_width = 144;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

arriaii_ram_block ram_block1a98(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[98]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a98_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a98.clk0_core_clock_enable = "ena0";
defparam ram_block1a98.clk0_input_clock_enable = "ena2";
defparam ram_block1a98.clk1_core_clock_enable = "ena3";
defparam ram_block1a98.clk1_input_clock_enable = "ena3";
defparam ram_block1a98.clk1_output_clock_enable = "ena1";
defparam ram_block1a98.clock_duty_cycle_dependence = "on";
defparam ram_block1a98.data_interleave_offset_in_bits = 1;
defparam ram_block1a98.data_interleave_width_in_bits = 1;
defparam ram_block1a98.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a98.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a98.operation_mode = "dual_port";
defparam ram_block1a98.port_a_address_clear = "none";
defparam ram_block1a98.port_a_address_width = 8;
defparam ram_block1a98.port_a_data_out_clear = "none";
defparam ram_block1a98.port_a_data_out_clock = "none";
defparam ram_block1a98.port_a_data_width = 1;
defparam ram_block1a98.port_a_first_address = 0;
defparam ram_block1a98.port_a_first_bit_number = 98;
defparam ram_block1a98.port_a_last_address = 255;
defparam ram_block1a98.port_a_logical_ram_depth = 256;
defparam ram_block1a98.port_a_logical_ram_width = 144;
defparam ram_block1a98.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a98.port_b_address_clear = "none";
defparam ram_block1a98.port_b_address_clock = "clock1";
defparam ram_block1a98.port_b_address_width = 8;
defparam ram_block1a98.port_b_data_out_clear = "none";
defparam ram_block1a98.port_b_data_out_clock = "clock1";
defparam ram_block1a98.port_b_data_width = 1;
defparam ram_block1a98.port_b_first_address = 0;
defparam ram_block1a98.port_b_first_bit_number = 98;
defparam ram_block1a98.port_b_last_address = 255;
defparam ram_block1a98.port_b_logical_ram_depth = 256;
defparam ram_block1a98.port_b_logical_ram_width = 144;
defparam ram_block1a98.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a98.port_b_read_enable_clock = "clock1";
defparam ram_block1a98.ram_block_type = "auto";

arriaii_ram_block ram_block1a34(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[34]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a34_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a34.clk0_core_clock_enable = "ena0";
defparam ram_block1a34.clk0_input_clock_enable = "ena2";
defparam ram_block1a34.clk1_core_clock_enable = "ena3";
defparam ram_block1a34.clk1_input_clock_enable = "ena3";
defparam ram_block1a34.clk1_output_clock_enable = "ena1";
defparam ram_block1a34.clock_duty_cycle_dependence = "on";
defparam ram_block1a34.data_interleave_offset_in_bits = 1;
defparam ram_block1a34.data_interleave_width_in_bits = 1;
defparam ram_block1a34.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a34.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a34.operation_mode = "dual_port";
defparam ram_block1a34.port_a_address_clear = "none";
defparam ram_block1a34.port_a_address_width = 8;
defparam ram_block1a34.port_a_data_out_clear = "none";
defparam ram_block1a34.port_a_data_out_clock = "none";
defparam ram_block1a34.port_a_data_width = 1;
defparam ram_block1a34.port_a_first_address = 0;
defparam ram_block1a34.port_a_first_bit_number = 34;
defparam ram_block1a34.port_a_last_address = 255;
defparam ram_block1a34.port_a_logical_ram_depth = 256;
defparam ram_block1a34.port_a_logical_ram_width = 144;
defparam ram_block1a34.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a34.port_b_address_clear = "none";
defparam ram_block1a34.port_b_address_clock = "clock1";
defparam ram_block1a34.port_b_address_width = 8;
defparam ram_block1a34.port_b_data_out_clear = "none";
defparam ram_block1a34.port_b_data_out_clock = "clock1";
defparam ram_block1a34.port_b_data_width = 1;
defparam ram_block1a34.port_b_first_address = 0;
defparam ram_block1a34.port_b_first_bit_number = 34;
defparam ram_block1a34.port_b_last_address = 255;
defparam ram_block1a34.port_b_logical_ram_depth = 256;
defparam ram_block1a34.port_b_logical_ram_width = 144;
defparam ram_block1a34.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a34.port_b_read_enable_clock = "clock1";
defparam ram_block1a34.ram_block_type = "auto";

arriaii_ram_block ram_block1a66(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[66]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a66_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a66.clk0_core_clock_enable = "ena0";
defparam ram_block1a66.clk0_input_clock_enable = "ena2";
defparam ram_block1a66.clk1_core_clock_enable = "ena3";
defparam ram_block1a66.clk1_input_clock_enable = "ena3";
defparam ram_block1a66.clk1_output_clock_enable = "ena1";
defparam ram_block1a66.clock_duty_cycle_dependence = "on";
defparam ram_block1a66.data_interleave_offset_in_bits = 1;
defparam ram_block1a66.data_interleave_width_in_bits = 1;
defparam ram_block1a66.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a66.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a66.operation_mode = "dual_port";
defparam ram_block1a66.port_a_address_clear = "none";
defparam ram_block1a66.port_a_address_width = 8;
defparam ram_block1a66.port_a_data_out_clear = "none";
defparam ram_block1a66.port_a_data_out_clock = "none";
defparam ram_block1a66.port_a_data_width = 1;
defparam ram_block1a66.port_a_first_address = 0;
defparam ram_block1a66.port_a_first_bit_number = 66;
defparam ram_block1a66.port_a_last_address = 255;
defparam ram_block1a66.port_a_logical_ram_depth = 256;
defparam ram_block1a66.port_a_logical_ram_width = 144;
defparam ram_block1a66.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a66.port_b_address_clear = "none";
defparam ram_block1a66.port_b_address_clock = "clock1";
defparam ram_block1a66.port_b_address_width = 8;
defparam ram_block1a66.port_b_data_out_clear = "none";
defparam ram_block1a66.port_b_data_out_clock = "clock1";
defparam ram_block1a66.port_b_data_width = 1;
defparam ram_block1a66.port_b_first_address = 0;
defparam ram_block1a66.port_b_first_bit_number = 66;
defparam ram_block1a66.port_b_last_address = 255;
defparam ram_block1a66.port_b_logical_ram_depth = 256;
defparam ram_block1a66.port_b_logical_ram_width = 144;
defparam ram_block1a66.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a66.port_b_read_enable_clock = "clock1";
defparam ram_block1a66.ram_block_type = "auto";

arriaii_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena2";
defparam ram_block1a2.clk1_core_clock_enable = "ena3";
defparam ram_block1a2.clk1_input_clock_enable = "ena3";
defparam ram_block1a2.clk1_output_clock_enable = "ena1";
defparam ram_block1a2.clock_duty_cycle_dependence = "on";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 8;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 255;
defparam ram_block1a2.port_a_logical_ram_depth = 256;
defparam ram_block1a2.port_a_logical_ram_width = 144;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 8;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock1";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 255;
defparam ram_block1a2.port_b_logical_ram_depth = 256;
defparam ram_block1a2.port_b_logical_ram_width = 144;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

arriaii_ram_block ram_block1a99(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[99]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a99_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a99.clk0_core_clock_enable = "ena0";
defparam ram_block1a99.clk0_input_clock_enable = "ena2";
defparam ram_block1a99.clk1_core_clock_enable = "ena3";
defparam ram_block1a99.clk1_input_clock_enable = "ena3";
defparam ram_block1a99.clk1_output_clock_enable = "ena1";
defparam ram_block1a99.clock_duty_cycle_dependence = "on";
defparam ram_block1a99.data_interleave_offset_in_bits = 1;
defparam ram_block1a99.data_interleave_width_in_bits = 1;
defparam ram_block1a99.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a99.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a99.operation_mode = "dual_port";
defparam ram_block1a99.port_a_address_clear = "none";
defparam ram_block1a99.port_a_address_width = 8;
defparam ram_block1a99.port_a_data_out_clear = "none";
defparam ram_block1a99.port_a_data_out_clock = "none";
defparam ram_block1a99.port_a_data_width = 1;
defparam ram_block1a99.port_a_first_address = 0;
defparam ram_block1a99.port_a_first_bit_number = 99;
defparam ram_block1a99.port_a_last_address = 255;
defparam ram_block1a99.port_a_logical_ram_depth = 256;
defparam ram_block1a99.port_a_logical_ram_width = 144;
defparam ram_block1a99.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a99.port_b_address_clear = "none";
defparam ram_block1a99.port_b_address_clock = "clock1";
defparam ram_block1a99.port_b_address_width = 8;
defparam ram_block1a99.port_b_data_out_clear = "none";
defparam ram_block1a99.port_b_data_out_clock = "clock1";
defparam ram_block1a99.port_b_data_width = 1;
defparam ram_block1a99.port_b_first_address = 0;
defparam ram_block1a99.port_b_first_bit_number = 99;
defparam ram_block1a99.port_b_last_address = 255;
defparam ram_block1a99.port_b_logical_ram_depth = 256;
defparam ram_block1a99.port_b_logical_ram_width = 144;
defparam ram_block1a99.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a99.port_b_read_enable_clock = "clock1";
defparam ram_block1a99.ram_block_type = "auto";

arriaii_ram_block ram_block1a35(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[35]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a35_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a35.clk0_core_clock_enable = "ena0";
defparam ram_block1a35.clk0_input_clock_enable = "ena2";
defparam ram_block1a35.clk1_core_clock_enable = "ena3";
defparam ram_block1a35.clk1_input_clock_enable = "ena3";
defparam ram_block1a35.clk1_output_clock_enable = "ena1";
defparam ram_block1a35.clock_duty_cycle_dependence = "on";
defparam ram_block1a35.data_interleave_offset_in_bits = 1;
defparam ram_block1a35.data_interleave_width_in_bits = 1;
defparam ram_block1a35.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a35.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a35.operation_mode = "dual_port";
defparam ram_block1a35.port_a_address_clear = "none";
defparam ram_block1a35.port_a_address_width = 8;
defparam ram_block1a35.port_a_data_out_clear = "none";
defparam ram_block1a35.port_a_data_out_clock = "none";
defparam ram_block1a35.port_a_data_width = 1;
defparam ram_block1a35.port_a_first_address = 0;
defparam ram_block1a35.port_a_first_bit_number = 35;
defparam ram_block1a35.port_a_last_address = 255;
defparam ram_block1a35.port_a_logical_ram_depth = 256;
defparam ram_block1a35.port_a_logical_ram_width = 144;
defparam ram_block1a35.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a35.port_b_address_clear = "none";
defparam ram_block1a35.port_b_address_clock = "clock1";
defparam ram_block1a35.port_b_address_width = 8;
defparam ram_block1a35.port_b_data_out_clear = "none";
defparam ram_block1a35.port_b_data_out_clock = "clock1";
defparam ram_block1a35.port_b_data_width = 1;
defparam ram_block1a35.port_b_first_address = 0;
defparam ram_block1a35.port_b_first_bit_number = 35;
defparam ram_block1a35.port_b_last_address = 255;
defparam ram_block1a35.port_b_logical_ram_depth = 256;
defparam ram_block1a35.port_b_logical_ram_width = 144;
defparam ram_block1a35.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a35.port_b_read_enable_clock = "clock1";
defparam ram_block1a35.ram_block_type = "auto";

arriaii_ram_block ram_block1a67(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[67]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a67_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a67.clk0_core_clock_enable = "ena0";
defparam ram_block1a67.clk0_input_clock_enable = "ena2";
defparam ram_block1a67.clk1_core_clock_enable = "ena3";
defparam ram_block1a67.clk1_input_clock_enable = "ena3";
defparam ram_block1a67.clk1_output_clock_enable = "ena1";
defparam ram_block1a67.clock_duty_cycle_dependence = "on";
defparam ram_block1a67.data_interleave_offset_in_bits = 1;
defparam ram_block1a67.data_interleave_width_in_bits = 1;
defparam ram_block1a67.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a67.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a67.operation_mode = "dual_port";
defparam ram_block1a67.port_a_address_clear = "none";
defparam ram_block1a67.port_a_address_width = 8;
defparam ram_block1a67.port_a_data_out_clear = "none";
defparam ram_block1a67.port_a_data_out_clock = "none";
defparam ram_block1a67.port_a_data_width = 1;
defparam ram_block1a67.port_a_first_address = 0;
defparam ram_block1a67.port_a_first_bit_number = 67;
defparam ram_block1a67.port_a_last_address = 255;
defparam ram_block1a67.port_a_logical_ram_depth = 256;
defparam ram_block1a67.port_a_logical_ram_width = 144;
defparam ram_block1a67.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a67.port_b_address_clear = "none";
defparam ram_block1a67.port_b_address_clock = "clock1";
defparam ram_block1a67.port_b_address_width = 8;
defparam ram_block1a67.port_b_data_out_clear = "none";
defparam ram_block1a67.port_b_data_out_clock = "clock1";
defparam ram_block1a67.port_b_data_width = 1;
defparam ram_block1a67.port_b_first_address = 0;
defparam ram_block1a67.port_b_first_bit_number = 67;
defparam ram_block1a67.port_b_last_address = 255;
defparam ram_block1a67.port_b_logical_ram_depth = 256;
defparam ram_block1a67.port_b_logical_ram_width = 144;
defparam ram_block1a67.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a67.port_b_read_enable_clock = "clock1";
defparam ram_block1a67.ram_block_type = "auto";

arriaii_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena2";
defparam ram_block1a3.clk1_core_clock_enable = "ena3";
defparam ram_block1a3.clk1_input_clock_enable = "ena3";
defparam ram_block1a3.clk1_output_clock_enable = "ena1";
defparam ram_block1a3.clock_duty_cycle_dependence = "on";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 8;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 255;
defparam ram_block1a3.port_a_logical_ram_depth = 256;
defparam ram_block1a3.port_a_logical_ram_width = 144;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 8;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock1";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 255;
defparam ram_block1a3.port_b_logical_ram_depth = 256;
defparam ram_block1a3.port_b_logical_ram_width = 144;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

arriaii_ram_block ram_block1a100(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[100]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a100_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a100.clk0_core_clock_enable = "ena0";
defparam ram_block1a100.clk0_input_clock_enable = "ena2";
defparam ram_block1a100.clk1_core_clock_enable = "ena3";
defparam ram_block1a100.clk1_input_clock_enable = "ena3";
defparam ram_block1a100.clk1_output_clock_enable = "ena1";
defparam ram_block1a100.clock_duty_cycle_dependence = "on";
defparam ram_block1a100.data_interleave_offset_in_bits = 1;
defparam ram_block1a100.data_interleave_width_in_bits = 1;
defparam ram_block1a100.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a100.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a100.operation_mode = "dual_port";
defparam ram_block1a100.port_a_address_clear = "none";
defparam ram_block1a100.port_a_address_width = 8;
defparam ram_block1a100.port_a_data_out_clear = "none";
defparam ram_block1a100.port_a_data_out_clock = "none";
defparam ram_block1a100.port_a_data_width = 1;
defparam ram_block1a100.port_a_first_address = 0;
defparam ram_block1a100.port_a_first_bit_number = 100;
defparam ram_block1a100.port_a_last_address = 255;
defparam ram_block1a100.port_a_logical_ram_depth = 256;
defparam ram_block1a100.port_a_logical_ram_width = 144;
defparam ram_block1a100.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a100.port_b_address_clear = "none";
defparam ram_block1a100.port_b_address_clock = "clock1";
defparam ram_block1a100.port_b_address_width = 8;
defparam ram_block1a100.port_b_data_out_clear = "none";
defparam ram_block1a100.port_b_data_out_clock = "clock1";
defparam ram_block1a100.port_b_data_width = 1;
defparam ram_block1a100.port_b_first_address = 0;
defparam ram_block1a100.port_b_first_bit_number = 100;
defparam ram_block1a100.port_b_last_address = 255;
defparam ram_block1a100.port_b_logical_ram_depth = 256;
defparam ram_block1a100.port_b_logical_ram_width = 144;
defparam ram_block1a100.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a100.port_b_read_enable_clock = "clock1";
defparam ram_block1a100.ram_block_type = "auto";

arriaii_ram_block ram_block1a36(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[36]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a36_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a36.clk0_core_clock_enable = "ena0";
defparam ram_block1a36.clk0_input_clock_enable = "ena2";
defparam ram_block1a36.clk1_core_clock_enable = "ena3";
defparam ram_block1a36.clk1_input_clock_enable = "ena3";
defparam ram_block1a36.clk1_output_clock_enable = "ena1";
defparam ram_block1a36.clock_duty_cycle_dependence = "on";
defparam ram_block1a36.data_interleave_offset_in_bits = 1;
defparam ram_block1a36.data_interleave_width_in_bits = 1;
defparam ram_block1a36.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a36.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a36.operation_mode = "dual_port";
defparam ram_block1a36.port_a_address_clear = "none";
defparam ram_block1a36.port_a_address_width = 8;
defparam ram_block1a36.port_a_data_out_clear = "none";
defparam ram_block1a36.port_a_data_out_clock = "none";
defparam ram_block1a36.port_a_data_width = 1;
defparam ram_block1a36.port_a_first_address = 0;
defparam ram_block1a36.port_a_first_bit_number = 36;
defparam ram_block1a36.port_a_last_address = 255;
defparam ram_block1a36.port_a_logical_ram_depth = 256;
defparam ram_block1a36.port_a_logical_ram_width = 144;
defparam ram_block1a36.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a36.port_b_address_clear = "none";
defparam ram_block1a36.port_b_address_clock = "clock1";
defparam ram_block1a36.port_b_address_width = 8;
defparam ram_block1a36.port_b_data_out_clear = "none";
defparam ram_block1a36.port_b_data_out_clock = "clock1";
defparam ram_block1a36.port_b_data_width = 1;
defparam ram_block1a36.port_b_first_address = 0;
defparam ram_block1a36.port_b_first_bit_number = 36;
defparam ram_block1a36.port_b_last_address = 255;
defparam ram_block1a36.port_b_logical_ram_depth = 256;
defparam ram_block1a36.port_b_logical_ram_width = 144;
defparam ram_block1a36.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a36.port_b_read_enable_clock = "clock1";
defparam ram_block1a36.ram_block_type = "auto";

arriaii_ram_block ram_block1a68(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[68]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a68_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a68.clk0_core_clock_enable = "ena0";
defparam ram_block1a68.clk0_input_clock_enable = "ena2";
defparam ram_block1a68.clk1_core_clock_enable = "ena3";
defparam ram_block1a68.clk1_input_clock_enable = "ena3";
defparam ram_block1a68.clk1_output_clock_enable = "ena1";
defparam ram_block1a68.clock_duty_cycle_dependence = "on";
defparam ram_block1a68.data_interleave_offset_in_bits = 1;
defparam ram_block1a68.data_interleave_width_in_bits = 1;
defparam ram_block1a68.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a68.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a68.operation_mode = "dual_port";
defparam ram_block1a68.port_a_address_clear = "none";
defparam ram_block1a68.port_a_address_width = 8;
defparam ram_block1a68.port_a_data_out_clear = "none";
defparam ram_block1a68.port_a_data_out_clock = "none";
defparam ram_block1a68.port_a_data_width = 1;
defparam ram_block1a68.port_a_first_address = 0;
defparam ram_block1a68.port_a_first_bit_number = 68;
defparam ram_block1a68.port_a_last_address = 255;
defparam ram_block1a68.port_a_logical_ram_depth = 256;
defparam ram_block1a68.port_a_logical_ram_width = 144;
defparam ram_block1a68.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a68.port_b_address_clear = "none";
defparam ram_block1a68.port_b_address_clock = "clock1";
defparam ram_block1a68.port_b_address_width = 8;
defparam ram_block1a68.port_b_data_out_clear = "none";
defparam ram_block1a68.port_b_data_out_clock = "clock1";
defparam ram_block1a68.port_b_data_width = 1;
defparam ram_block1a68.port_b_first_address = 0;
defparam ram_block1a68.port_b_first_bit_number = 68;
defparam ram_block1a68.port_b_last_address = 255;
defparam ram_block1a68.port_b_logical_ram_depth = 256;
defparam ram_block1a68.port_b_logical_ram_width = 144;
defparam ram_block1a68.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a68.port_b_read_enable_clock = "clock1";
defparam ram_block1a68.ram_block_type = "auto";

arriaii_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena2";
defparam ram_block1a4.clk1_core_clock_enable = "ena3";
defparam ram_block1a4.clk1_input_clock_enable = "ena3";
defparam ram_block1a4.clk1_output_clock_enable = "ena1";
defparam ram_block1a4.clock_duty_cycle_dependence = "on";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 8;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 255;
defparam ram_block1a4.port_a_logical_ram_depth = 256;
defparam ram_block1a4.port_a_logical_ram_width = 144;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 8;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock1";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 255;
defparam ram_block1a4.port_b_logical_ram_depth = 256;
defparam ram_block1a4.port_b_logical_ram_width = 144;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

arriaii_ram_block ram_block1a101(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[101]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a101_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a101.clk0_core_clock_enable = "ena0";
defparam ram_block1a101.clk0_input_clock_enable = "ena2";
defparam ram_block1a101.clk1_core_clock_enable = "ena3";
defparam ram_block1a101.clk1_input_clock_enable = "ena3";
defparam ram_block1a101.clk1_output_clock_enable = "ena1";
defparam ram_block1a101.clock_duty_cycle_dependence = "on";
defparam ram_block1a101.data_interleave_offset_in_bits = 1;
defparam ram_block1a101.data_interleave_width_in_bits = 1;
defparam ram_block1a101.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a101.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a101.operation_mode = "dual_port";
defparam ram_block1a101.port_a_address_clear = "none";
defparam ram_block1a101.port_a_address_width = 8;
defparam ram_block1a101.port_a_data_out_clear = "none";
defparam ram_block1a101.port_a_data_out_clock = "none";
defparam ram_block1a101.port_a_data_width = 1;
defparam ram_block1a101.port_a_first_address = 0;
defparam ram_block1a101.port_a_first_bit_number = 101;
defparam ram_block1a101.port_a_last_address = 255;
defparam ram_block1a101.port_a_logical_ram_depth = 256;
defparam ram_block1a101.port_a_logical_ram_width = 144;
defparam ram_block1a101.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a101.port_b_address_clear = "none";
defparam ram_block1a101.port_b_address_clock = "clock1";
defparam ram_block1a101.port_b_address_width = 8;
defparam ram_block1a101.port_b_data_out_clear = "none";
defparam ram_block1a101.port_b_data_out_clock = "clock1";
defparam ram_block1a101.port_b_data_width = 1;
defparam ram_block1a101.port_b_first_address = 0;
defparam ram_block1a101.port_b_first_bit_number = 101;
defparam ram_block1a101.port_b_last_address = 255;
defparam ram_block1a101.port_b_logical_ram_depth = 256;
defparam ram_block1a101.port_b_logical_ram_width = 144;
defparam ram_block1a101.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a101.port_b_read_enable_clock = "clock1";
defparam ram_block1a101.ram_block_type = "auto";

arriaii_ram_block ram_block1a37(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[37]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a37_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a37.clk0_core_clock_enable = "ena0";
defparam ram_block1a37.clk0_input_clock_enable = "ena2";
defparam ram_block1a37.clk1_core_clock_enable = "ena3";
defparam ram_block1a37.clk1_input_clock_enable = "ena3";
defparam ram_block1a37.clk1_output_clock_enable = "ena1";
defparam ram_block1a37.clock_duty_cycle_dependence = "on";
defparam ram_block1a37.data_interleave_offset_in_bits = 1;
defparam ram_block1a37.data_interleave_width_in_bits = 1;
defparam ram_block1a37.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a37.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a37.operation_mode = "dual_port";
defparam ram_block1a37.port_a_address_clear = "none";
defparam ram_block1a37.port_a_address_width = 8;
defparam ram_block1a37.port_a_data_out_clear = "none";
defparam ram_block1a37.port_a_data_out_clock = "none";
defparam ram_block1a37.port_a_data_width = 1;
defparam ram_block1a37.port_a_first_address = 0;
defparam ram_block1a37.port_a_first_bit_number = 37;
defparam ram_block1a37.port_a_last_address = 255;
defparam ram_block1a37.port_a_logical_ram_depth = 256;
defparam ram_block1a37.port_a_logical_ram_width = 144;
defparam ram_block1a37.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a37.port_b_address_clear = "none";
defparam ram_block1a37.port_b_address_clock = "clock1";
defparam ram_block1a37.port_b_address_width = 8;
defparam ram_block1a37.port_b_data_out_clear = "none";
defparam ram_block1a37.port_b_data_out_clock = "clock1";
defparam ram_block1a37.port_b_data_width = 1;
defparam ram_block1a37.port_b_first_address = 0;
defparam ram_block1a37.port_b_first_bit_number = 37;
defparam ram_block1a37.port_b_last_address = 255;
defparam ram_block1a37.port_b_logical_ram_depth = 256;
defparam ram_block1a37.port_b_logical_ram_width = 144;
defparam ram_block1a37.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a37.port_b_read_enable_clock = "clock1";
defparam ram_block1a37.ram_block_type = "auto";

arriaii_ram_block ram_block1a69(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[69]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a69_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a69.clk0_core_clock_enable = "ena0";
defparam ram_block1a69.clk0_input_clock_enable = "ena2";
defparam ram_block1a69.clk1_core_clock_enable = "ena3";
defparam ram_block1a69.clk1_input_clock_enable = "ena3";
defparam ram_block1a69.clk1_output_clock_enable = "ena1";
defparam ram_block1a69.clock_duty_cycle_dependence = "on";
defparam ram_block1a69.data_interleave_offset_in_bits = 1;
defparam ram_block1a69.data_interleave_width_in_bits = 1;
defparam ram_block1a69.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a69.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a69.operation_mode = "dual_port";
defparam ram_block1a69.port_a_address_clear = "none";
defparam ram_block1a69.port_a_address_width = 8;
defparam ram_block1a69.port_a_data_out_clear = "none";
defparam ram_block1a69.port_a_data_out_clock = "none";
defparam ram_block1a69.port_a_data_width = 1;
defparam ram_block1a69.port_a_first_address = 0;
defparam ram_block1a69.port_a_first_bit_number = 69;
defparam ram_block1a69.port_a_last_address = 255;
defparam ram_block1a69.port_a_logical_ram_depth = 256;
defparam ram_block1a69.port_a_logical_ram_width = 144;
defparam ram_block1a69.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a69.port_b_address_clear = "none";
defparam ram_block1a69.port_b_address_clock = "clock1";
defparam ram_block1a69.port_b_address_width = 8;
defparam ram_block1a69.port_b_data_out_clear = "none";
defparam ram_block1a69.port_b_data_out_clock = "clock1";
defparam ram_block1a69.port_b_data_width = 1;
defparam ram_block1a69.port_b_first_address = 0;
defparam ram_block1a69.port_b_first_bit_number = 69;
defparam ram_block1a69.port_b_last_address = 255;
defparam ram_block1a69.port_b_logical_ram_depth = 256;
defparam ram_block1a69.port_b_logical_ram_width = 144;
defparam ram_block1a69.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a69.port_b_read_enable_clock = "clock1";
defparam ram_block1a69.ram_block_type = "auto";

arriaii_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena2";
defparam ram_block1a5.clk1_core_clock_enable = "ena3";
defparam ram_block1a5.clk1_input_clock_enable = "ena3";
defparam ram_block1a5.clk1_output_clock_enable = "ena1";
defparam ram_block1a5.clock_duty_cycle_dependence = "on";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 8;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 255;
defparam ram_block1a5.port_a_logical_ram_depth = 256;
defparam ram_block1a5.port_a_logical_ram_width = 144;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 8;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 255;
defparam ram_block1a5.port_b_logical_ram_depth = 256;
defparam ram_block1a5.port_b_logical_ram_width = 144;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

arriaii_ram_block ram_block1a102(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[102]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a102_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a102.clk0_core_clock_enable = "ena0";
defparam ram_block1a102.clk0_input_clock_enable = "ena2";
defparam ram_block1a102.clk1_core_clock_enable = "ena3";
defparam ram_block1a102.clk1_input_clock_enable = "ena3";
defparam ram_block1a102.clk1_output_clock_enable = "ena1";
defparam ram_block1a102.clock_duty_cycle_dependence = "on";
defparam ram_block1a102.data_interleave_offset_in_bits = 1;
defparam ram_block1a102.data_interleave_width_in_bits = 1;
defparam ram_block1a102.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a102.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a102.operation_mode = "dual_port";
defparam ram_block1a102.port_a_address_clear = "none";
defparam ram_block1a102.port_a_address_width = 8;
defparam ram_block1a102.port_a_data_out_clear = "none";
defparam ram_block1a102.port_a_data_out_clock = "none";
defparam ram_block1a102.port_a_data_width = 1;
defparam ram_block1a102.port_a_first_address = 0;
defparam ram_block1a102.port_a_first_bit_number = 102;
defparam ram_block1a102.port_a_last_address = 255;
defparam ram_block1a102.port_a_logical_ram_depth = 256;
defparam ram_block1a102.port_a_logical_ram_width = 144;
defparam ram_block1a102.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a102.port_b_address_clear = "none";
defparam ram_block1a102.port_b_address_clock = "clock1";
defparam ram_block1a102.port_b_address_width = 8;
defparam ram_block1a102.port_b_data_out_clear = "none";
defparam ram_block1a102.port_b_data_out_clock = "clock1";
defparam ram_block1a102.port_b_data_width = 1;
defparam ram_block1a102.port_b_first_address = 0;
defparam ram_block1a102.port_b_first_bit_number = 102;
defparam ram_block1a102.port_b_last_address = 255;
defparam ram_block1a102.port_b_logical_ram_depth = 256;
defparam ram_block1a102.port_b_logical_ram_width = 144;
defparam ram_block1a102.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a102.port_b_read_enable_clock = "clock1";
defparam ram_block1a102.ram_block_type = "auto";

arriaii_ram_block ram_block1a38(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[38]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a38_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a38.clk0_core_clock_enable = "ena0";
defparam ram_block1a38.clk0_input_clock_enable = "ena2";
defparam ram_block1a38.clk1_core_clock_enable = "ena3";
defparam ram_block1a38.clk1_input_clock_enable = "ena3";
defparam ram_block1a38.clk1_output_clock_enable = "ena1";
defparam ram_block1a38.clock_duty_cycle_dependence = "on";
defparam ram_block1a38.data_interleave_offset_in_bits = 1;
defparam ram_block1a38.data_interleave_width_in_bits = 1;
defparam ram_block1a38.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a38.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a38.operation_mode = "dual_port";
defparam ram_block1a38.port_a_address_clear = "none";
defparam ram_block1a38.port_a_address_width = 8;
defparam ram_block1a38.port_a_data_out_clear = "none";
defparam ram_block1a38.port_a_data_out_clock = "none";
defparam ram_block1a38.port_a_data_width = 1;
defparam ram_block1a38.port_a_first_address = 0;
defparam ram_block1a38.port_a_first_bit_number = 38;
defparam ram_block1a38.port_a_last_address = 255;
defparam ram_block1a38.port_a_logical_ram_depth = 256;
defparam ram_block1a38.port_a_logical_ram_width = 144;
defparam ram_block1a38.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a38.port_b_address_clear = "none";
defparam ram_block1a38.port_b_address_clock = "clock1";
defparam ram_block1a38.port_b_address_width = 8;
defparam ram_block1a38.port_b_data_out_clear = "none";
defparam ram_block1a38.port_b_data_out_clock = "clock1";
defparam ram_block1a38.port_b_data_width = 1;
defparam ram_block1a38.port_b_first_address = 0;
defparam ram_block1a38.port_b_first_bit_number = 38;
defparam ram_block1a38.port_b_last_address = 255;
defparam ram_block1a38.port_b_logical_ram_depth = 256;
defparam ram_block1a38.port_b_logical_ram_width = 144;
defparam ram_block1a38.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a38.port_b_read_enable_clock = "clock1";
defparam ram_block1a38.ram_block_type = "auto";

arriaii_ram_block ram_block1a70(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[70]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a70_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a70.clk0_core_clock_enable = "ena0";
defparam ram_block1a70.clk0_input_clock_enable = "ena2";
defparam ram_block1a70.clk1_core_clock_enable = "ena3";
defparam ram_block1a70.clk1_input_clock_enable = "ena3";
defparam ram_block1a70.clk1_output_clock_enable = "ena1";
defparam ram_block1a70.clock_duty_cycle_dependence = "on";
defparam ram_block1a70.data_interleave_offset_in_bits = 1;
defparam ram_block1a70.data_interleave_width_in_bits = 1;
defparam ram_block1a70.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a70.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a70.operation_mode = "dual_port";
defparam ram_block1a70.port_a_address_clear = "none";
defparam ram_block1a70.port_a_address_width = 8;
defparam ram_block1a70.port_a_data_out_clear = "none";
defparam ram_block1a70.port_a_data_out_clock = "none";
defparam ram_block1a70.port_a_data_width = 1;
defparam ram_block1a70.port_a_first_address = 0;
defparam ram_block1a70.port_a_first_bit_number = 70;
defparam ram_block1a70.port_a_last_address = 255;
defparam ram_block1a70.port_a_logical_ram_depth = 256;
defparam ram_block1a70.port_a_logical_ram_width = 144;
defparam ram_block1a70.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a70.port_b_address_clear = "none";
defparam ram_block1a70.port_b_address_clock = "clock1";
defparam ram_block1a70.port_b_address_width = 8;
defparam ram_block1a70.port_b_data_out_clear = "none";
defparam ram_block1a70.port_b_data_out_clock = "clock1";
defparam ram_block1a70.port_b_data_width = 1;
defparam ram_block1a70.port_b_first_address = 0;
defparam ram_block1a70.port_b_first_bit_number = 70;
defparam ram_block1a70.port_b_last_address = 255;
defparam ram_block1a70.port_b_logical_ram_depth = 256;
defparam ram_block1a70.port_b_logical_ram_width = 144;
defparam ram_block1a70.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a70.port_b_read_enable_clock = "clock1";
defparam ram_block1a70.ram_block_type = "auto";

arriaii_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena2";
defparam ram_block1a6.clk1_core_clock_enable = "ena3";
defparam ram_block1a6.clk1_input_clock_enable = "ena3";
defparam ram_block1a6.clk1_output_clock_enable = "ena1";
defparam ram_block1a6.clock_duty_cycle_dependence = "on";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 8;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 255;
defparam ram_block1a6.port_a_logical_ram_depth = 256;
defparam ram_block1a6.port_a_logical_ram_width = 144;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 8;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 255;
defparam ram_block1a6.port_b_logical_ram_depth = 256;
defparam ram_block1a6.port_b_logical_ram_width = 144;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

arriaii_ram_block ram_block1a103(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[103]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a103_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a103.clk0_core_clock_enable = "ena0";
defparam ram_block1a103.clk0_input_clock_enable = "ena2";
defparam ram_block1a103.clk1_core_clock_enable = "ena3";
defparam ram_block1a103.clk1_input_clock_enable = "ena3";
defparam ram_block1a103.clk1_output_clock_enable = "ena1";
defparam ram_block1a103.clock_duty_cycle_dependence = "on";
defparam ram_block1a103.data_interleave_offset_in_bits = 1;
defparam ram_block1a103.data_interleave_width_in_bits = 1;
defparam ram_block1a103.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a103.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a103.operation_mode = "dual_port";
defparam ram_block1a103.port_a_address_clear = "none";
defparam ram_block1a103.port_a_address_width = 8;
defparam ram_block1a103.port_a_data_out_clear = "none";
defparam ram_block1a103.port_a_data_out_clock = "none";
defparam ram_block1a103.port_a_data_width = 1;
defparam ram_block1a103.port_a_first_address = 0;
defparam ram_block1a103.port_a_first_bit_number = 103;
defparam ram_block1a103.port_a_last_address = 255;
defparam ram_block1a103.port_a_logical_ram_depth = 256;
defparam ram_block1a103.port_a_logical_ram_width = 144;
defparam ram_block1a103.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a103.port_b_address_clear = "none";
defparam ram_block1a103.port_b_address_clock = "clock1";
defparam ram_block1a103.port_b_address_width = 8;
defparam ram_block1a103.port_b_data_out_clear = "none";
defparam ram_block1a103.port_b_data_out_clock = "clock1";
defparam ram_block1a103.port_b_data_width = 1;
defparam ram_block1a103.port_b_first_address = 0;
defparam ram_block1a103.port_b_first_bit_number = 103;
defparam ram_block1a103.port_b_last_address = 255;
defparam ram_block1a103.port_b_logical_ram_depth = 256;
defparam ram_block1a103.port_b_logical_ram_width = 144;
defparam ram_block1a103.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a103.port_b_read_enable_clock = "clock1";
defparam ram_block1a103.ram_block_type = "auto";

arriaii_ram_block ram_block1a39(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[39]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a39_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a39.clk0_core_clock_enable = "ena0";
defparam ram_block1a39.clk0_input_clock_enable = "ena2";
defparam ram_block1a39.clk1_core_clock_enable = "ena3";
defparam ram_block1a39.clk1_input_clock_enable = "ena3";
defparam ram_block1a39.clk1_output_clock_enable = "ena1";
defparam ram_block1a39.clock_duty_cycle_dependence = "on";
defparam ram_block1a39.data_interleave_offset_in_bits = 1;
defparam ram_block1a39.data_interleave_width_in_bits = 1;
defparam ram_block1a39.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a39.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a39.operation_mode = "dual_port";
defparam ram_block1a39.port_a_address_clear = "none";
defparam ram_block1a39.port_a_address_width = 8;
defparam ram_block1a39.port_a_data_out_clear = "none";
defparam ram_block1a39.port_a_data_out_clock = "none";
defparam ram_block1a39.port_a_data_width = 1;
defparam ram_block1a39.port_a_first_address = 0;
defparam ram_block1a39.port_a_first_bit_number = 39;
defparam ram_block1a39.port_a_last_address = 255;
defparam ram_block1a39.port_a_logical_ram_depth = 256;
defparam ram_block1a39.port_a_logical_ram_width = 144;
defparam ram_block1a39.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a39.port_b_address_clear = "none";
defparam ram_block1a39.port_b_address_clock = "clock1";
defparam ram_block1a39.port_b_address_width = 8;
defparam ram_block1a39.port_b_data_out_clear = "none";
defparam ram_block1a39.port_b_data_out_clock = "clock1";
defparam ram_block1a39.port_b_data_width = 1;
defparam ram_block1a39.port_b_first_address = 0;
defparam ram_block1a39.port_b_first_bit_number = 39;
defparam ram_block1a39.port_b_last_address = 255;
defparam ram_block1a39.port_b_logical_ram_depth = 256;
defparam ram_block1a39.port_b_logical_ram_width = 144;
defparam ram_block1a39.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a39.port_b_read_enable_clock = "clock1";
defparam ram_block1a39.ram_block_type = "auto";

arriaii_ram_block ram_block1a71(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[71]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a71_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a71.clk0_core_clock_enable = "ena0";
defparam ram_block1a71.clk0_input_clock_enable = "ena2";
defparam ram_block1a71.clk1_core_clock_enable = "ena3";
defparam ram_block1a71.clk1_input_clock_enable = "ena3";
defparam ram_block1a71.clk1_output_clock_enable = "ena1";
defparam ram_block1a71.clock_duty_cycle_dependence = "on";
defparam ram_block1a71.data_interleave_offset_in_bits = 1;
defparam ram_block1a71.data_interleave_width_in_bits = 1;
defparam ram_block1a71.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a71.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a71.operation_mode = "dual_port";
defparam ram_block1a71.port_a_address_clear = "none";
defparam ram_block1a71.port_a_address_width = 8;
defparam ram_block1a71.port_a_data_out_clear = "none";
defparam ram_block1a71.port_a_data_out_clock = "none";
defparam ram_block1a71.port_a_data_width = 1;
defparam ram_block1a71.port_a_first_address = 0;
defparam ram_block1a71.port_a_first_bit_number = 71;
defparam ram_block1a71.port_a_last_address = 255;
defparam ram_block1a71.port_a_logical_ram_depth = 256;
defparam ram_block1a71.port_a_logical_ram_width = 144;
defparam ram_block1a71.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a71.port_b_address_clear = "none";
defparam ram_block1a71.port_b_address_clock = "clock1";
defparam ram_block1a71.port_b_address_width = 8;
defparam ram_block1a71.port_b_data_out_clear = "none";
defparam ram_block1a71.port_b_data_out_clock = "clock1";
defparam ram_block1a71.port_b_data_width = 1;
defparam ram_block1a71.port_b_first_address = 0;
defparam ram_block1a71.port_b_first_bit_number = 71;
defparam ram_block1a71.port_b_last_address = 255;
defparam ram_block1a71.port_b_logical_ram_depth = 256;
defparam ram_block1a71.port_b_logical_ram_width = 144;
defparam ram_block1a71.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a71.port_b_read_enable_clock = "clock1";
defparam ram_block1a71.ram_block_type = "auto";

arriaii_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena2";
defparam ram_block1a7.clk1_core_clock_enable = "ena3";
defparam ram_block1a7.clk1_input_clock_enable = "ena3";
defparam ram_block1a7.clk1_output_clock_enable = "ena1";
defparam ram_block1a7.clock_duty_cycle_dependence = "on";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 8;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 255;
defparam ram_block1a7.port_a_logical_ram_depth = 256;
defparam ram_block1a7.port_a_logical_ram_width = 144;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 8;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 255;
defparam ram_block1a7.port_b_logical_ram_depth = 256;
defparam ram_block1a7.port_b_logical_ram_width = 144;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

arriaii_ram_block ram_block1a104(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[104]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a104_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a104.clk0_core_clock_enable = "ena0";
defparam ram_block1a104.clk0_input_clock_enable = "ena2";
defparam ram_block1a104.clk1_core_clock_enable = "ena3";
defparam ram_block1a104.clk1_input_clock_enable = "ena3";
defparam ram_block1a104.clk1_output_clock_enable = "ena1";
defparam ram_block1a104.clock_duty_cycle_dependence = "on";
defparam ram_block1a104.data_interleave_offset_in_bits = 1;
defparam ram_block1a104.data_interleave_width_in_bits = 1;
defparam ram_block1a104.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a104.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a104.operation_mode = "dual_port";
defparam ram_block1a104.port_a_address_clear = "none";
defparam ram_block1a104.port_a_address_width = 8;
defparam ram_block1a104.port_a_data_out_clear = "none";
defparam ram_block1a104.port_a_data_out_clock = "none";
defparam ram_block1a104.port_a_data_width = 1;
defparam ram_block1a104.port_a_first_address = 0;
defparam ram_block1a104.port_a_first_bit_number = 104;
defparam ram_block1a104.port_a_last_address = 255;
defparam ram_block1a104.port_a_logical_ram_depth = 256;
defparam ram_block1a104.port_a_logical_ram_width = 144;
defparam ram_block1a104.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a104.port_b_address_clear = "none";
defparam ram_block1a104.port_b_address_clock = "clock1";
defparam ram_block1a104.port_b_address_width = 8;
defparam ram_block1a104.port_b_data_out_clear = "none";
defparam ram_block1a104.port_b_data_out_clock = "clock1";
defparam ram_block1a104.port_b_data_width = 1;
defparam ram_block1a104.port_b_first_address = 0;
defparam ram_block1a104.port_b_first_bit_number = 104;
defparam ram_block1a104.port_b_last_address = 255;
defparam ram_block1a104.port_b_logical_ram_depth = 256;
defparam ram_block1a104.port_b_logical_ram_width = 144;
defparam ram_block1a104.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a104.port_b_read_enable_clock = "clock1";
defparam ram_block1a104.ram_block_type = "auto";

arriaii_ram_block ram_block1a40(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[40]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a40_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a40.clk0_core_clock_enable = "ena0";
defparam ram_block1a40.clk0_input_clock_enable = "ena2";
defparam ram_block1a40.clk1_core_clock_enable = "ena3";
defparam ram_block1a40.clk1_input_clock_enable = "ena3";
defparam ram_block1a40.clk1_output_clock_enable = "ena1";
defparam ram_block1a40.clock_duty_cycle_dependence = "on";
defparam ram_block1a40.data_interleave_offset_in_bits = 1;
defparam ram_block1a40.data_interleave_width_in_bits = 1;
defparam ram_block1a40.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a40.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a40.operation_mode = "dual_port";
defparam ram_block1a40.port_a_address_clear = "none";
defparam ram_block1a40.port_a_address_width = 8;
defparam ram_block1a40.port_a_data_out_clear = "none";
defparam ram_block1a40.port_a_data_out_clock = "none";
defparam ram_block1a40.port_a_data_width = 1;
defparam ram_block1a40.port_a_first_address = 0;
defparam ram_block1a40.port_a_first_bit_number = 40;
defparam ram_block1a40.port_a_last_address = 255;
defparam ram_block1a40.port_a_logical_ram_depth = 256;
defparam ram_block1a40.port_a_logical_ram_width = 144;
defparam ram_block1a40.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a40.port_b_address_clear = "none";
defparam ram_block1a40.port_b_address_clock = "clock1";
defparam ram_block1a40.port_b_address_width = 8;
defparam ram_block1a40.port_b_data_out_clear = "none";
defparam ram_block1a40.port_b_data_out_clock = "clock1";
defparam ram_block1a40.port_b_data_width = 1;
defparam ram_block1a40.port_b_first_address = 0;
defparam ram_block1a40.port_b_first_bit_number = 40;
defparam ram_block1a40.port_b_last_address = 255;
defparam ram_block1a40.port_b_logical_ram_depth = 256;
defparam ram_block1a40.port_b_logical_ram_width = 144;
defparam ram_block1a40.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a40.port_b_read_enable_clock = "clock1";
defparam ram_block1a40.ram_block_type = "auto";

arriaii_ram_block ram_block1a72(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[72]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a72_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a72.clk0_core_clock_enable = "ena0";
defparam ram_block1a72.clk0_input_clock_enable = "ena2";
defparam ram_block1a72.clk1_core_clock_enable = "ena3";
defparam ram_block1a72.clk1_input_clock_enable = "ena3";
defparam ram_block1a72.clk1_output_clock_enable = "ena1";
defparam ram_block1a72.clock_duty_cycle_dependence = "on";
defparam ram_block1a72.data_interleave_offset_in_bits = 1;
defparam ram_block1a72.data_interleave_width_in_bits = 1;
defparam ram_block1a72.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a72.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a72.operation_mode = "dual_port";
defparam ram_block1a72.port_a_address_clear = "none";
defparam ram_block1a72.port_a_address_width = 8;
defparam ram_block1a72.port_a_data_out_clear = "none";
defparam ram_block1a72.port_a_data_out_clock = "none";
defparam ram_block1a72.port_a_data_width = 1;
defparam ram_block1a72.port_a_first_address = 0;
defparam ram_block1a72.port_a_first_bit_number = 72;
defparam ram_block1a72.port_a_last_address = 255;
defparam ram_block1a72.port_a_logical_ram_depth = 256;
defparam ram_block1a72.port_a_logical_ram_width = 144;
defparam ram_block1a72.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a72.port_b_address_clear = "none";
defparam ram_block1a72.port_b_address_clock = "clock1";
defparam ram_block1a72.port_b_address_width = 8;
defparam ram_block1a72.port_b_data_out_clear = "none";
defparam ram_block1a72.port_b_data_out_clock = "clock1";
defparam ram_block1a72.port_b_data_width = 1;
defparam ram_block1a72.port_b_first_address = 0;
defparam ram_block1a72.port_b_first_bit_number = 72;
defparam ram_block1a72.port_b_last_address = 255;
defparam ram_block1a72.port_b_logical_ram_depth = 256;
defparam ram_block1a72.port_b_logical_ram_width = 144;
defparam ram_block1a72.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a72.port_b_read_enable_clock = "clock1";
defparam ram_block1a72.ram_block_type = "auto";

arriaii_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena2";
defparam ram_block1a8.clk1_core_clock_enable = "ena3";
defparam ram_block1a8.clk1_input_clock_enable = "ena3";
defparam ram_block1a8.clk1_output_clock_enable = "ena1";
defparam ram_block1a8.clock_duty_cycle_dependence = "on";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 8;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 255;
defparam ram_block1a8.port_a_logical_ram_depth = 256;
defparam ram_block1a8.port_a_logical_ram_width = 144;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 8;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 255;
defparam ram_block1a8.port_b_logical_ram_depth = 256;
defparam ram_block1a8.port_b_logical_ram_width = 144;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

arriaii_ram_block ram_block1a105(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[105]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a105_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a105.clk0_core_clock_enable = "ena0";
defparam ram_block1a105.clk0_input_clock_enable = "ena2";
defparam ram_block1a105.clk1_core_clock_enable = "ena3";
defparam ram_block1a105.clk1_input_clock_enable = "ena3";
defparam ram_block1a105.clk1_output_clock_enable = "ena1";
defparam ram_block1a105.clock_duty_cycle_dependence = "on";
defparam ram_block1a105.data_interleave_offset_in_bits = 1;
defparam ram_block1a105.data_interleave_width_in_bits = 1;
defparam ram_block1a105.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a105.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a105.operation_mode = "dual_port";
defparam ram_block1a105.port_a_address_clear = "none";
defparam ram_block1a105.port_a_address_width = 8;
defparam ram_block1a105.port_a_data_out_clear = "none";
defparam ram_block1a105.port_a_data_out_clock = "none";
defparam ram_block1a105.port_a_data_width = 1;
defparam ram_block1a105.port_a_first_address = 0;
defparam ram_block1a105.port_a_first_bit_number = 105;
defparam ram_block1a105.port_a_last_address = 255;
defparam ram_block1a105.port_a_logical_ram_depth = 256;
defparam ram_block1a105.port_a_logical_ram_width = 144;
defparam ram_block1a105.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a105.port_b_address_clear = "none";
defparam ram_block1a105.port_b_address_clock = "clock1";
defparam ram_block1a105.port_b_address_width = 8;
defparam ram_block1a105.port_b_data_out_clear = "none";
defparam ram_block1a105.port_b_data_out_clock = "clock1";
defparam ram_block1a105.port_b_data_width = 1;
defparam ram_block1a105.port_b_first_address = 0;
defparam ram_block1a105.port_b_first_bit_number = 105;
defparam ram_block1a105.port_b_last_address = 255;
defparam ram_block1a105.port_b_logical_ram_depth = 256;
defparam ram_block1a105.port_b_logical_ram_width = 144;
defparam ram_block1a105.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a105.port_b_read_enable_clock = "clock1";
defparam ram_block1a105.ram_block_type = "auto";

arriaii_ram_block ram_block1a41(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[41]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a41_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a41.clk0_core_clock_enable = "ena0";
defparam ram_block1a41.clk0_input_clock_enable = "ena2";
defparam ram_block1a41.clk1_core_clock_enable = "ena3";
defparam ram_block1a41.clk1_input_clock_enable = "ena3";
defparam ram_block1a41.clk1_output_clock_enable = "ena1";
defparam ram_block1a41.clock_duty_cycle_dependence = "on";
defparam ram_block1a41.data_interleave_offset_in_bits = 1;
defparam ram_block1a41.data_interleave_width_in_bits = 1;
defparam ram_block1a41.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a41.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a41.operation_mode = "dual_port";
defparam ram_block1a41.port_a_address_clear = "none";
defparam ram_block1a41.port_a_address_width = 8;
defparam ram_block1a41.port_a_data_out_clear = "none";
defparam ram_block1a41.port_a_data_out_clock = "none";
defparam ram_block1a41.port_a_data_width = 1;
defparam ram_block1a41.port_a_first_address = 0;
defparam ram_block1a41.port_a_first_bit_number = 41;
defparam ram_block1a41.port_a_last_address = 255;
defparam ram_block1a41.port_a_logical_ram_depth = 256;
defparam ram_block1a41.port_a_logical_ram_width = 144;
defparam ram_block1a41.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a41.port_b_address_clear = "none";
defparam ram_block1a41.port_b_address_clock = "clock1";
defparam ram_block1a41.port_b_address_width = 8;
defparam ram_block1a41.port_b_data_out_clear = "none";
defparam ram_block1a41.port_b_data_out_clock = "clock1";
defparam ram_block1a41.port_b_data_width = 1;
defparam ram_block1a41.port_b_first_address = 0;
defparam ram_block1a41.port_b_first_bit_number = 41;
defparam ram_block1a41.port_b_last_address = 255;
defparam ram_block1a41.port_b_logical_ram_depth = 256;
defparam ram_block1a41.port_b_logical_ram_width = 144;
defparam ram_block1a41.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a41.port_b_read_enable_clock = "clock1";
defparam ram_block1a41.ram_block_type = "auto";

arriaii_ram_block ram_block1a73(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[73]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a73_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a73.clk0_core_clock_enable = "ena0";
defparam ram_block1a73.clk0_input_clock_enable = "ena2";
defparam ram_block1a73.clk1_core_clock_enable = "ena3";
defparam ram_block1a73.clk1_input_clock_enable = "ena3";
defparam ram_block1a73.clk1_output_clock_enable = "ena1";
defparam ram_block1a73.clock_duty_cycle_dependence = "on";
defparam ram_block1a73.data_interleave_offset_in_bits = 1;
defparam ram_block1a73.data_interleave_width_in_bits = 1;
defparam ram_block1a73.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a73.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a73.operation_mode = "dual_port";
defparam ram_block1a73.port_a_address_clear = "none";
defparam ram_block1a73.port_a_address_width = 8;
defparam ram_block1a73.port_a_data_out_clear = "none";
defparam ram_block1a73.port_a_data_out_clock = "none";
defparam ram_block1a73.port_a_data_width = 1;
defparam ram_block1a73.port_a_first_address = 0;
defparam ram_block1a73.port_a_first_bit_number = 73;
defparam ram_block1a73.port_a_last_address = 255;
defparam ram_block1a73.port_a_logical_ram_depth = 256;
defparam ram_block1a73.port_a_logical_ram_width = 144;
defparam ram_block1a73.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a73.port_b_address_clear = "none";
defparam ram_block1a73.port_b_address_clock = "clock1";
defparam ram_block1a73.port_b_address_width = 8;
defparam ram_block1a73.port_b_data_out_clear = "none";
defparam ram_block1a73.port_b_data_out_clock = "clock1";
defparam ram_block1a73.port_b_data_width = 1;
defparam ram_block1a73.port_b_first_address = 0;
defparam ram_block1a73.port_b_first_bit_number = 73;
defparam ram_block1a73.port_b_last_address = 255;
defparam ram_block1a73.port_b_logical_ram_depth = 256;
defparam ram_block1a73.port_b_logical_ram_width = 144;
defparam ram_block1a73.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a73.port_b_read_enable_clock = "clock1";
defparam ram_block1a73.ram_block_type = "auto";

arriaii_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena2";
defparam ram_block1a9.clk1_core_clock_enable = "ena3";
defparam ram_block1a9.clk1_input_clock_enable = "ena3";
defparam ram_block1a9.clk1_output_clock_enable = "ena1";
defparam ram_block1a9.clock_duty_cycle_dependence = "on";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 8;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 255;
defparam ram_block1a9.port_a_logical_ram_depth = 256;
defparam ram_block1a9.port_a_logical_ram_width = 144;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 8;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 255;
defparam ram_block1a9.port_b_logical_ram_depth = 256;
defparam ram_block1a9.port_b_logical_ram_width = 144;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

arriaii_ram_block ram_block1a106(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[106]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a106_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a106.clk0_core_clock_enable = "ena0";
defparam ram_block1a106.clk0_input_clock_enable = "ena2";
defparam ram_block1a106.clk1_core_clock_enable = "ena3";
defparam ram_block1a106.clk1_input_clock_enable = "ena3";
defparam ram_block1a106.clk1_output_clock_enable = "ena1";
defparam ram_block1a106.clock_duty_cycle_dependence = "on";
defparam ram_block1a106.data_interleave_offset_in_bits = 1;
defparam ram_block1a106.data_interleave_width_in_bits = 1;
defparam ram_block1a106.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a106.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a106.operation_mode = "dual_port";
defparam ram_block1a106.port_a_address_clear = "none";
defparam ram_block1a106.port_a_address_width = 8;
defparam ram_block1a106.port_a_data_out_clear = "none";
defparam ram_block1a106.port_a_data_out_clock = "none";
defparam ram_block1a106.port_a_data_width = 1;
defparam ram_block1a106.port_a_first_address = 0;
defparam ram_block1a106.port_a_first_bit_number = 106;
defparam ram_block1a106.port_a_last_address = 255;
defparam ram_block1a106.port_a_logical_ram_depth = 256;
defparam ram_block1a106.port_a_logical_ram_width = 144;
defparam ram_block1a106.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a106.port_b_address_clear = "none";
defparam ram_block1a106.port_b_address_clock = "clock1";
defparam ram_block1a106.port_b_address_width = 8;
defparam ram_block1a106.port_b_data_out_clear = "none";
defparam ram_block1a106.port_b_data_out_clock = "clock1";
defparam ram_block1a106.port_b_data_width = 1;
defparam ram_block1a106.port_b_first_address = 0;
defparam ram_block1a106.port_b_first_bit_number = 106;
defparam ram_block1a106.port_b_last_address = 255;
defparam ram_block1a106.port_b_logical_ram_depth = 256;
defparam ram_block1a106.port_b_logical_ram_width = 144;
defparam ram_block1a106.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a106.port_b_read_enable_clock = "clock1";
defparam ram_block1a106.ram_block_type = "auto";

arriaii_ram_block ram_block1a42(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[42]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a42_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a42.clk0_core_clock_enable = "ena0";
defparam ram_block1a42.clk0_input_clock_enable = "ena2";
defparam ram_block1a42.clk1_core_clock_enable = "ena3";
defparam ram_block1a42.clk1_input_clock_enable = "ena3";
defparam ram_block1a42.clk1_output_clock_enable = "ena1";
defparam ram_block1a42.clock_duty_cycle_dependence = "on";
defparam ram_block1a42.data_interleave_offset_in_bits = 1;
defparam ram_block1a42.data_interleave_width_in_bits = 1;
defparam ram_block1a42.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a42.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a42.operation_mode = "dual_port";
defparam ram_block1a42.port_a_address_clear = "none";
defparam ram_block1a42.port_a_address_width = 8;
defparam ram_block1a42.port_a_data_out_clear = "none";
defparam ram_block1a42.port_a_data_out_clock = "none";
defparam ram_block1a42.port_a_data_width = 1;
defparam ram_block1a42.port_a_first_address = 0;
defparam ram_block1a42.port_a_first_bit_number = 42;
defparam ram_block1a42.port_a_last_address = 255;
defparam ram_block1a42.port_a_logical_ram_depth = 256;
defparam ram_block1a42.port_a_logical_ram_width = 144;
defparam ram_block1a42.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a42.port_b_address_clear = "none";
defparam ram_block1a42.port_b_address_clock = "clock1";
defparam ram_block1a42.port_b_address_width = 8;
defparam ram_block1a42.port_b_data_out_clear = "none";
defparam ram_block1a42.port_b_data_out_clock = "clock1";
defparam ram_block1a42.port_b_data_width = 1;
defparam ram_block1a42.port_b_first_address = 0;
defparam ram_block1a42.port_b_first_bit_number = 42;
defparam ram_block1a42.port_b_last_address = 255;
defparam ram_block1a42.port_b_logical_ram_depth = 256;
defparam ram_block1a42.port_b_logical_ram_width = 144;
defparam ram_block1a42.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a42.port_b_read_enable_clock = "clock1";
defparam ram_block1a42.ram_block_type = "auto";

arriaii_ram_block ram_block1a74(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[74]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a74_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a74.clk0_core_clock_enable = "ena0";
defparam ram_block1a74.clk0_input_clock_enable = "ena2";
defparam ram_block1a74.clk1_core_clock_enable = "ena3";
defparam ram_block1a74.clk1_input_clock_enable = "ena3";
defparam ram_block1a74.clk1_output_clock_enable = "ena1";
defparam ram_block1a74.clock_duty_cycle_dependence = "on";
defparam ram_block1a74.data_interleave_offset_in_bits = 1;
defparam ram_block1a74.data_interleave_width_in_bits = 1;
defparam ram_block1a74.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a74.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a74.operation_mode = "dual_port";
defparam ram_block1a74.port_a_address_clear = "none";
defparam ram_block1a74.port_a_address_width = 8;
defparam ram_block1a74.port_a_data_out_clear = "none";
defparam ram_block1a74.port_a_data_out_clock = "none";
defparam ram_block1a74.port_a_data_width = 1;
defparam ram_block1a74.port_a_first_address = 0;
defparam ram_block1a74.port_a_first_bit_number = 74;
defparam ram_block1a74.port_a_last_address = 255;
defparam ram_block1a74.port_a_logical_ram_depth = 256;
defparam ram_block1a74.port_a_logical_ram_width = 144;
defparam ram_block1a74.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a74.port_b_address_clear = "none";
defparam ram_block1a74.port_b_address_clock = "clock1";
defparam ram_block1a74.port_b_address_width = 8;
defparam ram_block1a74.port_b_data_out_clear = "none";
defparam ram_block1a74.port_b_data_out_clock = "clock1";
defparam ram_block1a74.port_b_data_width = 1;
defparam ram_block1a74.port_b_first_address = 0;
defparam ram_block1a74.port_b_first_bit_number = 74;
defparam ram_block1a74.port_b_last_address = 255;
defparam ram_block1a74.port_b_logical_ram_depth = 256;
defparam ram_block1a74.port_b_logical_ram_width = 144;
defparam ram_block1a74.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a74.port_b_read_enable_clock = "clock1";
defparam ram_block1a74.ram_block_type = "auto";

arriaii_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena2";
defparam ram_block1a10.clk1_core_clock_enable = "ena3";
defparam ram_block1a10.clk1_input_clock_enable = "ena3";
defparam ram_block1a10.clk1_output_clock_enable = "ena1";
defparam ram_block1a10.clock_duty_cycle_dependence = "on";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 8;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 255;
defparam ram_block1a10.port_a_logical_ram_depth = 256;
defparam ram_block1a10.port_a_logical_ram_width = 144;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 8;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 255;
defparam ram_block1a10.port_b_logical_ram_depth = 256;
defparam ram_block1a10.port_b_logical_ram_width = 144;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

arriaii_ram_block ram_block1a107(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[107]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a107_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a107.clk0_core_clock_enable = "ena0";
defparam ram_block1a107.clk0_input_clock_enable = "ena2";
defparam ram_block1a107.clk1_core_clock_enable = "ena3";
defparam ram_block1a107.clk1_input_clock_enable = "ena3";
defparam ram_block1a107.clk1_output_clock_enable = "ena1";
defparam ram_block1a107.clock_duty_cycle_dependence = "on";
defparam ram_block1a107.data_interleave_offset_in_bits = 1;
defparam ram_block1a107.data_interleave_width_in_bits = 1;
defparam ram_block1a107.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a107.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a107.operation_mode = "dual_port";
defparam ram_block1a107.port_a_address_clear = "none";
defparam ram_block1a107.port_a_address_width = 8;
defparam ram_block1a107.port_a_data_out_clear = "none";
defparam ram_block1a107.port_a_data_out_clock = "none";
defparam ram_block1a107.port_a_data_width = 1;
defparam ram_block1a107.port_a_first_address = 0;
defparam ram_block1a107.port_a_first_bit_number = 107;
defparam ram_block1a107.port_a_last_address = 255;
defparam ram_block1a107.port_a_logical_ram_depth = 256;
defparam ram_block1a107.port_a_logical_ram_width = 144;
defparam ram_block1a107.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a107.port_b_address_clear = "none";
defparam ram_block1a107.port_b_address_clock = "clock1";
defparam ram_block1a107.port_b_address_width = 8;
defparam ram_block1a107.port_b_data_out_clear = "none";
defparam ram_block1a107.port_b_data_out_clock = "clock1";
defparam ram_block1a107.port_b_data_width = 1;
defparam ram_block1a107.port_b_first_address = 0;
defparam ram_block1a107.port_b_first_bit_number = 107;
defparam ram_block1a107.port_b_last_address = 255;
defparam ram_block1a107.port_b_logical_ram_depth = 256;
defparam ram_block1a107.port_b_logical_ram_width = 144;
defparam ram_block1a107.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a107.port_b_read_enable_clock = "clock1";
defparam ram_block1a107.ram_block_type = "auto";

arriaii_ram_block ram_block1a43(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[43]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a43_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a43.clk0_core_clock_enable = "ena0";
defparam ram_block1a43.clk0_input_clock_enable = "ena2";
defparam ram_block1a43.clk1_core_clock_enable = "ena3";
defparam ram_block1a43.clk1_input_clock_enable = "ena3";
defparam ram_block1a43.clk1_output_clock_enable = "ena1";
defparam ram_block1a43.clock_duty_cycle_dependence = "on";
defparam ram_block1a43.data_interleave_offset_in_bits = 1;
defparam ram_block1a43.data_interleave_width_in_bits = 1;
defparam ram_block1a43.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a43.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a43.operation_mode = "dual_port";
defparam ram_block1a43.port_a_address_clear = "none";
defparam ram_block1a43.port_a_address_width = 8;
defparam ram_block1a43.port_a_data_out_clear = "none";
defparam ram_block1a43.port_a_data_out_clock = "none";
defparam ram_block1a43.port_a_data_width = 1;
defparam ram_block1a43.port_a_first_address = 0;
defparam ram_block1a43.port_a_first_bit_number = 43;
defparam ram_block1a43.port_a_last_address = 255;
defparam ram_block1a43.port_a_logical_ram_depth = 256;
defparam ram_block1a43.port_a_logical_ram_width = 144;
defparam ram_block1a43.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a43.port_b_address_clear = "none";
defparam ram_block1a43.port_b_address_clock = "clock1";
defparam ram_block1a43.port_b_address_width = 8;
defparam ram_block1a43.port_b_data_out_clear = "none";
defparam ram_block1a43.port_b_data_out_clock = "clock1";
defparam ram_block1a43.port_b_data_width = 1;
defparam ram_block1a43.port_b_first_address = 0;
defparam ram_block1a43.port_b_first_bit_number = 43;
defparam ram_block1a43.port_b_last_address = 255;
defparam ram_block1a43.port_b_logical_ram_depth = 256;
defparam ram_block1a43.port_b_logical_ram_width = 144;
defparam ram_block1a43.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a43.port_b_read_enable_clock = "clock1";
defparam ram_block1a43.ram_block_type = "auto";

arriaii_ram_block ram_block1a75(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[75]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a75_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a75.clk0_core_clock_enable = "ena0";
defparam ram_block1a75.clk0_input_clock_enable = "ena2";
defparam ram_block1a75.clk1_core_clock_enable = "ena3";
defparam ram_block1a75.clk1_input_clock_enable = "ena3";
defparam ram_block1a75.clk1_output_clock_enable = "ena1";
defparam ram_block1a75.clock_duty_cycle_dependence = "on";
defparam ram_block1a75.data_interleave_offset_in_bits = 1;
defparam ram_block1a75.data_interleave_width_in_bits = 1;
defparam ram_block1a75.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a75.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a75.operation_mode = "dual_port";
defparam ram_block1a75.port_a_address_clear = "none";
defparam ram_block1a75.port_a_address_width = 8;
defparam ram_block1a75.port_a_data_out_clear = "none";
defparam ram_block1a75.port_a_data_out_clock = "none";
defparam ram_block1a75.port_a_data_width = 1;
defparam ram_block1a75.port_a_first_address = 0;
defparam ram_block1a75.port_a_first_bit_number = 75;
defparam ram_block1a75.port_a_last_address = 255;
defparam ram_block1a75.port_a_logical_ram_depth = 256;
defparam ram_block1a75.port_a_logical_ram_width = 144;
defparam ram_block1a75.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a75.port_b_address_clear = "none";
defparam ram_block1a75.port_b_address_clock = "clock1";
defparam ram_block1a75.port_b_address_width = 8;
defparam ram_block1a75.port_b_data_out_clear = "none";
defparam ram_block1a75.port_b_data_out_clock = "clock1";
defparam ram_block1a75.port_b_data_width = 1;
defparam ram_block1a75.port_b_first_address = 0;
defparam ram_block1a75.port_b_first_bit_number = 75;
defparam ram_block1a75.port_b_last_address = 255;
defparam ram_block1a75.port_b_logical_ram_depth = 256;
defparam ram_block1a75.port_b_logical_ram_width = 144;
defparam ram_block1a75.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a75.port_b_read_enable_clock = "clock1";
defparam ram_block1a75.ram_block_type = "auto";

arriaii_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena2";
defparam ram_block1a11.clk1_core_clock_enable = "ena3";
defparam ram_block1a11.clk1_input_clock_enable = "ena3";
defparam ram_block1a11.clk1_output_clock_enable = "ena1";
defparam ram_block1a11.clock_duty_cycle_dependence = "on";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 8;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 255;
defparam ram_block1a11.port_a_logical_ram_depth = 256;
defparam ram_block1a11.port_a_logical_ram_width = 144;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 8;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 255;
defparam ram_block1a11.port_b_logical_ram_depth = 256;
defparam ram_block1a11.port_b_logical_ram_width = 144;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

arriaii_ram_block ram_block1a108(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[108]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a108_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a108.clk0_core_clock_enable = "ena0";
defparam ram_block1a108.clk0_input_clock_enable = "ena2";
defparam ram_block1a108.clk1_core_clock_enable = "ena3";
defparam ram_block1a108.clk1_input_clock_enable = "ena3";
defparam ram_block1a108.clk1_output_clock_enable = "ena1";
defparam ram_block1a108.clock_duty_cycle_dependence = "on";
defparam ram_block1a108.data_interleave_offset_in_bits = 1;
defparam ram_block1a108.data_interleave_width_in_bits = 1;
defparam ram_block1a108.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a108.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a108.operation_mode = "dual_port";
defparam ram_block1a108.port_a_address_clear = "none";
defparam ram_block1a108.port_a_address_width = 8;
defparam ram_block1a108.port_a_data_out_clear = "none";
defparam ram_block1a108.port_a_data_out_clock = "none";
defparam ram_block1a108.port_a_data_width = 1;
defparam ram_block1a108.port_a_first_address = 0;
defparam ram_block1a108.port_a_first_bit_number = 108;
defparam ram_block1a108.port_a_last_address = 255;
defparam ram_block1a108.port_a_logical_ram_depth = 256;
defparam ram_block1a108.port_a_logical_ram_width = 144;
defparam ram_block1a108.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a108.port_b_address_clear = "none";
defparam ram_block1a108.port_b_address_clock = "clock1";
defparam ram_block1a108.port_b_address_width = 8;
defparam ram_block1a108.port_b_data_out_clear = "none";
defparam ram_block1a108.port_b_data_out_clock = "clock1";
defparam ram_block1a108.port_b_data_width = 1;
defparam ram_block1a108.port_b_first_address = 0;
defparam ram_block1a108.port_b_first_bit_number = 108;
defparam ram_block1a108.port_b_last_address = 255;
defparam ram_block1a108.port_b_logical_ram_depth = 256;
defparam ram_block1a108.port_b_logical_ram_width = 144;
defparam ram_block1a108.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a108.port_b_read_enable_clock = "clock1";
defparam ram_block1a108.ram_block_type = "auto";

arriaii_ram_block ram_block1a44(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[44]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a44_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a44.clk0_core_clock_enable = "ena0";
defparam ram_block1a44.clk0_input_clock_enable = "ena2";
defparam ram_block1a44.clk1_core_clock_enable = "ena3";
defparam ram_block1a44.clk1_input_clock_enable = "ena3";
defparam ram_block1a44.clk1_output_clock_enable = "ena1";
defparam ram_block1a44.clock_duty_cycle_dependence = "on";
defparam ram_block1a44.data_interleave_offset_in_bits = 1;
defparam ram_block1a44.data_interleave_width_in_bits = 1;
defparam ram_block1a44.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a44.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a44.operation_mode = "dual_port";
defparam ram_block1a44.port_a_address_clear = "none";
defparam ram_block1a44.port_a_address_width = 8;
defparam ram_block1a44.port_a_data_out_clear = "none";
defparam ram_block1a44.port_a_data_out_clock = "none";
defparam ram_block1a44.port_a_data_width = 1;
defparam ram_block1a44.port_a_first_address = 0;
defparam ram_block1a44.port_a_first_bit_number = 44;
defparam ram_block1a44.port_a_last_address = 255;
defparam ram_block1a44.port_a_logical_ram_depth = 256;
defparam ram_block1a44.port_a_logical_ram_width = 144;
defparam ram_block1a44.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a44.port_b_address_clear = "none";
defparam ram_block1a44.port_b_address_clock = "clock1";
defparam ram_block1a44.port_b_address_width = 8;
defparam ram_block1a44.port_b_data_out_clear = "none";
defparam ram_block1a44.port_b_data_out_clock = "clock1";
defparam ram_block1a44.port_b_data_width = 1;
defparam ram_block1a44.port_b_first_address = 0;
defparam ram_block1a44.port_b_first_bit_number = 44;
defparam ram_block1a44.port_b_last_address = 255;
defparam ram_block1a44.port_b_logical_ram_depth = 256;
defparam ram_block1a44.port_b_logical_ram_width = 144;
defparam ram_block1a44.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a44.port_b_read_enable_clock = "clock1";
defparam ram_block1a44.ram_block_type = "auto";

arriaii_ram_block ram_block1a76(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[76]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a76_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a76.clk0_core_clock_enable = "ena0";
defparam ram_block1a76.clk0_input_clock_enable = "ena2";
defparam ram_block1a76.clk1_core_clock_enable = "ena3";
defparam ram_block1a76.clk1_input_clock_enable = "ena3";
defparam ram_block1a76.clk1_output_clock_enable = "ena1";
defparam ram_block1a76.clock_duty_cycle_dependence = "on";
defparam ram_block1a76.data_interleave_offset_in_bits = 1;
defparam ram_block1a76.data_interleave_width_in_bits = 1;
defparam ram_block1a76.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a76.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a76.operation_mode = "dual_port";
defparam ram_block1a76.port_a_address_clear = "none";
defparam ram_block1a76.port_a_address_width = 8;
defparam ram_block1a76.port_a_data_out_clear = "none";
defparam ram_block1a76.port_a_data_out_clock = "none";
defparam ram_block1a76.port_a_data_width = 1;
defparam ram_block1a76.port_a_first_address = 0;
defparam ram_block1a76.port_a_first_bit_number = 76;
defparam ram_block1a76.port_a_last_address = 255;
defparam ram_block1a76.port_a_logical_ram_depth = 256;
defparam ram_block1a76.port_a_logical_ram_width = 144;
defparam ram_block1a76.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a76.port_b_address_clear = "none";
defparam ram_block1a76.port_b_address_clock = "clock1";
defparam ram_block1a76.port_b_address_width = 8;
defparam ram_block1a76.port_b_data_out_clear = "none";
defparam ram_block1a76.port_b_data_out_clock = "clock1";
defparam ram_block1a76.port_b_data_width = 1;
defparam ram_block1a76.port_b_first_address = 0;
defparam ram_block1a76.port_b_first_bit_number = 76;
defparam ram_block1a76.port_b_last_address = 255;
defparam ram_block1a76.port_b_logical_ram_depth = 256;
defparam ram_block1a76.port_b_logical_ram_width = 144;
defparam ram_block1a76.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a76.port_b_read_enable_clock = "clock1";
defparam ram_block1a76.ram_block_type = "auto";

arriaii_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena2";
defparam ram_block1a12.clk1_core_clock_enable = "ena3";
defparam ram_block1a12.clk1_input_clock_enable = "ena3";
defparam ram_block1a12.clk1_output_clock_enable = "ena1";
defparam ram_block1a12.clock_duty_cycle_dependence = "on";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 8;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 255;
defparam ram_block1a12.port_a_logical_ram_depth = 256;
defparam ram_block1a12.port_a_logical_ram_width = 144;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 8;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 255;
defparam ram_block1a12.port_b_logical_ram_depth = 256;
defparam ram_block1a12.port_b_logical_ram_width = 144;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

arriaii_ram_block ram_block1a109(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[109]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a109_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a109.clk0_core_clock_enable = "ena0";
defparam ram_block1a109.clk0_input_clock_enable = "ena2";
defparam ram_block1a109.clk1_core_clock_enable = "ena3";
defparam ram_block1a109.clk1_input_clock_enable = "ena3";
defparam ram_block1a109.clk1_output_clock_enable = "ena1";
defparam ram_block1a109.clock_duty_cycle_dependence = "on";
defparam ram_block1a109.data_interleave_offset_in_bits = 1;
defparam ram_block1a109.data_interleave_width_in_bits = 1;
defparam ram_block1a109.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a109.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a109.operation_mode = "dual_port";
defparam ram_block1a109.port_a_address_clear = "none";
defparam ram_block1a109.port_a_address_width = 8;
defparam ram_block1a109.port_a_data_out_clear = "none";
defparam ram_block1a109.port_a_data_out_clock = "none";
defparam ram_block1a109.port_a_data_width = 1;
defparam ram_block1a109.port_a_first_address = 0;
defparam ram_block1a109.port_a_first_bit_number = 109;
defparam ram_block1a109.port_a_last_address = 255;
defparam ram_block1a109.port_a_logical_ram_depth = 256;
defparam ram_block1a109.port_a_logical_ram_width = 144;
defparam ram_block1a109.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a109.port_b_address_clear = "none";
defparam ram_block1a109.port_b_address_clock = "clock1";
defparam ram_block1a109.port_b_address_width = 8;
defparam ram_block1a109.port_b_data_out_clear = "none";
defparam ram_block1a109.port_b_data_out_clock = "clock1";
defparam ram_block1a109.port_b_data_width = 1;
defparam ram_block1a109.port_b_first_address = 0;
defparam ram_block1a109.port_b_first_bit_number = 109;
defparam ram_block1a109.port_b_last_address = 255;
defparam ram_block1a109.port_b_logical_ram_depth = 256;
defparam ram_block1a109.port_b_logical_ram_width = 144;
defparam ram_block1a109.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a109.port_b_read_enable_clock = "clock1";
defparam ram_block1a109.ram_block_type = "auto";

arriaii_ram_block ram_block1a45(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[45]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a45_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a45.clk0_core_clock_enable = "ena0";
defparam ram_block1a45.clk0_input_clock_enable = "ena2";
defparam ram_block1a45.clk1_core_clock_enable = "ena3";
defparam ram_block1a45.clk1_input_clock_enable = "ena3";
defparam ram_block1a45.clk1_output_clock_enable = "ena1";
defparam ram_block1a45.clock_duty_cycle_dependence = "on";
defparam ram_block1a45.data_interleave_offset_in_bits = 1;
defparam ram_block1a45.data_interleave_width_in_bits = 1;
defparam ram_block1a45.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a45.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a45.operation_mode = "dual_port";
defparam ram_block1a45.port_a_address_clear = "none";
defparam ram_block1a45.port_a_address_width = 8;
defparam ram_block1a45.port_a_data_out_clear = "none";
defparam ram_block1a45.port_a_data_out_clock = "none";
defparam ram_block1a45.port_a_data_width = 1;
defparam ram_block1a45.port_a_first_address = 0;
defparam ram_block1a45.port_a_first_bit_number = 45;
defparam ram_block1a45.port_a_last_address = 255;
defparam ram_block1a45.port_a_logical_ram_depth = 256;
defparam ram_block1a45.port_a_logical_ram_width = 144;
defparam ram_block1a45.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a45.port_b_address_clear = "none";
defparam ram_block1a45.port_b_address_clock = "clock1";
defparam ram_block1a45.port_b_address_width = 8;
defparam ram_block1a45.port_b_data_out_clear = "none";
defparam ram_block1a45.port_b_data_out_clock = "clock1";
defparam ram_block1a45.port_b_data_width = 1;
defparam ram_block1a45.port_b_first_address = 0;
defparam ram_block1a45.port_b_first_bit_number = 45;
defparam ram_block1a45.port_b_last_address = 255;
defparam ram_block1a45.port_b_logical_ram_depth = 256;
defparam ram_block1a45.port_b_logical_ram_width = 144;
defparam ram_block1a45.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a45.port_b_read_enable_clock = "clock1";
defparam ram_block1a45.ram_block_type = "auto";

arriaii_ram_block ram_block1a77(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[77]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a77_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a77.clk0_core_clock_enable = "ena0";
defparam ram_block1a77.clk0_input_clock_enable = "ena2";
defparam ram_block1a77.clk1_core_clock_enable = "ena3";
defparam ram_block1a77.clk1_input_clock_enable = "ena3";
defparam ram_block1a77.clk1_output_clock_enable = "ena1";
defparam ram_block1a77.clock_duty_cycle_dependence = "on";
defparam ram_block1a77.data_interleave_offset_in_bits = 1;
defparam ram_block1a77.data_interleave_width_in_bits = 1;
defparam ram_block1a77.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a77.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a77.operation_mode = "dual_port";
defparam ram_block1a77.port_a_address_clear = "none";
defparam ram_block1a77.port_a_address_width = 8;
defparam ram_block1a77.port_a_data_out_clear = "none";
defparam ram_block1a77.port_a_data_out_clock = "none";
defparam ram_block1a77.port_a_data_width = 1;
defparam ram_block1a77.port_a_first_address = 0;
defparam ram_block1a77.port_a_first_bit_number = 77;
defparam ram_block1a77.port_a_last_address = 255;
defparam ram_block1a77.port_a_logical_ram_depth = 256;
defparam ram_block1a77.port_a_logical_ram_width = 144;
defparam ram_block1a77.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a77.port_b_address_clear = "none";
defparam ram_block1a77.port_b_address_clock = "clock1";
defparam ram_block1a77.port_b_address_width = 8;
defparam ram_block1a77.port_b_data_out_clear = "none";
defparam ram_block1a77.port_b_data_out_clock = "clock1";
defparam ram_block1a77.port_b_data_width = 1;
defparam ram_block1a77.port_b_first_address = 0;
defparam ram_block1a77.port_b_first_bit_number = 77;
defparam ram_block1a77.port_b_last_address = 255;
defparam ram_block1a77.port_b_logical_ram_depth = 256;
defparam ram_block1a77.port_b_logical_ram_width = 144;
defparam ram_block1a77.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a77.port_b_read_enable_clock = "clock1";
defparam ram_block1a77.ram_block_type = "auto";

arriaii_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena2";
defparam ram_block1a13.clk1_core_clock_enable = "ena3";
defparam ram_block1a13.clk1_input_clock_enable = "ena3";
defparam ram_block1a13.clk1_output_clock_enable = "ena1";
defparam ram_block1a13.clock_duty_cycle_dependence = "on";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 8;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 255;
defparam ram_block1a13.port_a_logical_ram_depth = 256;
defparam ram_block1a13.port_a_logical_ram_width = 144;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 8;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 255;
defparam ram_block1a13.port_b_logical_ram_depth = 256;
defparam ram_block1a13.port_b_logical_ram_width = 144;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

arriaii_ram_block ram_block1a110(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[110]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a110_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a110.clk0_core_clock_enable = "ena0";
defparam ram_block1a110.clk0_input_clock_enable = "ena2";
defparam ram_block1a110.clk1_core_clock_enable = "ena3";
defparam ram_block1a110.clk1_input_clock_enable = "ena3";
defparam ram_block1a110.clk1_output_clock_enable = "ena1";
defparam ram_block1a110.clock_duty_cycle_dependence = "on";
defparam ram_block1a110.data_interleave_offset_in_bits = 1;
defparam ram_block1a110.data_interleave_width_in_bits = 1;
defparam ram_block1a110.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a110.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a110.operation_mode = "dual_port";
defparam ram_block1a110.port_a_address_clear = "none";
defparam ram_block1a110.port_a_address_width = 8;
defparam ram_block1a110.port_a_data_out_clear = "none";
defparam ram_block1a110.port_a_data_out_clock = "none";
defparam ram_block1a110.port_a_data_width = 1;
defparam ram_block1a110.port_a_first_address = 0;
defparam ram_block1a110.port_a_first_bit_number = 110;
defparam ram_block1a110.port_a_last_address = 255;
defparam ram_block1a110.port_a_logical_ram_depth = 256;
defparam ram_block1a110.port_a_logical_ram_width = 144;
defparam ram_block1a110.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a110.port_b_address_clear = "none";
defparam ram_block1a110.port_b_address_clock = "clock1";
defparam ram_block1a110.port_b_address_width = 8;
defparam ram_block1a110.port_b_data_out_clear = "none";
defparam ram_block1a110.port_b_data_out_clock = "clock1";
defparam ram_block1a110.port_b_data_width = 1;
defparam ram_block1a110.port_b_first_address = 0;
defparam ram_block1a110.port_b_first_bit_number = 110;
defparam ram_block1a110.port_b_last_address = 255;
defparam ram_block1a110.port_b_logical_ram_depth = 256;
defparam ram_block1a110.port_b_logical_ram_width = 144;
defparam ram_block1a110.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a110.port_b_read_enable_clock = "clock1";
defparam ram_block1a110.ram_block_type = "auto";

arriaii_ram_block ram_block1a46(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[46]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a46_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a46.clk0_core_clock_enable = "ena0";
defparam ram_block1a46.clk0_input_clock_enable = "ena2";
defparam ram_block1a46.clk1_core_clock_enable = "ena3";
defparam ram_block1a46.clk1_input_clock_enable = "ena3";
defparam ram_block1a46.clk1_output_clock_enable = "ena1";
defparam ram_block1a46.clock_duty_cycle_dependence = "on";
defparam ram_block1a46.data_interleave_offset_in_bits = 1;
defparam ram_block1a46.data_interleave_width_in_bits = 1;
defparam ram_block1a46.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a46.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a46.operation_mode = "dual_port";
defparam ram_block1a46.port_a_address_clear = "none";
defparam ram_block1a46.port_a_address_width = 8;
defparam ram_block1a46.port_a_data_out_clear = "none";
defparam ram_block1a46.port_a_data_out_clock = "none";
defparam ram_block1a46.port_a_data_width = 1;
defparam ram_block1a46.port_a_first_address = 0;
defparam ram_block1a46.port_a_first_bit_number = 46;
defparam ram_block1a46.port_a_last_address = 255;
defparam ram_block1a46.port_a_logical_ram_depth = 256;
defparam ram_block1a46.port_a_logical_ram_width = 144;
defparam ram_block1a46.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a46.port_b_address_clear = "none";
defparam ram_block1a46.port_b_address_clock = "clock1";
defparam ram_block1a46.port_b_address_width = 8;
defparam ram_block1a46.port_b_data_out_clear = "none";
defparam ram_block1a46.port_b_data_out_clock = "clock1";
defparam ram_block1a46.port_b_data_width = 1;
defparam ram_block1a46.port_b_first_address = 0;
defparam ram_block1a46.port_b_first_bit_number = 46;
defparam ram_block1a46.port_b_last_address = 255;
defparam ram_block1a46.port_b_logical_ram_depth = 256;
defparam ram_block1a46.port_b_logical_ram_width = 144;
defparam ram_block1a46.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a46.port_b_read_enable_clock = "clock1";
defparam ram_block1a46.ram_block_type = "auto";

arriaii_ram_block ram_block1a78(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[78]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a78_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a78.clk0_core_clock_enable = "ena0";
defparam ram_block1a78.clk0_input_clock_enable = "ena2";
defparam ram_block1a78.clk1_core_clock_enable = "ena3";
defparam ram_block1a78.clk1_input_clock_enable = "ena3";
defparam ram_block1a78.clk1_output_clock_enable = "ena1";
defparam ram_block1a78.clock_duty_cycle_dependence = "on";
defparam ram_block1a78.data_interleave_offset_in_bits = 1;
defparam ram_block1a78.data_interleave_width_in_bits = 1;
defparam ram_block1a78.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a78.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a78.operation_mode = "dual_port";
defparam ram_block1a78.port_a_address_clear = "none";
defparam ram_block1a78.port_a_address_width = 8;
defparam ram_block1a78.port_a_data_out_clear = "none";
defparam ram_block1a78.port_a_data_out_clock = "none";
defparam ram_block1a78.port_a_data_width = 1;
defparam ram_block1a78.port_a_first_address = 0;
defparam ram_block1a78.port_a_first_bit_number = 78;
defparam ram_block1a78.port_a_last_address = 255;
defparam ram_block1a78.port_a_logical_ram_depth = 256;
defparam ram_block1a78.port_a_logical_ram_width = 144;
defparam ram_block1a78.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a78.port_b_address_clear = "none";
defparam ram_block1a78.port_b_address_clock = "clock1";
defparam ram_block1a78.port_b_address_width = 8;
defparam ram_block1a78.port_b_data_out_clear = "none";
defparam ram_block1a78.port_b_data_out_clock = "clock1";
defparam ram_block1a78.port_b_data_width = 1;
defparam ram_block1a78.port_b_first_address = 0;
defparam ram_block1a78.port_b_first_bit_number = 78;
defparam ram_block1a78.port_b_last_address = 255;
defparam ram_block1a78.port_b_logical_ram_depth = 256;
defparam ram_block1a78.port_b_logical_ram_width = 144;
defparam ram_block1a78.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a78.port_b_read_enable_clock = "clock1";
defparam ram_block1a78.ram_block_type = "auto";

arriaii_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena2";
defparam ram_block1a14.clk1_core_clock_enable = "ena3";
defparam ram_block1a14.clk1_input_clock_enable = "ena3";
defparam ram_block1a14.clk1_output_clock_enable = "ena1";
defparam ram_block1a14.clock_duty_cycle_dependence = "on";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 8;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 255;
defparam ram_block1a14.port_a_logical_ram_depth = 256;
defparam ram_block1a14.port_a_logical_ram_width = 144;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 8;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 255;
defparam ram_block1a14.port_b_logical_ram_depth = 256;
defparam ram_block1a14.port_b_logical_ram_width = 144;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

arriaii_ram_block ram_block1a111(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[111]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a111_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a111.clk0_core_clock_enable = "ena0";
defparam ram_block1a111.clk0_input_clock_enable = "ena2";
defparam ram_block1a111.clk1_core_clock_enable = "ena3";
defparam ram_block1a111.clk1_input_clock_enable = "ena3";
defparam ram_block1a111.clk1_output_clock_enable = "ena1";
defparam ram_block1a111.clock_duty_cycle_dependence = "on";
defparam ram_block1a111.data_interleave_offset_in_bits = 1;
defparam ram_block1a111.data_interleave_width_in_bits = 1;
defparam ram_block1a111.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a111.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a111.operation_mode = "dual_port";
defparam ram_block1a111.port_a_address_clear = "none";
defparam ram_block1a111.port_a_address_width = 8;
defparam ram_block1a111.port_a_data_out_clear = "none";
defparam ram_block1a111.port_a_data_out_clock = "none";
defparam ram_block1a111.port_a_data_width = 1;
defparam ram_block1a111.port_a_first_address = 0;
defparam ram_block1a111.port_a_first_bit_number = 111;
defparam ram_block1a111.port_a_last_address = 255;
defparam ram_block1a111.port_a_logical_ram_depth = 256;
defparam ram_block1a111.port_a_logical_ram_width = 144;
defparam ram_block1a111.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a111.port_b_address_clear = "none";
defparam ram_block1a111.port_b_address_clock = "clock1";
defparam ram_block1a111.port_b_address_width = 8;
defparam ram_block1a111.port_b_data_out_clear = "none";
defparam ram_block1a111.port_b_data_out_clock = "clock1";
defparam ram_block1a111.port_b_data_width = 1;
defparam ram_block1a111.port_b_first_address = 0;
defparam ram_block1a111.port_b_first_bit_number = 111;
defparam ram_block1a111.port_b_last_address = 255;
defparam ram_block1a111.port_b_logical_ram_depth = 256;
defparam ram_block1a111.port_b_logical_ram_width = 144;
defparam ram_block1a111.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a111.port_b_read_enable_clock = "clock1";
defparam ram_block1a111.ram_block_type = "auto";

arriaii_ram_block ram_block1a47(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[47]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a47_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a47.clk0_core_clock_enable = "ena0";
defparam ram_block1a47.clk0_input_clock_enable = "ena2";
defparam ram_block1a47.clk1_core_clock_enable = "ena3";
defparam ram_block1a47.clk1_input_clock_enable = "ena3";
defparam ram_block1a47.clk1_output_clock_enable = "ena1";
defparam ram_block1a47.clock_duty_cycle_dependence = "on";
defparam ram_block1a47.data_interleave_offset_in_bits = 1;
defparam ram_block1a47.data_interleave_width_in_bits = 1;
defparam ram_block1a47.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a47.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a47.operation_mode = "dual_port";
defparam ram_block1a47.port_a_address_clear = "none";
defparam ram_block1a47.port_a_address_width = 8;
defparam ram_block1a47.port_a_data_out_clear = "none";
defparam ram_block1a47.port_a_data_out_clock = "none";
defparam ram_block1a47.port_a_data_width = 1;
defparam ram_block1a47.port_a_first_address = 0;
defparam ram_block1a47.port_a_first_bit_number = 47;
defparam ram_block1a47.port_a_last_address = 255;
defparam ram_block1a47.port_a_logical_ram_depth = 256;
defparam ram_block1a47.port_a_logical_ram_width = 144;
defparam ram_block1a47.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a47.port_b_address_clear = "none";
defparam ram_block1a47.port_b_address_clock = "clock1";
defparam ram_block1a47.port_b_address_width = 8;
defparam ram_block1a47.port_b_data_out_clear = "none";
defparam ram_block1a47.port_b_data_out_clock = "clock1";
defparam ram_block1a47.port_b_data_width = 1;
defparam ram_block1a47.port_b_first_address = 0;
defparam ram_block1a47.port_b_first_bit_number = 47;
defparam ram_block1a47.port_b_last_address = 255;
defparam ram_block1a47.port_b_logical_ram_depth = 256;
defparam ram_block1a47.port_b_logical_ram_width = 144;
defparam ram_block1a47.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a47.port_b_read_enable_clock = "clock1";
defparam ram_block1a47.ram_block_type = "auto";

arriaii_ram_block ram_block1a79(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[79]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a79_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a79.clk0_core_clock_enable = "ena0";
defparam ram_block1a79.clk0_input_clock_enable = "ena2";
defparam ram_block1a79.clk1_core_clock_enable = "ena3";
defparam ram_block1a79.clk1_input_clock_enable = "ena3";
defparam ram_block1a79.clk1_output_clock_enable = "ena1";
defparam ram_block1a79.clock_duty_cycle_dependence = "on";
defparam ram_block1a79.data_interleave_offset_in_bits = 1;
defparam ram_block1a79.data_interleave_width_in_bits = 1;
defparam ram_block1a79.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a79.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a79.operation_mode = "dual_port";
defparam ram_block1a79.port_a_address_clear = "none";
defparam ram_block1a79.port_a_address_width = 8;
defparam ram_block1a79.port_a_data_out_clear = "none";
defparam ram_block1a79.port_a_data_out_clock = "none";
defparam ram_block1a79.port_a_data_width = 1;
defparam ram_block1a79.port_a_first_address = 0;
defparam ram_block1a79.port_a_first_bit_number = 79;
defparam ram_block1a79.port_a_last_address = 255;
defparam ram_block1a79.port_a_logical_ram_depth = 256;
defparam ram_block1a79.port_a_logical_ram_width = 144;
defparam ram_block1a79.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a79.port_b_address_clear = "none";
defparam ram_block1a79.port_b_address_clock = "clock1";
defparam ram_block1a79.port_b_address_width = 8;
defparam ram_block1a79.port_b_data_out_clear = "none";
defparam ram_block1a79.port_b_data_out_clock = "clock1";
defparam ram_block1a79.port_b_data_width = 1;
defparam ram_block1a79.port_b_first_address = 0;
defparam ram_block1a79.port_b_first_bit_number = 79;
defparam ram_block1a79.port_b_last_address = 255;
defparam ram_block1a79.port_b_logical_ram_depth = 256;
defparam ram_block1a79.port_b_logical_ram_width = 144;
defparam ram_block1a79.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a79.port_b_read_enable_clock = "clock1";
defparam ram_block1a79.ram_block_type = "auto";

arriaii_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena2";
defparam ram_block1a15.clk1_core_clock_enable = "ena3";
defparam ram_block1a15.clk1_input_clock_enable = "ena3";
defparam ram_block1a15.clk1_output_clock_enable = "ena1";
defparam ram_block1a15.clock_duty_cycle_dependence = "on";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 8;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 255;
defparam ram_block1a15.port_a_logical_ram_depth = 256;
defparam ram_block1a15.port_a_logical_ram_width = 144;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 8;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 255;
defparam ram_block1a15.port_b_logical_ram_depth = 256;
defparam ram_block1a15.port_b_logical_ram_width = 144;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

arriaii_ram_block ram_block1a112(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[112]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a112_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a112.clk0_core_clock_enable = "ena0";
defparam ram_block1a112.clk0_input_clock_enable = "ena2";
defparam ram_block1a112.clk1_core_clock_enable = "ena3";
defparam ram_block1a112.clk1_input_clock_enable = "ena3";
defparam ram_block1a112.clk1_output_clock_enable = "ena1";
defparam ram_block1a112.clock_duty_cycle_dependence = "on";
defparam ram_block1a112.data_interleave_offset_in_bits = 1;
defparam ram_block1a112.data_interleave_width_in_bits = 1;
defparam ram_block1a112.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a112.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a112.operation_mode = "dual_port";
defparam ram_block1a112.port_a_address_clear = "none";
defparam ram_block1a112.port_a_address_width = 8;
defparam ram_block1a112.port_a_data_out_clear = "none";
defparam ram_block1a112.port_a_data_out_clock = "none";
defparam ram_block1a112.port_a_data_width = 1;
defparam ram_block1a112.port_a_first_address = 0;
defparam ram_block1a112.port_a_first_bit_number = 112;
defparam ram_block1a112.port_a_last_address = 255;
defparam ram_block1a112.port_a_logical_ram_depth = 256;
defparam ram_block1a112.port_a_logical_ram_width = 144;
defparam ram_block1a112.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a112.port_b_address_clear = "none";
defparam ram_block1a112.port_b_address_clock = "clock1";
defparam ram_block1a112.port_b_address_width = 8;
defparam ram_block1a112.port_b_data_out_clear = "none";
defparam ram_block1a112.port_b_data_out_clock = "clock1";
defparam ram_block1a112.port_b_data_width = 1;
defparam ram_block1a112.port_b_first_address = 0;
defparam ram_block1a112.port_b_first_bit_number = 112;
defparam ram_block1a112.port_b_last_address = 255;
defparam ram_block1a112.port_b_logical_ram_depth = 256;
defparam ram_block1a112.port_b_logical_ram_width = 144;
defparam ram_block1a112.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a112.port_b_read_enable_clock = "clock1";
defparam ram_block1a112.ram_block_type = "auto";

arriaii_ram_block ram_block1a48(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[48]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a48_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a48.clk0_core_clock_enable = "ena0";
defparam ram_block1a48.clk0_input_clock_enable = "ena2";
defparam ram_block1a48.clk1_core_clock_enable = "ena3";
defparam ram_block1a48.clk1_input_clock_enable = "ena3";
defparam ram_block1a48.clk1_output_clock_enable = "ena1";
defparam ram_block1a48.clock_duty_cycle_dependence = "on";
defparam ram_block1a48.data_interleave_offset_in_bits = 1;
defparam ram_block1a48.data_interleave_width_in_bits = 1;
defparam ram_block1a48.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a48.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a48.operation_mode = "dual_port";
defparam ram_block1a48.port_a_address_clear = "none";
defparam ram_block1a48.port_a_address_width = 8;
defparam ram_block1a48.port_a_data_out_clear = "none";
defparam ram_block1a48.port_a_data_out_clock = "none";
defparam ram_block1a48.port_a_data_width = 1;
defparam ram_block1a48.port_a_first_address = 0;
defparam ram_block1a48.port_a_first_bit_number = 48;
defparam ram_block1a48.port_a_last_address = 255;
defparam ram_block1a48.port_a_logical_ram_depth = 256;
defparam ram_block1a48.port_a_logical_ram_width = 144;
defparam ram_block1a48.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a48.port_b_address_clear = "none";
defparam ram_block1a48.port_b_address_clock = "clock1";
defparam ram_block1a48.port_b_address_width = 8;
defparam ram_block1a48.port_b_data_out_clear = "none";
defparam ram_block1a48.port_b_data_out_clock = "clock1";
defparam ram_block1a48.port_b_data_width = 1;
defparam ram_block1a48.port_b_first_address = 0;
defparam ram_block1a48.port_b_first_bit_number = 48;
defparam ram_block1a48.port_b_last_address = 255;
defparam ram_block1a48.port_b_logical_ram_depth = 256;
defparam ram_block1a48.port_b_logical_ram_width = 144;
defparam ram_block1a48.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a48.port_b_read_enable_clock = "clock1";
defparam ram_block1a48.ram_block_type = "auto";

arriaii_ram_block ram_block1a80(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[80]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a80_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a80.clk0_core_clock_enable = "ena0";
defparam ram_block1a80.clk0_input_clock_enable = "ena2";
defparam ram_block1a80.clk1_core_clock_enable = "ena3";
defparam ram_block1a80.clk1_input_clock_enable = "ena3";
defparam ram_block1a80.clk1_output_clock_enable = "ena1";
defparam ram_block1a80.clock_duty_cycle_dependence = "on";
defparam ram_block1a80.data_interleave_offset_in_bits = 1;
defparam ram_block1a80.data_interleave_width_in_bits = 1;
defparam ram_block1a80.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a80.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a80.operation_mode = "dual_port";
defparam ram_block1a80.port_a_address_clear = "none";
defparam ram_block1a80.port_a_address_width = 8;
defparam ram_block1a80.port_a_data_out_clear = "none";
defparam ram_block1a80.port_a_data_out_clock = "none";
defparam ram_block1a80.port_a_data_width = 1;
defparam ram_block1a80.port_a_first_address = 0;
defparam ram_block1a80.port_a_first_bit_number = 80;
defparam ram_block1a80.port_a_last_address = 255;
defparam ram_block1a80.port_a_logical_ram_depth = 256;
defparam ram_block1a80.port_a_logical_ram_width = 144;
defparam ram_block1a80.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a80.port_b_address_clear = "none";
defparam ram_block1a80.port_b_address_clock = "clock1";
defparam ram_block1a80.port_b_address_width = 8;
defparam ram_block1a80.port_b_data_out_clear = "none";
defparam ram_block1a80.port_b_data_out_clock = "clock1";
defparam ram_block1a80.port_b_data_width = 1;
defparam ram_block1a80.port_b_first_address = 0;
defparam ram_block1a80.port_b_first_bit_number = 80;
defparam ram_block1a80.port_b_last_address = 255;
defparam ram_block1a80.port_b_logical_ram_depth = 256;
defparam ram_block1a80.port_b_logical_ram_width = 144;
defparam ram_block1a80.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a80.port_b_read_enable_clock = "clock1";
defparam ram_block1a80.ram_block_type = "auto";

arriaii_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena2";
defparam ram_block1a16.clk1_core_clock_enable = "ena3";
defparam ram_block1a16.clk1_input_clock_enable = "ena3";
defparam ram_block1a16.clk1_output_clock_enable = "ena1";
defparam ram_block1a16.clock_duty_cycle_dependence = "on";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 8;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 255;
defparam ram_block1a16.port_a_logical_ram_depth = 256;
defparam ram_block1a16.port_a_logical_ram_width = 144;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 8;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 255;
defparam ram_block1a16.port_b_logical_ram_depth = 256;
defparam ram_block1a16.port_b_logical_ram_width = 144;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

arriaii_ram_block ram_block1a113(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[113]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a113_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a113.clk0_core_clock_enable = "ena0";
defparam ram_block1a113.clk0_input_clock_enable = "ena2";
defparam ram_block1a113.clk1_core_clock_enable = "ena3";
defparam ram_block1a113.clk1_input_clock_enable = "ena3";
defparam ram_block1a113.clk1_output_clock_enable = "ena1";
defparam ram_block1a113.clock_duty_cycle_dependence = "on";
defparam ram_block1a113.data_interleave_offset_in_bits = 1;
defparam ram_block1a113.data_interleave_width_in_bits = 1;
defparam ram_block1a113.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a113.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a113.operation_mode = "dual_port";
defparam ram_block1a113.port_a_address_clear = "none";
defparam ram_block1a113.port_a_address_width = 8;
defparam ram_block1a113.port_a_data_out_clear = "none";
defparam ram_block1a113.port_a_data_out_clock = "none";
defparam ram_block1a113.port_a_data_width = 1;
defparam ram_block1a113.port_a_first_address = 0;
defparam ram_block1a113.port_a_first_bit_number = 113;
defparam ram_block1a113.port_a_last_address = 255;
defparam ram_block1a113.port_a_logical_ram_depth = 256;
defparam ram_block1a113.port_a_logical_ram_width = 144;
defparam ram_block1a113.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a113.port_b_address_clear = "none";
defparam ram_block1a113.port_b_address_clock = "clock1";
defparam ram_block1a113.port_b_address_width = 8;
defparam ram_block1a113.port_b_data_out_clear = "none";
defparam ram_block1a113.port_b_data_out_clock = "clock1";
defparam ram_block1a113.port_b_data_width = 1;
defparam ram_block1a113.port_b_first_address = 0;
defparam ram_block1a113.port_b_first_bit_number = 113;
defparam ram_block1a113.port_b_last_address = 255;
defparam ram_block1a113.port_b_logical_ram_depth = 256;
defparam ram_block1a113.port_b_logical_ram_width = 144;
defparam ram_block1a113.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a113.port_b_read_enable_clock = "clock1";
defparam ram_block1a113.ram_block_type = "auto";

arriaii_ram_block ram_block1a49(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[49]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a49_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a49.clk0_core_clock_enable = "ena0";
defparam ram_block1a49.clk0_input_clock_enable = "ena2";
defparam ram_block1a49.clk1_core_clock_enable = "ena3";
defparam ram_block1a49.clk1_input_clock_enable = "ena3";
defparam ram_block1a49.clk1_output_clock_enable = "ena1";
defparam ram_block1a49.clock_duty_cycle_dependence = "on";
defparam ram_block1a49.data_interleave_offset_in_bits = 1;
defparam ram_block1a49.data_interleave_width_in_bits = 1;
defparam ram_block1a49.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a49.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a49.operation_mode = "dual_port";
defparam ram_block1a49.port_a_address_clear = "none";
defparam ram_block1a49.port_a_address_width = 8;
defparam ram_block1a49.port_a_data_out_clear = "none";
defparam ram_block1a49.port_a_data_out_clock = "none";
defparam ram_block1a49.port_a_data_width = 1;
defparam ram_block1a49.port_a_first_address = 0;
defparam ram_block1a49.port_a_first_bit_number = 49;
defparam ram_block1a49.port_a_last_address = 255;
defparam ram_block1a49.port_a_logical_ram_depth = 256;
defparam ram_block1a49.port_a_logical_ram_width = 144;
defparam ram_block1a49.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a49.port_b_address_clear = "none";
defparam ram_block1a49.port_b_address_clock = "clock1";
defparam ram_block1a49.port_b_address_width = 8;
defparam ram_block1a49.port_b_data_out_clear = "none";
defparam ram_block1a49.port_b_data_out_clock = "clock1";
defparam ram_block1a49.port_b_data_width = 1;
defparam ram_block1a49.port_b_first_address = 0;
defparam ram_block1a49.port_b_first_bit_number = 49;
defparam ram_block1a49.port_b_last_address = 255;
defparam ram_block1a49.port_b_logical_ram_depth = 256;
defparam ram_block1a49.port_b_logical_ram_width = 144;
defparam ram_block1a49.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a49.port_b_read_enable_clock = "clock1";
defparam ram_block1a49.ram_block_type = "auto";

arriaii_ram_block ram_block1a81(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[81]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a81_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a81.clk0_core_clock_enable = "ena0";
defparam ram_block1a81.clk0_input_clock_enable = "ena2";
defparam ram_block1a81.clk1_core_clock_enable = "ena3";
defparam ram_block1a81.clk1_input_clock_enable = "ena3";
defparam ram_block1a81.clk1_output_clock_enable = "ena1";
defparam ram_block1a81.clock_duty_cycle_dependence = "on";
defparam ram_block1a81.data_interleave_offset_in_bits = 1;
defparam ram_block1a81.data_interleave_width_in_bits = 1;
defparam ram_block1a81.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a81.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a81.operation_mode = "dual_port";
defparam ram_block1a81.port_a_address_clear = "none";
defparam ram_block1a81.port_a_address_width = 8;
defparam ram_block1a81.port_a_data_out_clear = "none";
defparam ram_block1a81.port_a_data_out_clock = "none";
defparam ram_block1a81.port_a_data_width = 1;
defparam ram_block1a81.port_a_first_address = 0;
defparam ram_block1a81.port_a_first_bit_number = 81;
defparam ram_block1a81.port_a_last_address = 255;
defparam ram_block1a81.port_a_logical_ram_depth = 256;
defparam ram_block1a81.port_a_logical_ram_width = 144;
defparam ram_block1a81.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a81.port_b_address_clear = "none";
defparam ram_block1a81.port_b_address_clock = "clock1";
defparam ram_block1a81.port_b_address_width = 8;
defparam ram_block1a81.port_b_data_out_clear = "none";
defparam ram_block1a81.port_b_data_out_clock = "clock1";
defparam ram_block1a81.port_b_data_width = 1;
defparam ram_block1a81.port_b_first_address = 0;
defparam ram_block1a81.port_b_first_bit_number = 81;
defparam ram_block1a81.port_b_last_address = 255;
defparam ram_block1a81.port_b_logical_ram_depth = 256;
defparam ram_block1a81.port_b_logical_ram_width = 144;
defparam ram_block1a81.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a81.port_b_read_enable_clock = "clock1";
defparam ram_block1a81.ram_block_type = "auto";

arriaii_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena2";
defparam ram_block1a17.clk1_core_clock_enable = "ena3";
defparam ram_block1a17.clk1_input_clock_enable = "ena3";
defparam ram_block1a17.clk1_output_clock_enable = "ena1";
defparam ram_block1a17.clock_duty_cycle_dependence = "on";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 8;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 255;
defparam ram_block1a17.port_a_logical_ram_depth = 256;
defparam ram_block1a17.port_a_logical_ram_width = 144;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 8;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 255;
defparam ram_block1a17.port_b_logical_ram_depth = 256;
defparam ram_block1a17.port_b_logical_ram_width = 144;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

arriaii_ram_block ram_block1a114(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[114]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a114_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a114.clk0_core_clock_enable = "ena0";
defparam ram_block1a114.clk0_input_clock_enable = "ena2";
defparam ram_block1a114.clk1_core_clock_enable = "ena3";
defparam ram_block1a114.clk1_input_clock_enable = "ena3";
defparam ram_block1a114.clk1_output_clock_enable = "ena1";
defparam ram_block1a114.clock_duty_cycle_dependence = "on";
defparam ram_block1a114.data_interleave_offset_in_bits = 1;
defparam ram_block1a114.data_interleave_width_in_bits = 1;
defparam ram_block1a114.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a114.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a114.operation_mode = "dual_port";
defparam ram_block1a114.port_a_address_clear = "none";
defparam ram_block1a114.port_a_address_width = 8;
defparam ram_block1a114.port_a_data_out_clear = "none";
defparam ram_block1a114.port_a_data_out_clock = "none";
defparam ram_block1a114.port_a_data_width = 1;
defparam ram_block1a114.port_a_first_address = 0;
defparam ram_block1a114.port_a_first_bit_number = 114;
defparam ram_block1a114.port_a_last_address = 255;
defparam ram_block1a114.port_a_logical_ram_depth = 256;
defparam ram_block1a114.port_a_logical_ram_width = 144;
defparam ram_block1a114.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a114.port_b_address_clear = "none";
defparam ram_block1a114.port_b_address_clock = "clock1";
defparam ram_block1a114.port_b_address_width = 8;
defparam ram_block1a114.port_b_data_out_clear = "none";
defparam ram_block1a114.port_b_data_out_clock = "clock1";
defparam ram_block1a114.port_b_data_width = 1;
defparam ram_block1a114.port_b_first_address = 0;
defparam ram_block1a114.port_b_first_bit_number = 114;
defparam ram_block1a114.port_b_last_address = 255;
defparam ram_block1a114.port_b_logical_ram_depth = 256;
defparam ram_block1a114.port_b_logical_ram_width = 144;
defparam ram_block1a114.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a114.port_b_read_enable_clock = "clock1";
defparam ram_block1a114.ram_block_type = "auto";

arriaii_ram_block ram_block1a50(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[50]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a50_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a50.clk0_core_clock_enable = "ena0";
defparam ram_block1a50.clk0_input_clock_enable = "ena2";
defparam ram_block1a50.clk1_core_clock_enable = "ena3";
defparam ram_block1a50.clk1_input_clock_enable = "ena3";
defparam ram_block1a50.clk1_output_clock_enable = "ena1";
defparam ram_block1a50.clock_duty_cycle_dependence = "on";
defparam ram_block1a50.data_interleave_offset_in_bits = 1;
defparam ram_block1a50.data_interleave_width_in_bits = 1;
defparam ram_block1a50.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a50.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a50.operation_mode = "dual_port";
defparam ram_block1a50.port_a_address_clear = "none";
defparam ram_block1a50.port_a_address_width = 8;
defparam ram_block1a50.port_a_data_out_clear = "none";
defparam ram_block1a50.port_a_data_out_clock = "none";
defparam ram_block1a50.port_a_data_width = 1;
defparam ram_block1a50.port_a_first_address = 0;
defparam ram_block1a50.port_a_first_bit_number = 50;
defparam ram_block1a50.port_a_last_address = 255;
defparam ram_block1a50.port_a_logical_ram_depth = 256;
defparam ram_block1a50.port_a_logical_ram_width = 144;
defparam ram_block1a50.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a50.port_b_address_clear = "none";
defparam ram_block1a50.port_b_address_clock = "clock1";
defparam ram_block1a50.port_b_address_width = 8;
defparam ram_block1a50.port_b_data_out_clear = "none";
defparam ram_block1a50.port_b_data_out_clock = "clock1";
defparam ram_block1a50.port_b_data_width = 1;
defparam ram_block1a50.port_b_first_address = 0;
defparam ram_block1a50.port_b_first_bit_number = 50;
defparam ram_block1a50.port_b_last_address = 255;
defparam ram_block1a50.port_b_logical_ram_depth = 256;
defparam ram_block1a50.port_b_logical_ram_width = 144;
defparam ram_block1a50.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a50.port_b_read_enable_clock = "clock1";
defparam ram_block1a50.ram_block_type = "auto";

arriaii_ram_block ram_block1a82(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[82]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a82_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a82.clk0_core_clock_enable = "ena0";
defparam ram_block1a82.clk0_input_clock_enable = "ena2";
defparam ram_block1a82.clk1_core_clock_enable = "ena3";
defparam ram_block1a82.clk1_input_clock_enable = "ena3";
defparam ram_block1a82.clk1_output_clock_enable = "ena1";
defparam ram_block1a82.clock_duty_cycle_dependence = "on";
defparam ram_block1a82.data_interleave_offset_in_bits = 1;
defparam ram_block1a82.data_interleave_width_in_bits = 1;
defparam ram_block1a82.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a82.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a82.operation_mode = "dual_port";
defparam ram_block1a82.port_a_address_clear = "none";
defparam ram_block1a82.port_a_address_width = 8;
defparam ram_block1a82.port_a_data_out_clear = "none";
defparam ram_block1a82.port_a_data_out_clock = "none";
defparam ram_block1a82.port_a_data_width = 1;
defparam ram_block1a82.port_a_first_address = 0;
defparam ram_block1a82.port_a_first_bit_number = 82;
defparam ram_block1a82.port_a_last_address = 255;
defparam ram_block1a82.port_a_logical_ram_depth = 256;
defparam ram_block1a82.port_a_logical_ram_width = 144;
defparam ram_block1a82.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a82.port_b_address_clear = "none";
defparam ram_block1a82.port_b_address_clock = "clock1";
defparam ram_block1a82.port_b_address_width = 8;
defparam ram_block1a82.port_b_data_out_clear = "none";
defparam ram_block1a82.port_b_data_out_clock = "clock1";
defparam ram_block1a82.port_b_data_width = 1;
defparam ram_block1a82.port_b_first_address = 0;
defparam ram_block1a82.port_b_first_bit_number = 82;
defparam ram_block1a82.port_b_last_address = 255;
defparam ram_block1a82.port_b_logical_ram_depth = 256;
defparam ram_block1a82.port_b_logical_ram_width = 144;
defparam ram_block1a82.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a82.port_b_read_enable_clock = "clock1";
defparam ram_block1a82.ram_block_type = "auto";

arriaii_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena2";
defparam ram_block1a18.clk1_core_clock_enable = "ena3";
defparam ram_block1a18.clk1_input_clock_enable = "ena3";
defparam ram_block1a18.clk1_output_clock_enable = "ena1";
defparam ram_block1a18.clock_duty_cycle_dependence = "on";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 8;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 255;
defparam ram_block1a18.port_a_logical_ram_depth = 256;
defparam ram_block1a18.port_a_logical_ram_width = 144;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 8;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 255;
defparam ram_block1a18.port_b_logical_ram_depth = 256;
defparam ram_block1a18.port_b_logical_ram_width = 144;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

arriaii_ram_block ram_block1a115(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[115]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a115_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a115.clk0_core_clock_enable = "ena0";
defparam ram_block1a115.clk0_input_clock_enable = "ena2";
defparam ram_block1a115.clk1_core_clock_enable = "ena3";
defparam ram_block1a115.clk1_input_clock_enable = "ena3";
defparam ram_block1a115.clk1_output_clock_enable = "ena1";
defparam ram_block1a115.clock_duty_cycle_dependence = "on";
defparam ram_block1a115.data_interleave_offset_in_bits = 1;
defparam ram_block1a115.data_interleave_width_in_bits = 1;
defparam ram_block1a115.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a115.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a115.operation_mode = "dual_port";
defparam ram_block1a115.port_a_address_clear = "none";
defparam ram_block1a115.port_a_address_width = 8;
defparam ram_block1a115.port_a_data_out_clear = "none";
defparam ram_block1a115.port_a_data_out_clock = "none";
defparam ram_block1a115.port_a_data_width = 1;
defparam ram_block1a115.port_a_first_address = 0;
defparam ram_block1a115.port_a_first_bit_number = 115;
defparam ram_block1a115.port_a_last_address = 255;
defparam ram_block1a115.port_a_logical_ram_depth = 256;
defparam ram_block1a115.port_a_logical_ram_width = 144;
defparam ram_block1a115.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a115.port_b_address_clear = "none";
defparam ram_block1a115.port_b_address_clock = "clock1";
defparam ram_block1a115.port_b_address_width = 8;
defparam ram_block1a115.port_b_data_out_clear = "none";
defparam ram_block1a115.port_b_data_out_clock = "clock1";
defparam ram_block1a115.port_b_data_width = 1;
defparam ram_block1a115.port_b_first_address = 0;
defparam ram_block1a115.port_b_first_bit_number = 115;
defparam ram_block1a115.port_b_last_address = 255;
defparam ram_block1a115.port_b_logical_ram_depth = 256;
defparam ram_block1a115.port_b_logical_ram_width = 144;
defparam ram_block1a115.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a115.port_b_read_enable_clock = "clock1";
defparam ram_block1a115.ram_block_type = "auto";

arriaii_ram_block ram_block1a51(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[51]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a51_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a51.clk0_core_clock_enable = "ena0";
defparam ram_block1a51.clk0_input_clock_enable = "ena2";
defparam ram_block1a51.clk1_core_clock_enable = "ena3";
defparam ram_block1a51.clk1_input_clock_enable = "ena3";
defparam ram_block1a51.clk1_output_clock_enable = "ena1";
defparam ram_block1a51.clock_duty_cycle_dependence = "on";
defparam ram_block1a51.data_interleave_offset_in_bits = 1;
defparam ram_block1a51.data_interleave_width_in_bits = 1;
defparam ram_block1a51.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a51.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a51.operation_mode = "dual_port";
defparam ram_block1a51.port_a_address_clear = "none";
defparam ram_block1a51.port_a_address_width = 8;
defparam ram_block1a51.port_a_data_out_clear = "none";
defparam ram_block1a51.port_a_data_out_clock = "none";
defparam ram_block1a51.port_a_data_width = 1;
defparam ram_block1a51.port_a_first_address = 0;
defparam ram_block1a51.port_a_first_bit_number = 51;
defparam ram_block1a51.port_a_last_address = 255;
defparam ram_block1a51.port_a_logical_ram_depth = 256;
defparam ram_block1a51.port_a_logical_ram_width = 144;
defparam ram_block1a51.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a51.port_b_address_clear = "none";
defparam ram_block1a51.port_b_address_clock = "clock1";
defparam ram_block1a51.port_b_address_width = 8;
defparam ram_block1a51.port_b_data_out_clear = "none";
defparam ram_block1a51.port_b_data_out_clock = "clock1";
defparam ram_block1a51.port_b_data_width = 1;
defparam ram_block1a51.port_b_first_address = 0;
defparam ram_block1a51.port_b_first_bit_number = 51;
defparam ram_block1a51.port_b_last_address = 255;
defparam ram_block1a51.port_b_logical_ram_depth = 256;
defparam ram_block1a51.port_b_logical_ram_width = 144;
defparam ram_block1a51.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a51.port_b_read_enable_clock = "clock1";
defparam ram_block1a51.ram_block_type = "auto";

arriaii_ram_block ram_block1a83(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[83]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a83_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a83.clk0_core_clock_enable = "ena0";
defparam ram_block1a83.clk0_input_clock_enable = "ena2";
defparam ram_block1a83.clk1_core_clock_enable = "ena3";
defparam ram_block1a83.clk1_input_clock_enable = "ena3";
defparam ram_block1a83.clk1_output_clock_enable = "ena1";
defparam ram_block1a83.clock_duty_cycle_dependence = "on";
defparam ram_block1a83.data_interleave_offset_in_bits = 1;
defparam ram_block1a83.data_interleave_width_in_bits = 1;
defparam ram_block1a83.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a83.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a83.operation_mode = "dual_port";
defparam ram_block1a83.port_a_address_clear = "none";
defparam ram_block1a83.port_a_address_width = 8;
defparam ram_block1a83.port_a_data_out_clear = "none";
defparam ram_block1a83.port_a_data_out_clock = "none";
defparam ram_block1a83.port_a_data_width = 1;
defparam ram_block1a83.port_a_first_address = 0;
defparam ram_block1a83.port_a_first_bit_number = 83;
defparam ram_block1a83.port_a_last_address = 255;
defparam ram_block1a83.port_a_logical_ram_depth = 256;
defparam ram_block1a83.port_a_logical_ram_width = 144;
defparam ram_block1a83.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a83.port_b_address_clear = "none";
defparam ram_block1a83.port_b_address_clock = "clock1";
defparam ram_block1a83.port_b_address_width = 8;
defparam ram_block1a83.port_b_data_out_clear = "none";
defparam ram_block1a83.port_b_data_out_clock = "clock1";
defparam ram_block1a83.port_b_data_width = 1;
defparam ram_block1a83.port_b_first_address = 0;
defparam ram_block1a83.port_b_first_bit_number = 83;
defparam ram_block1a83.port_b_last_address = 255;
defparam ram_block1a83.port_b_logical_ram_depth = 256;
defparam ram_block1a83.port_b_logical_ram_width = 144;
defparam ram_block1a83.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a83.port_b_read_enable_clock = "clock1";
defparam ram_block1a83.ram_block_type = "auto";

arriaii_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena2";
defparam ram_block1a19.clk1_core_clock_enable = "ena3";
defparam ram_block1a19.clk1_input_clock_enable = "ena3";
defparam ram_block1a19.clk1_output_clock_enable = "ena1";
defparam ram_block1a19.clock_duty_cycle_dependence = "on";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 8;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 255;
defparam ram_block1a19.port_a_logical_ram_depth = 256;
defparam ram_block1a19.port_a_logical_ram_width = 144;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 8;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "clock1";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 255;
defparam ram_block1a19.port_b_logical_ram_depth = 256;
defparam ram_block1a19.port_b_logical_ram_width = 144;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

arriaii_ram_block ram_block1a116(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[116]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a116_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a116.clk0_core_clock_enable = "ena0";
defparam ram_block1a116.clk0_input_clock_enable = "ena2";
defparam ram_block1a116.clk1_core_clock_enable = "ena3";
defparam ram_block1a116.clk1_input_clock_enable = "ena3";
defparam ram_block1a116.clk1_output_clock_enable = "ena1";
defparam ram_block1a116.clock_duty_cycle_dependence = "on";
defparam ram_block1a116.data_interleave_offset_in_bits = 1;
defparam ram_block1a116.data_interleave_width_in_bits = 1;
defparam ram_block1a116.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a116.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a116.operation_mode = "dual_port";
defparam ram_block1a116.port_a_address_clear = "none";
defparam ram_block1a116.port_a_address_width = 8;
defparam ram_block1a116.port_a_data_out_clear = "none";
defparam ram_block1a116.port_a_data_out_clock = "none";
defparam ram_block1a116.port_a_data_width = 1;
defparam ram_block1a116.port_a_first_address = 0;
defparam ram_block1a116.port_a_first_bit_number = 116;
defparam ram_block1a116.port_a_last_address = 255;
defparam ram_block1a116.port_a_logical_ram_depth = 256;
defparam ram_block1a116.port_a_logical_ram_width = 144;
defparam ram_block1a116.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a116.port_b_address_clear = "none";
defparam ram_block1a116.port_b_address_clock = "clock1";
defparam ram_block1a116.port_b_address_width = 8;
defparam ram_block1a116.port_b_data_out_clear = "none";
defparam ram_block1a116.port_b_data_out_clock = "clock1";
defparam ram_block1a116.port_b_data_width = 1;
defparam ram_block1a116.port_b_first_address = 0;
defparam ram_block1a116.port_b_first_bit_number = 116;
defparam ram_block1a116.port_b_last_address = 255;
defparam ram_block1a116.port_b_logical_ram_depth = 256;
defparam ram_block1a116.port_b_logical_ram_width = 144;
defparam ram_block1a116.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a116.port_b_read_enable_clock = "clock1";
defparam ram_block1a116.ram_block_type = "auto";

arriaii_ram_block ram_block1a52(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[52]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a52_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a52.clk0_core_clock_enable = "ena0";
defparam ram_block1a52.clk0_input_clock_enable = "ena2";
defparam ram_block1a52.clk1_core_clock_enable = "ena3";
defparam ram_block1a52.clk1_input_clock_enable = "ena3";
defparam ram_block1a52.clk1_output_clock_enable = "ena1";
defparam ram_block1a52.clock_duty_cycle_dependence = "on";
defparam ram_block1a52.data_interleave_offset_in_bits = 1;
defparam ram_block1a52.data_interleave_width_in_bits = 1;
defparam ram_block1a52.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a52.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a52.operation_mode = "dual_port";
defparam ram_block1a52.port_a_address_clear = "none";
defparam ram_block1a52.port_a_address_width = 8;
defparam ram_block1a52.port_a_data_out_clear = "none";
defparam ram_block1a52.port_a_data_out_clock = "none";
defparam ram_block1a52.port_a_data_width = 1;
defparam ram_block1a52.port_a_first_address = 0;
defparam ram_block1a52.port_a_first_bit_number = 52;
defparam ram_block1a52.port_a_last_address = 255;
defparam ram_block1a52.port_a_logical_ram_depth = 256;
defparam ram_block1a52.port_a_logical_ram_width = 144;
defparam ram_block1a52.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a52.port_b_address_clear = "none";
defparam ram_block1a52.port_b_address_clock = "clock1";
defparam ram_block1a52.port_b_address_width = 8;
defparam ram_block1a52.port_b_data_out_clear = "none";
defparam ram_block1a52.port_b_data_out_clock = "clock1";
defparam ram_block1a52.port_b_data_width = 1;
defparam ram_block1a52.port_b_first_address = 0;
defparam ram_block1a52.port_b_first_bit_number = 52;
defparam ram_block1a52.port_b_last_address = 255;
defparam ram_block1a52.port_b_logical_ram_depth = 256;
defparam ram_block1a52.port_b_logical_ram_width = 144;
defparam ram_block1a52.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a52.port_b_read_enable_clock = "clock1";
defparam ram_block1a52.ram_block_type = "auto";

arriaii_ram_block ram_block1a84(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[84]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a84_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a84.clk0_core_clock_enable = "ena0";
defparam ram_block1a84.clk0_input_clock_enable = "ena2";
defparam ram_block1a84.clk1_core_clock_enable = "ena3";
defparam ram_block1a84.clk1_input_clock_enable = "ena3";
defparam ram_block1a84.clk1_output_clock_enable = "ena1";
defparam ram_block1a84.clock_duty_cycle_dependence = "on";
defparam ram_block1a84.data_interleave_offset_in_bits = 1;
defparam ram_block1a84.data_interleave_width_in_bits = 1;
defparam ram_block1a84.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a84.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a84.operation_mode = "dual_port";
defparam ram_block1a84.port_a_address_clear = "none";
defparam ram_block1a84.port_a_address_width = 8;
defparam ram_block1a84.port_a_data_out_clear = "none";
defparam ram_block1a84.port_a_data_out_clock = "none";
defparam ram_block1a84.port_a_data_width = 1;
defparam ram_block1a84.port_a_first_address = 0;
defparam ram_block1a84.port_a_first_bit_number = 84;
defparam ram_block1a84.port_a_last_address = 255;
defparam ram_block1a84.port_a_logical_ram_depth = 256;
defparam ram_block1a84.port_a_logical_ram_width = 144;
defparam ram_block1a84.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a84.port_b_address_clear = "none";
defparam ram_block1a84.port_b_address_clock = "clock1";
defparam ram_block1a84.port_b_address_width = 8;
defparam ram_block1a84.port_b_data_out_clear = "none";
defparam ram_block1a84.port_b_data_out_clock = "clock1";
defparam ram_block1a84.port_b_data_width = 1;
defparam ram_block1a84.port_b_first_address = 0;
defparam ram_block1a84.port_b_first_bit_number = 84;
defparam ram_block1a84.port_b_last_address = 255;
defparam ram_block1a84.port_b_logical_ram_depth = 256;
defparam ram_block1a84.port_b_logical_ram_width = 144;
defparam ram_block1a84.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a84.port_b_read_enable_clock = "clock1";
defparam ram_block1a84.ram_block_type = "auto";

arriaii_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena2";
defparam ram_block1a20.clk1_core_clock_enable = "ena3";
defparam ram_block1a20.clk1_input_clock_enable = "ena3";
defparam ram_block1a20.clk1_output_clock_enable = "ena1";
defparam ram_block1a20.clock_duty_cycle_dependence = "on";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 8;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 255;
defparam ram_block1a20.port_a_logical_ram_depth = 256;
defparam ram_block1a20.port_a_logical_ram_width = 144;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 8;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "clock1";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 255;
defparam ram_block1a20.port_b_logical_ram_depth = 256;
defparam ram_block1a20.port_b_logical_ram_width = 144;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

arriaii_ram_block ram_block1a117(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[117]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a117_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a117.clk0_core_clock_enable = "ena0";
defparam ram_block1a117.clk0_input_clock_enable = "ena2";
defparam ram_block1a117.clk1_core_clock_enable = "ena3";
defparam ram_block1a117.clk1_input_clock_enable = "ena3";
defparam ram_block1a117.clk1_output_clock_enable = "ena1";
defparam ram_block1a117.clock_duty_cycle_dependence = "on";
defparam ram_block1a117.data_interleave_offset_in_bits = 1;
defparam ram_block1a117.data_interleave_width_in_bits = 1;
defparam ram_block1a117.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a117.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a117.operation_mode = "dual_port";
defparam ram_block1a117.port_a_address_clear = "none";
defparam ram_block1a117.port_a_address_width = 8;
defparam ram_block1a117.port_a_data_out_clear = "none";
defparam ram_block1a117.port_a_data_out_clock = "none";
defparam ram_block1a117.port_a_data_width = 1;
defparam ram_block1a117.port_a_first_address = 0;
defparam ram_block1a117.port_a_first_bit_number = 117;
defparam ram_block1a117.port_a_last_address = 255;
defparam ram_block1a117.port_a_logical_ram_depth = 256;
defparam ram_block1a117.port_a_logical_ram_width = 144;
defparam ram_block1a117.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a117.port_b_address_clear = "none";
defparam ram_block1a117.port_b_address_clock = "clock1";
defparam ram_block1a117.port_b_address_width = 8;
defparam ram_block1a117.port_b_data_out_clear = "none";
defparam ram_block1a117.port_b_data_out_clock = "clock1";
defparam ram_block1a117.port_b_data_width = 1;
defparam ram_block1a117.port_b_first_address = 0;
defparam ram_block1a117.port_b_first_bit_number = 117;
defparam ram_block1a117.port_b_last_address = 255;
defparam ram_block1a117.port_b_logical_ram_depth = 256;
defparam ram_block1a117.port_b_logical_ram_width = 144;
defparam ram_block1a117.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a117.port_b_read_enable_clock = "clock1";
defparam ram_block1a117.ram_block_type = "auto";

arriaii_ram_block ram_block1a53(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[53]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a53_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a53.clk0_core_clock_enable = "ena0";
defparam ram_block1a53.clk0_input_clock_enable = "ena2";
defparam ram_block1a53.clk1_core_clock_enable = "ena3";
defparam ram_block1a53.clk1_input_clock_enable = "ena3";
defparam ram_block1a53.clk1_output_clock_enable = "ena1";
defparam ram_block1a53.clock_duty_cycle_dependence = "on";
defparam ram_block1a53.data_interleave_offset_in_bits = 1;
defparam ram_block1a53.data_interleave_width_in_bits = 1;
defparam ram_block1a53.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a53.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a53.operation_mode = "dual_port";
defparam ram_block1a53.port_a_address_clear = "none";
defparam ram_block1a53.port_a_address_width = 8;
defparam ram_block1a53.port_a_data_out_clear = "none";
defparam ram_block1a53.port_a_data_out_clock = "none";
defparam ram_block1a53.port_a_data_width = 1;
defparam ram_block1a53.port_a_first_address = 0;
defparam ram_block1a53.port_a_first_bit_number = 53;
defparam ram_block1a53.port_a_last_address = 255;
defparam ram_block1a53.port_a_logical_ram_depth = 256;
defparam ram_block1a53.port_a_logical_ram_width = 144;
defparam ram_block1a53.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a53.port_b_address_clear = "none";
defparam ram_block1a53.port_b_address_clock = "clock1";
defparam ram_block1a53.port_b_address_width = 8;
defparam ram_block1a53.port_b_data_out_clear = "none";
defparam ram_block1a53.port_b_data_out_clock = "clock1";
defparam ram_block1a53.port_b_data_width = 1;
defparam ram_block1a53.port_b_first_address = 0;
defparam ram_block1a53.port_b_first_bit_number = 53;
defparam ram_block1a53.port_b_last_address = 255;
defparam ram_block1a53.port_b_logical_ram_depth = 256;
defparam ram_block1a53.port_b_logical_ram_width = 144;
defparam ram_block1a53.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a53.port_b_read_enable_clock = "clock1";
defparam ram_block1a53.ram_block_type = "auto";

arriaii_ram_block ram_block1a85(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[85]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a85_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a85.clk0_core_clock_enable = "ena0";
defparam ram_block1a85.clk0_input_clock_enable = "ena2";
defparam ram_block1a85.clk1_core_clock_enable = "ena3";
defparam ram_block1a85.clk1_input_clock_enable = "ena3";
defparam ram_block1a85.clk1_output_clock_enable = "ena1";
defparam ram_block1a85.clock_duty_cycle_dependence = "on";
defparam ram_block1a85.data_interleave_offset_in_bits = 1;
defparam ram_block1a85.data_interleave_width_in_bits = 1;
defparam ram_block1a85.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a85.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a85.operation_mode = "dual_port";
defparam ram_block1a85.port_a_address_clear = "none";
defparam ram_block1a85.port_a_address_width = 8;
defparam ram_block1a85.port_a_data_out_clear = "none";
defparam ram_block1a85.port_a_data_out_clock = "none";
defparam ram_block1a85.port_a_data_width = 1;
defparam ram_block1a85.port_a_first_address = 0;
defparam ram_block1a85.port_a_first_bit_number = 85;
defparam ram_block1a85.port_a_last_address = 255;
defparam ram_block1a85.port_a_logical_ram_depth = 256;
defparam ram_block1a85.port_a_logical_ram_width = 144;
defparam ram_block1a85.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a85.port_b_address_clear = "none";
defparam ram_block1a85.port_b_address_clock = "clock1";
defparam ram_block1a85.port_b_address_width = 8;
defparam ram_block1a85.port_b_data_out_clear = "none";
defparam ram_block1a85.port_b_data_out_clock = "clock1";
defparam ram_block1a85.port_b_data_width = 1;
defparam ram_block1a85.port_b_first_address = 0;
defparam ram_block1a85.port_b_first_bit_number = 85;
defparam ram_block1a85.port_b_last_address = 255;
defparam ram_block1a85.port_b_logical_ram_depth = 256;
defparam ram_block1a85.port_b_logical_ram_width = 144;
defparam ram_block1a85.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a85.port_b_read_enable_clock = "clock1";
defparam ram_block1a85.ram_block_type = "auto";

arriaii_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena2";
defparam ram_block1a21.clk1_core_clock_enable = "ena3";
defparam ram_block1a21.clk1_input_clock_enable = "ena3";
defparam ram_block1a21.clk1_output_clock_enable = "ena1";
defparam ram_block1a21.clock_duty_cycle_dependence = "on";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 8;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 255;
defparam ram_block1a21.port_a_logical_ram_depth = 256;
defparam ram_block1a21.port_a_logical_ram_width = 144;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 8;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "clock1";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 255;
defparam ram_block1a21.port_b_logical_ram_depth = 256;
defparam ram_block1a21.port_b_logical_ram_width = 144;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

arriaii_ram_block ram_block1a118(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[118]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a118_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a118.clk0_core_clock_enable = "ena0";
defparam ram_block1a118.clk0_input_clock_enable = "ena2";
defparam ram_block1a118.clk1_core_clock_enable = "ena3";
defparam ram_block1a118.clk1_input_clock_enable = "ena3";
defparam ram_block1a118.clk1_output_clock_enable = "ena1";
defparam ram_block1a118.clock_duty_cycle_dependence = "on";
defparam ram_block1a118.data_interleave_offset_in_bits = 1;
defparam ram_block1a118.data_interleave_width_in_bits = 1;
defparam ram_block1a118.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a118.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a118.operation_mode = "dual_port";
defparam ram_block1a118.port_a_address_clear = "none";
defparam ram_block1a118.port_a_address_width = 8;
defparam ram_block1a118.port_a_data_out_clear = "none";
defparam ram_block1a118.port_a_data_out_clock = "none";
defparam ram_block1a118.port_a_data_width = 1;
defparam ram_block1a118.port_a_first_address = 0;
defparam ram_block1a118.port_a_first_bit_number = 118;
defparam ram_block1a118.port_a_last_address = 255;
defparam ram_block1a118.port_a_logical_ram_depth = 256;
defparam ram_block1a118.port_a_logical_ram_width = 144;
defparam ram_block1a118.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a118.port_b_address_clear = "none";
defparam ram_block1a118.port_b_address_clock = "clock1";
defparam ram_block1a118.port_b_address_width = 8;
defparam ram_block1a118.port_b_data_out_clear = "none";
defparam ram_block1a118.port_b_data_out_clock = "clock1";
defparam ram_block1a118.port_b_data_width = 1;
defparam ram_block1a118.port_b_first_address = 0;
defparam ram_block1a118.port_b_first_bit_number = 118;
defparam ram_block1a118.port_b_last_address = 255;
defparam ram_block1a118.port_b_logical_ram_depth = 256;
defparam ram_block1a118.port_b_logical_ram_width = 144;
defparam ram_block1a118.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a118.port_b_read_enable_clock = "clock1";
defparam ram_block1a118.ram_block_type = "auto";

arriaii_ram_block ram_block1a54(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[54]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a54_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a54.clk0_core_clock_enable = "ena0";
defparam ram_block1a54.clk0_input_clock_enable = "ena2";
defparam ram_block1a54.clk1_core_clock_enable = "ena3";
defparam ram_block1a54.clk1_input_clock_enable = "ena3";
defparam ram_block1a54.clk1_output_clock_enable = "ena1";
defparam ram_block1a54.clock_duty_cycle_dependence = "on";
defparam ram_block1a54.data_interleave_offset_in_bits = 1;
defparam ram_block1a54.data_interleave_width_in_bits = 1;
defparam ram_block1a54.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a54.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a54.operation_mode = "dual_port";
defparam ram_block1a54.port_a_address_clear = "none";
defparam ram_block1a54.port_a_address_width = 8;
defparam ram_block1a54.port_a_data_out_clear = "none";
defparam ram_block1a54.port_a_data_out_clock = "none";
defparam ram_block1a54.port_a_data_width = 1;
defparam ram_block1a54.port_a_first_address = 0;
defparam ram_block1a54.port_a_first_bit_number = 54;
defparam ram_block1a54.port_a_last_address = 255;
defparam ram_block1a54.port_a_logical_ram_depth = 256;
defparam ram_block1a54.port_a_logical_ram_width = 144;
defparam ram_block1a54.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a54.port_b_address_clear = "none";
defparam ram_block1a54.port_b_address_clock = "clock1";
defparam ram_block1a54.port_b_address_width = 8;
defparam ram_block1a54.port_b_data_out_clear = "none";
defparam ram_block1a54.port_b_data_out_clock = "clock1";
defparam ram_block1a54.port_b_data_width = 1;
defparam ram_block1a54.port_b_first_address = 0;
defparam ram_block1a54.port_b_first_bit_number = 54;
defparam ram_block1a54.port_b_last_address = 255;
defparam ram_block1a54.port_b_logical_ram_depth = 256;
defparam ram_block1a54.port_b_logical_ram_width = 144;
defparam ram_block1a54.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a54.port_b_read_enable_clock = "clock1";
defparam ram_block1a54.ram_block_type = "auto";

arriaii_ram_block ram_block1a86(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[86]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a86_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a86.clk0_core_clock_enable = "ena0";
defparam ram_block1a86.clk0_input_clock_enable = "ena2";
defparam ram_block1a86.clk1_core_clock_enable = "ena3";
defparam ram_block1a86.clk1_input_clock_enable = "ena3";
defparam ram_block1a86.clk1_output_clock_enable = "ena1";
defparam ram_block1a86.clock_duty_cycle_dependence = "on";
defparam ram_block1a86.data_interleave_offset_in_bits = 1;
defparam ram_block1a86.data_interleave_width_in_bits = 1;
defparam ram_block1a86.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a86.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a86.operation_mode = "dual_port";
defparam ram_block1a86.port_a_address_clear = "none";
defparam ram_block1a86.port_a_address_width = 8;
defparam ram_block1a86.port_a_data_out_clear = "none";
defparam ram_block1a86.port_a_data_out_clock = "none";
defparam ram_block1a86.port_a_data_width = 1;
defparam ram_block1a86.port_a_first_address = 0;
defparam ram_block1a86.port_a_first_bit_number = 86;
defparam ram_block1a86.port_a_last_address = 255;
defparam ram_block1a86.port_a_logical_ram_depth = 256;
defparam ram_block1a86.port_a_logical_ram_width = 144;
defparam ram_block1a86.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a86.port_b_address_clear = "none";
defparam ram_block1a86.port_b_address_clock = "clock1";
defparam ram_block1a86.port_b_address_width = 8;
defparam ram_block1a86.port_b_data_out_clear = "none";
defparam ram_block1a86.port_b_data_out_clock = "clock1";
defparam ram_block1a86.port_b_data_width = 1;
defparam ram_block1a86.port_b_first_address = 0;
defparam ram_block1a86.port_b_first_bit_number = 86;
defparam ram_block1a86.port_b_last_address = 255;
defparam ram_block1a86.port_b_logical_ram_depth = 256;
defparam ram_block1a86.port_b_logical_ram_width = 144;
defparam ram_block1a86.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a86.port_b_read_enable_clock = "clock1";
defparam ram_block1a86.ram_block_type = "auto";

arriaii_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena2";
defparam ram_block1a22.clk1_core_clock_enable = "ena3";
defparam ram_block1a22.clk1_input_clock_enable = "ena3";
defparam ram_block1a22.clk1_output_clock_enable = "ena1";
defparam ram_block1a22.clock_duty_cycle_dependence = "on";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 8;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 255;
defparam ram_block1a22.port_a_logical_ram_depth = 256;
defparam ram_block1a22.port_a_logical_ram_width = 144;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock1";
defparam ram_block1a22.port_b_address_width = 8;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "clock1";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 255;
defparam ram_block1a22.port_b_logical_ram_depth = 256;
defparam ram_block1a22.port_b_logical_ram_width = 144;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock1";
defparam ram_block1a22.ram_block_type = "auto";

arriaii_ram_block ram_block1a119(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[119]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a119_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a119.clk0_core_clock_enable = "ena0";
defparam ram_block1a119.clk0_input_clock_enable = "ena2";
defparam ram_block1a119.clk1_core_clock_enable = "ena3";
defparam ram_block1a119.clk1_input_clock_enable = "ena3";
defparam ram_block1a119.clk1_output_clock_enable = "ena1";
defparam ram_block1a119.clock_duty_cycle_dependence = "on";
defparam ram_block1a119.data_interleave_offset_in_bits = 1;
defparam ram_block1a119.data_interleave_width_in_bits = 1;
defparam ram_block1a119.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a119.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a119.operation_mode = "dual_port";
defparam ram_block1a119.port_a_address_clear = "none";
defparam ram_block1a119.port_a_address_width = 8;
defparam ram_block1a119.port_a_data_out_clear = "none";
defparam ram_block1a119.port_a_data_out_clock = "none";
defparam ram_block1a119.port_a_data_width = 1;
defparam ram_block1a119.port_a_first_address = 0;
defparam ram_block1a119.port_a_first_bit_number = 119;
defparam ram_block1a119.port_a_last_address = 255;
defparam ram_block1a119.port_a_logical_ram_depth = 256;
defparam ram_block1a119.port_a_logical_ram_width = 144;
defparam ram_block1a119.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a119.port_b_address_clear = "none";
defparam ram_block1a119.port_b_address_clock = "clock1";
defparam ram_block1a119.port_b_address_width = 8;
defparam ram_block1a119.port_b_data_out_clear = "none";
defparam ram_block1a119.port_b_data_out_clock = "clock1";
defparam ram_block1a119.port_b_data_width = 1;
defparam ram_block1a119.port_b_first_address = 0;
defparam ram_block1a119.port_b_first_bit_number = 119;
defparam ram_block1a119.port_b_last_address = 255;
defparam ram_block1a119.port_b_logical_ram_depth = 256;
defparam ram_block1a119.port_b_logical_ram_width = 144;
defparam ram_block1a119.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a119.port_b_read_enable_clock = "clock1";
defparam ram_block1a119.ram_block_type = "auto";

arriaii_ram_block ram_block1a55(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[55]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a55_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a55.clk0_core_clock_enable = "ena0";
defparam ram_block1a55.clk0_input_clock_enable = "ena2";
defparam ram_block1a55.clk1_core_clock_enable = "ena3";
defparam ram_block1a55.clk1_input_clock_enable = "ena3";
defparam ram_block1a55.clk1_output_clock_enable = "ena1";
defparam ram_block1a55.clock_duty_cycle_dependence = "on";
defparam ram_block1a55.data_interleave_offset_in_bits = 1;
defparam ram_block1a55.data_interleave_width_in_bits = 1;
defparam ram_block1a55.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a55.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a55.operation_mode = "dual_port";
defparam ram_block1a55.port_a_address_clear = "none";
defparam ram_block1a55.port_a_address_width = 8;
defparam ram_block1a55.port_a_data_out_clear = "none";
defparam ram_block1a55.port_a_data_out_clock = "none";
defparam ram_block1a55.port_a_data_width = 1;
defparam ram_block1a55.port_a_first_address = 0;
defparam ram_block1a55.port_a_first_bit_number = 55;
defparam ram_block1a55.port_a_last_address = 255;
defparam ram_block1a55.port_a_logical_ram_depth = 256;
defparam ram_block1a55.port_a_logical_ram_width = 144;
defparam ram_block1a55.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a55.port_b_address_clear = "none";
defparam ram_block1a55.port_b_address_clock = "clock1";
defparam ram_block1a55.port_b_address_width = 8;
defparam ram_block1a55.port_b_data_out_clear = "none";
defparam ram_block1a55.port_b_data_out_clock = "clock1";
defparam ram_block1a55.port_b_data_width = 1;
defparam ram_block1a55.port_b_first_address = 0;
defparam ram_block1a55.port_b_first_bit_number = 55;
defparam ram_block1a55.port_b_last_address = 255;
defparam ram_block1a55.port_b_logical_ram_depth = 256;
defparam ram_block1a55.port_b_logical_ram_width = 144;
defparam ram_block1a55.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a55.port_b_read_enable_clock = "clock1";
defparam ram_block1a55.ram_block_type = "auto";

arriaii_ram_block ram_block1a87(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[87]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a87_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a87.clk0_core_clock_enable = "ena0";
defparam ram_block1a87.clk0_input_clock_enable = "ena2";
defparam ram_block1a87.clk1_core_clock_enable = "ena3";
defparam ram_block1a87.clk1_input_clock_enable = "ena3";
defparam ram_block1a87.clk1_output_clock_enable = "ena1";
defparam ram_block1a87.clock_duty_cycle_dependence = "on";
defparam ram_block1a87.data_interleave_offset_in_bits = 1;
defparam ram_block1a87.data_interleave_width_in_bits = 1;
defparam ram_block1a87.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a87.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a87.operation_mode = "dual_port";
defparam ram_block1a87.port_a_address_clear = "none";
defparam ram_block1a87.port_a_address_width = 8;
defparam ram_block1a87.port_a_data_out_clear = "none";
defparam ram_block1a87.port_a_data_out_clock = "none";
defparam ram_block1a87.port_a_data_width = 1;
defparam ram_block1a87.port_a_first_address = 0;
defparam ram_block1a87.port_a_first_bit_number = 87;
defparam ram_block1a87.port_a_last_address = 255;
defparam ram_block1a87.port_a_logical_ram_depth = 256;
defparam ram_block1a87.port_a_logical_ram_width = 144;
defparam ram_block1a87.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a87.port_b_address_clear = "none";
defparam ram_block1a87.port_b_address_clock = "clock1";
defparam ram_block1a87.port_b_address_width = 8;
defparam ram_block1a87.port_b_data_out_clear = "none";
defparam ram_block1a87.port_b_data_out_clock = "clock1";
defparam ram_block1a87.port_b_data_width = 1;
defparam ram_block1a87.port_b_first_address = 0;
defparam ram_block1a87.port_b_first_bit_number = 87;
defparam ram_block1a87.port_b_last_address = 255;
defparam ram_block1a87.port_b_logical_ram_depth = 256;
defparam ram_block1a87.port_b_logical_ram_width = 144;
defparam ram_block1a87.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a87.port_b_read_enable_clock = "clock1";
defparam ram_block1a87.ram_block_type = "auto";

arriaii_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena2";
defparam ram_block1a23.clk1_core_clock_enable = "ena3";
defparam ram_block1a23.clk1_input_clock_enable = "ena3";
defparam ram_block1a23.clk1_output_clock_enable = "ena1";
defparam ram_block1a23.clock_duty_cycle_dependence = "on";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 8;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 255;
defparam ram_block1a23.port_a_logical_ram_depth = 256;
defparam ram_block1a23.port_a_logical_ram_width = 144;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock1";
defparam ram_block1a23.port_b_address_width = 8;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "clock1";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 255;
defparam ram_block1a23.port_b_logical_ram_depth = 256;
defparam ram_block1a23.port_b_logical_ram_width = 144;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock1";
defparam ram_block1a23.ram_block_type = "auto";

arriaii_ram_block ram_block1a120(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[120]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a120_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a120.clk0_core_clock_enable = "ena0";
defparam ram_block1a120.clk0_input_clock_enable = "ena2";
defparam ram_block1a120.clk1_core_clock_enable = "ena3";
defparam ram_block1a120.clk1_input_clock_enable = "ena3";
defparam ram_block1a120.clk1_output_clock_enable = "ena1";
defparam ram_block1a120.clock_duty_cycle_dependence = "on";
defparam ram_block1a120.data_interleave_offset_in_bits = 1;
defparam ram_block1a120.data_interleave_width_in_bits = 1;
defparam ram_block1a120.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a120.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a120.operation_mode = "dual_port";
defparam ram_block1a120.port_a_address_clear = "none";
defparam ram_block1a120.port_a_address_width = 8;
defparam ram_block1a120.port_a_data_out_clear = "none";
defparam ram_block1a120.port_a_data_out_clock = "none";
defparam ram_block1a120.port_a_data_width = 1;
defparam ram_block1a120.port_a_first_address = 0;
defparam ram_block1a120.port_a_first_bit_number = 120;
defparam ram_block1a120.port_a_last_address = 255;
defparam ram_block1a120.port_a_logical_ram_depth = 256;
defparam ram_block1a120.port_a_logical_ram_width = 144;
defparam ram_block1a120.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a120.port_b_address_clear = "none";
defparam ram_block1a120.port_b_address_clock = "clock1";
defparam ram_block1a120.port_b_address_width = 8;
defparam ram_block1a120.port_b_data_out_clear = "none";
defparam ram_block1a120.port_b_data_out_clock = "clock1";
defparam ram_block1a120.port_b_data_width = 1;
defparam ram_block1a120.port_b_first_address = 0;
defparam ram_block1a120.port_b_first_bit_number = 120;
defparam ram_block1a120.port_b_last_address = 255;
defparam ram_block1a120.port_b_logical_ram_depth = 256;
defparam ram_block1a120.port_b_logical_ram_width = 144;
defparam ram_block1a120.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a120.port_b_read_enable_clock = "clock1";
defparam ram_block1a120.ram_block_type = "auto";

arriaii_ram_block ram_block1a56(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[56]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a56_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a56.clk0_core_clock_enable = "ena0";
defparam ram_block1a56.clk0_input_clock_enable = "ena2";
defparam ram_block1a56.clk1_core_clock_enable = "ena3";
defparam ram_block1a56.clk1_input_clock_enable = "ena3";
defparam ram_block1a56.clk1_output_clock_enable = "ena1";
defparam ram_block1a56.clock_duty_cycle_dependence = "on";
defparam ram_block1a56.data_interleave_offset_in_bits = 1;
defparam ram_block1a56.data_interleave_width_in_bits = 1;
defparam ram_block1a56.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a56.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a56.operation_mode = "dual_port";
defparam ram_block1a56.port_a_address_clear = "none";
defparam ram_block1a56.port_a_address_width = 8;
defparam ram_block1a56.port_a_data_out_clear = "none";
defparam ram_block1a56.port_a_data_out_clock = "none";
defparam ram_block1a56.port_a_data_width = 1;
defparam ram_block1a56.port_a_first_address = 0;
defparam ram_block1a56.port_a_first_bit_number = 56;
defparam ram_block1a56.port_a_last_address = 255;
defparam ram_block1a56.port_a_logical_ram_depth = 256;
defparam ram_block1a56.port_a_logical_ram_width = 144;
defparam ram_block1a56.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a56.port_b_address_clear = "none";
defparam ram_block1a56.port_b_address_clock = "clock1";
defparam ram_block1a56.port_b_address_width = 8;
defparam ram_block1a56.port_b_data_out_clear = "none";
defparam ram_block1a56.port_b_data_out_clock = "clock1";
defparam ram_block1a56.port_b_data_width = 1;
defparam ram_block1a56.port_b_first_address = 0;
defparam ram_block1a56.port_b_first_bit_number = 56;
defparam ram_block1a56.port_b_last_address = 255;
defparam ram_block1a56.port_b_logical_ram_depth = 256;
defparam ram_block1a56.port_b_logical_ram_width = 144;
defparam ram_block1a56.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a56.port_b_read_enable_clock = "clock1";
defparam ram_block1a56.ram_block_type = "auto";

arriaii_ram_block ram_block1a88(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[88]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a88_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a88.clk0_core_clock_enable = "ena0";
defparam ram_block1a88.clk0_input_clock_enable = "ena2";
defparam ram_block1a88.clk1_core_clock_enable = "ena3";
defparam ram_block1a88.clk1_input_clock_enable = "ena3";
defparam ram_block1a88.clk1_output_clock_enable = "ena1";
defparam ram_block1a88.clock_duty_cycle_dependence = "on";
defparam ram_block1a88.data_interleave_offset_in_bits = 1;
defparam ram_block1a88.data_interleave_width_in_bits = 1;
defparam ram_block1a88.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a88.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a88.operation_mode = "dual_port";
defparam ram_block1a88.port_a_address_clear = "none";
defparam ram_block1a88.port_a_address_width = 8;
defparam ram_block1a88.port_a_data_out_clear = "none";
defparam ram_block1a88.port_a_data_out_clock = "none";
defparam ram_block1a88.port_a_data_width = 1;
defparam ram_block1a88.port_a_first_address = 0;
defparam ram_block1a88.port_a_first_bit_number = 88;
defparam ram_block1a88.port_a_last_address = 255;
defparam ram_block1a88.port_a_logical_ram_depth = 256;
defparam ram_block1a88.port_a_logical_ram_width = 144;
defparam ram_block1a88.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a88.port_b_address_clear = "none";
defparam ram_block1a88.port_b_address_clock = "clock1";
defparam ram_block1a88.port_b_address_width = 8;
defparam ram_block1a88.port_b_data_out_clear = "none";
defparam ram_block1a88.port_b_data_out_clock = "clock1";
defparam ram_block1a88.port_b_data_width = 1;
defparam ram_block1a88.port_b_first_address = 0;
defparam ram_block1a88.port_b_first_bit_number = 88;
defparam ram_block1a88.port_b_last_address = 255;
defparam ram_block1a88.port_b_logical_ram_depth = 256;
defparam ram_block1a88.port_b_logical_ram_width = 144;
defparam ram_block1a88.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a88.port_b_read_enable_clock = "clock1";
defparam ram_block1a88.ram_block_type = "auto";

arriaii_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk0_input_clock_enable = "ena2";
defparam ram_block1a24.clk1_core_clock_enable = "ena3";
defparam ram_block1a24.clk1_input_clock_enable = "ena3";
defparam ram_block1a24.clk1_output_clock_enable = "ena1";
defparam ram_block1a24.clock_duty_cycle_dependence = "on";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 8;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 255;
defparam ram_block1a24.port_a_logical_ram_depth = 256;
defparam ram_block1a24.port_a_logical_ram_width = 144;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock1";
defparam ram_block1a24.port_b_address_width = 8;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "clock1";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 255;
defparam ram_block1a24.port_b_logical_ram_depth = 256;
defparam ram_block1a24.port_b_logical_ram_width = 144;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock1";
defparam ram_block1a24.ram_block_type = "auto";

arriaii_ram_block ram_block1a121(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[121]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a121_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a121.clk0_core_clock_enable = "ena0";
defparam ram_block1a121.clk0_input_clock_enable = "ena2";
defparam ram_block1a121.clk1_core_clock_enable = "ena3";
defparam ram_block1a121.clk1_input_clock_enable = "ena3";
defparam ram_block1a121.clk1_output_clock_enable = "ena1";
defparam ram_block1a121.clock_duty_cycle_dependence = "on";
defparam ram_block1a121.data_interleave_offset_in_bits = 1;
defparam ram_block1a121.data_interleave_width_in_bits = 1;
defparam ram_block1a121.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a121.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a121.operation_mode = "dual_port";
defparam ram_block1a121.port_a_address_clear = "none";
defparam ram_block1a121.port_a_address_width = 8;
defparam ram_block1a121.port_a_data_out_clear = "none";
defparam ram_block1a121.port_a_data_out_clock = "none";
defparam ram_block1a121.port_a_data_width = 1;
defparam ram_block1a121.port_a_first_address = 0;
defparam ram_block1a121.port_a_first_bit_number = 121;
defparam ram_block1a121.port_a_last_address = 255;
defparam ram_block1a121.port_a_logical_ram_depth = 256;
defparam ram_block1a121.port_a_logical_ram_width = 144;
defparam ram_block1a121.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a121.port_b_address_clear = "none";
defparam ram_block1a121.port_b_address_clock = "clock1";
defparam ram_block1a121.port_b_address_width = 8;
defparam ram_block1a121.port_b_data_out_clear = "none";
defparam ram_block1a121.port_b_data_out_clock = "clock1";
defparam ram_block1a121.port_b_data_width = 1;
defparam ram_block1a121.port_b_first_address = 0;
defparam ram_block1a121.port_b_first_bit_number = 121;
defparam ram_block1a121.port_b_last_address = 255;
defparam ram_block1a121.port_b_logical_ram_depth = 256;
defparam ram_block1a121.port_b_logical_ram_width = 144;
defparam ram_block1a121.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a121.port_b_read_enable_clock = "clock1";
defparam ram_block1a121.ram_block_type = "auto";

arriaii_ram_block ram_block1a57(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[57]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a57_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a57.clk0_core_clock_enable = "ena0";
defparam ram_block1a57.clk0_input_clock_enable = "ena2";
defparam ram_block1a57.clk1_core_clock_enable = "ena3";
defparam ram_block1a57.clk1_input_clock_enable = "ena3";
defparam ram_block1a57.clk1_output_clock_enable = "ena1";
defparam ram_block1a57.clock_duty_cycle_dependence = "on";
defparam ram_block1a57.data_interleave_offset_in_bits = 1;
defparam ram_block1a57.data_interleave_width_in_bits = 1;
defparam ram_block1a57.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a57.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a57.operation_mode = "dual_port";
defparam ram_block1a57.port_a_address_clear = "none";
defparam ram_block1a57.port_a_address_width = 8;
defparam ram_block1a57.port_a_data_out_clear = "none";
defparam ram_block1a57.port_a_data_out_clock = "none";
defparam ram_block1a57.port_a_data_width = 1;
defparam ram_block1a57.port_a_first_address = 0;
defparam ram_block1a57.port_a_first_bit_number = 57;
defparam ram_block1a57.port_a_last_address = 255;
defparam ram_block1a57.port_a_logical_ram_depth = 256;
defparam ram_block1a57.port_a_logical_ram_width = 144;
defparam ram_block1a57.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a57.port_b_address_clear = "none";
defparam ram_block1a57.port_b_address_clock = "clock1";
defparam ram_block1a57.port_b_address_width = 8;
defparam ram_block1a57.port_b_data_out_clear = "none";
defparam ram_block1a57.port_b_data_out_clock = "clock1";
defparam ram_block1a57.port_b_data_width = 1;
defparam ram_block1a57.port_b_first_address = 0;
defparam ram_block1a57.port_b_first_bit_number = 57;
defparam ram_block1a57.port_b_last_address = 255;
defparam ram_block1a57.port_b_logical_ram_depth = 256;
defparam ram_block1a57.port_b_logical_ram_width = 144;
defparam ram_block1a57.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a57.port_b_read_enable_clock = "clock1";
defparam ram_block1a57.ram_block_type = "auto";

arriaii_ram_block ram_block1a89(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[89]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a89_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a89.clk0_core_clock_enable = "ena0";
defparam ram_block1a89.clk0_input_clock_enable = "ena2";
defparam ram_block1a89.clk1_core_clock_enable = "ena3";
defparam ram_block1a89.clk1_input_clock_enable = "ena3";
defparam ram_block1a89.clk1_output_clock_enable = "ena1";
defparam ram_block1a89.clock_duty_cycle_dependence = "on";
defparam ram_block1a89.data_interleave_offset_in_bits = 1;
defparam ram_block1a89.data_interleave_width_in_bits = 1;
defparam ram_block1a89.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a89.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a89.operation_mode = "dual_port";
defparam ram_block1a89.port_a_address_clear = "none";
defparam ram_block1a89.port_a_address_width = 8;
defparam ram_block1a89.port_a_data_out_clear = "none";
defparam ram_block1a89.port_a_data_out_clock = "none";
defparam ram_block1a89.port_a_data_width = 1;
defparam ram_block1a89.port_a_first_address = 0;
defparam ram_block1a89.port_a_first_bit_number = 89;
defparam ram_block1a89.port_a_last_address = 255;
defparam ram_block1a89.port_a_logical_ram_depth = 256;
defparam ram_block1a89.port_a_logical_ram_width = 144;
defparam ram_block1a89.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a89.port_b_address_clear = "none";
defparam ram_block1a89.port_b_address_clock = "clock1";
defparam ram_block1a89.port_b_address_width = 8;
defparam ram_block1a89.port_b_data_out_clear = "none";
defparam ram_block1a89.port_b_data_out_clock = "clock1";
defparam ram_block1a89.port_b_data_width = 1;
defparam ram_block1a89.port_b_first_address = 0;
defparam ram_block1a89.port_b_first_bit_number = 89;
defparam ram_block1a89.port_b_last_address = 255;
defparam ram_block1a89.port_b_logical_ram_depth = 256;
defparam ram_block1a89.port_b_logical_ram_width = 144;
defparam ram_block1a89.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a89.port_b_read_enable_clock = "clock1";
defparam ram_block1a89.ram_block_type = "auto";

arriaii_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk0_input_clock_enable = "ena2";
defparam ram_block1a25.clk1_core_clock_enable = "ena3";
defparam ram_block1a25.clk1_input_clock_enable = "ena3";
defparam ram_block1a25.clk1_output_clock_enable = "ena1";
defparam ram_block1a25.clock_duty_cycle_dependence = "on";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 8;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 255;
defparam ram_block1a25.port_a_logical_ram_depth = 256;
defparam ram_block1a25.port_a_logical_ram_width = 144;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock1";
defparam ram_block1a25.port_b_address_width = 8;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "clock1";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 255;
defparam ram_block1a25.port_b_logical_ram_depth = 256;
defparam ram_block1a25.port_b_logical_ram_width = 144;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock1";
defparam ram_block1a25.ram_block_type = "auto";

arriaii_ram_block ram_block1a122(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[122]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a122_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a122.clk0_core_clock_enable = "ena0";
defparam ram_block1a122.clk0_input_clock_enable = "ena2";
defparam ram_block1a122.clk1_core_clock_enable = "ena3";
defparam ram_block1a122.clk1_input_clock_enable = "ena3";
defparam ram_block1a122.clk1_output_clock_enable = "ena1";
defparam ram_block1a122.clock_duty_cycle_dependence = "on";
defparam ram_block1a122.data_interleave_offset_in_bits = 1;
defparam ram_block1a122.data_interleave_width_in_bits = 1;
defparam ram_block1a122.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a122.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a122.operation_mode = "dual_port";
defparam ram_block1a122.port_a_address_clear = "none";
defparam ram_block1a122.port_a_address_width = 8;
defparam ram_block1a122.port_a_data_out_clear = "none";
defparam ram_block1a122.port_a_data_out_clock = "none";
defparam ram_block1a122.port_a_data_width = 1;
defparam ram_block1a122.port_a_first_address = 0;
defparam ram_block1a122.port_a_first_bit_number = 122;
defparam ram_block1a122.port_a_last_address = 255;
defparam ram_block1a122.port_a_logical_ram_depth = 256;
defparam ram_block1a122.port_a_logical_ram_width = 144;
defparam ram_block1a122.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a122.port_b_address_clear = "none";
defparam ram_block1a122.port_b_address_clock = "clock1";
defparam ram_block1a122.port_b_address_width = 8;
defparam ram_block1a122.port_b_data_out_clear = "none";
defparam ram_block1a122.port_b_data_out_clock = "clock1";
defparam ram_block1a122.port_b_data_width = 1;
defparam ram_block1a122.port_b_first_address = 0;
defparam ram_block1a122.port_b_first_bit_number = 122;
defparam ram_block1a122.port_b_last_address = 255;
defparam ram_block1a122.port_b_logical_ram_depth = 256;
defparam ram_block1a122.port_b_logical_ram_width = 144;
defparam ram_block1a122.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a122.port_b_read_enable_clock = "clock1";
defparam ram_block1a122.ram_block_type = "auto";

arriaii_ram_block ram_block1a58(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[58]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a58_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a58.clk0_core_clock_enable = "ena0";
defparam ram_block1a58.clk0_input_clock_enable = "ena2";
defparam ram_block1a58.clk1_core_clock_enable = "ena3";
defparam ram_block1a58.clk1_input_clock_enable = "ena3";
defparam ram_block1a58.clk1_output_clock_enable = "ena1";
defparam ram_block1a58.clock_duty_cycle_dependence = "on";
defparam ram_block1a58.data_interleave_offset_in_bits = 1;
defparam ram_block1a58.data_interleave_width_in_bits = 1;
defparam ram_block1a58.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a58.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a58.operation_mode = "dual_port";
defparam ram_block1a58.port_a_address_clear = "none";
defparam ram_block1a58.port_a_address_width = 8;
defparam ram_block1a58.port_a_data_out_clear = "none";
defparam ram_block1a58.port_a_data_out_clock = "none";
defparam ram_block1a58.port_a_data_width = 1;
defparam ram_block1a58.port_a_first_address = 0;
defparam ram_block1a58.port_a_first_bit_number = 58;
defparam ram_block1a58.port_a_last_address = 255;
defparam ram_block1a58.port_a_logical_ram_depth = 256;
defparam ram_block1a58.port_a_logical_ram_width = 144;
defparam ram_block1a58.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a58.port_b_address_clear = "none";
defparam ram_block1a58.port_b_address_clock = "clock1";
defparam ram_block1a58.port_b_address_width = 8;
defparam ram_block1a58.port_b_data_out_clear = "none";
defparam ram_block1a58.port_b_data_out_clock = "clock1";
defparam ram_block1a58.port_b_data_width = 1;
defparam ram_block1a58.port_b_first_address = 0;
defparam ram_block1a58.port_b_first_bit_number = 58;
defparam ram_block1a58.port_b_last_address = 255;
defparam ram_block1a58.port_b_logical_ram_depth = 256;
defparam ram_block1a58.port_b_logical_ram_width = 144;
defparam ram_block1a58.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a58.port_b_read_enable_clock = "clock1";
defparam ram_block1a58.ram_block_type = "auto";

arriaii_ram_block ram_block1a90(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[90]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a90_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a90.clk0_core_clock_enable = "ena0";
defparam ram_block1a90.clk0_input_clock_enable = "ena2";
defparam ram_block1a90.clk1_core_clock_enable = "ena3";
defparam ram_block1a90.clk1_input_clock_enable = "ena3";
defparam ram_block1a90.clk1_output_clock_enable = "ena1";
defparam ram_block1a90.clock_duty_cycle_dependence = "on";
defparam ram_block1a90.data_interleave_offset_in_bits = 1;
defparam ram_block1a90.data_interleave_width_in_bits = 1;
defparam ram_block1a90.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a90.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a90.operation_mode = "dual_port";
defparam ram_block1a90.port_a_address_clear = "none";
defparam ram_block1a90.port_a_address_width = 8;
defparam ram_block1a90.port_a_data_out_clear = "none";
defparam ram_block1a90.port_a_data_out_clock = "none";
defparam ram_block1a90.port_a_data_width = 1;
defparam ram_block1a90.port_a_first_address = 0;
defparam ram_block1a90.port_a_first_bit_number = 90;
defparam ram_block1a90.port_a_last_address = 255;
defparam ram_block1a90.port_a_logical_ram_depth = 256;
defparam ram_block1a90.port_a_logical_ram_width = 144;
defparam ram_block1a90.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a90.port_b_address_clear = "none";
defparam ram_block1a90.port_b_address_clock = "clock1";
defparam ram_block1a90.port_b_address_width = 8;
defparam ram_block1a90.port_b_data_out_clear = "none";
defparam ram_block1a90.port_b_data_out_clock = "clock1";
defparam ram_block1a90.port_b_data_width = 1;
defparam ram_block1a90.port_b_first_address = 0;
defparam ram_block1a90.port_b_first_bit_number = 90;
defparam ram_block1a90.port_b_last_address = 255;
defparam ram_block1a90.port_b_logical_ram_depth = 256;
defparam ram_block1a90.port_b_logical_ram_width = 144;
defparam ram_block1a90.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a90.port_b_read_enable_clock = "clock1";
defparam ram_block1a90.ram_block_type = "auto";

arriaii_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk0_input_clock_enable = "ena2";
defparam ram_block1a26.clk1_core_clock_enable = "ena3";
defparam ram_block1a26.clk1_input_clock_enable = "ena3";
defparam ram_block1a26.clk1_output_clock_enable = "ena1";
defparam ram_block1a26.clock_duty_cycle_dependence = "on";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 8;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 255;
defparam ram_block1a26.port_a_logical_ram_depth = 256;
defparam ram_block1a26.port_a_logical_ram_width = 144;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock1";
defparam ram_block1a26.port_b_address_width = 8;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "clock1";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 255;
defparam ram_block1a26.port_b_logical_ram_depth = 256;
defparam ram_block1a26.port_b_logical_ram_width = 144;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock1";
defparam ram_block1a26.ram_block_type = "auto";

arriaii_ram_block ram_block1a123(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[123]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a123_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a123.clk0_core_clock_enable = "ena0";
defparam ram_block1a123.clk0_input_clock_enable = "ena2";
defparam ram_block1a123.clk1_core_clock_enable = "ena3";
defparam ram_block1a123.clk1_input_clock_enable = "ena3";
defparam ram_block1a123.clk1_output_clock_enable = "ena1";
defparam ram_block1a123.clock_duty_cycle_dependence = "on";
defparam ram_block1a123.data_interleave_offset_in_bits = 1;
defparam ram_block1a123.data_interleave_width_in_bits = 1;
defparam ram_block1a123.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a123.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a123.operation_mode = "dual_port";
defparam ram_block1a123.port_a_address_clear = "none";
defparam ram_block1a123.port_a_address_width = 8;
defparam ram_block1a123.port_a_data_out_clear = "none";
defparam ram_block1a123.port_a_data_out_clock = "none";
defparam ram_block1a123.port_a_data_width = 1;
defparam ram_block1a123.port_a_first_address = 0;
defparam ram_block1a123.port_a_first_bit_number = 123;
defparam ram_block1a123.port_a_last_address = 255;
defparam ram_block1a123.port_a_logical_ram_depth = 256;
defparam ram_block1a123.port_a_logical_ram_width = 144;
defparam ram_block1a123.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a123.port_b_address_clear = "none";
defparam ram_block1a123.port_b_address_clock = "clock1";
defparam ram_block1a123.port_b_address_width = 8;
defparam ram_block1a123.port_b_data_out_clear = "none";
defparam ram_block1a123.port_b_data_out_clock = "clock1";
defparam ram_block1a123.port_b_data_width = 1;
defparam ram_block1a123.port_b_first_address = 0;
defparam ram_block1a123.port_b_first_bit_number = 123;
defparam ram_block1a123.port_b_last_address = 255;
defparam ram_block1a123.port_b_logical_ram_depth = 256;
defparam ram_block1a123.port_b_logical_ram_width = 144;
defparam ram_block1a123.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a123.port_b_read_enable_clock = "clock1";
defparam ram_block1a123.ram_block_type = "auto";

arriaii_ram_block ram_block1a59(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[59]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a59_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a59.clk0_core_clock_enable = "ena0";
defparam ram_block1a59.clk0_input_clock_enable = "ena2";
defparam ram_block1a59.clk1_core_clock_enable = "ena3";
defparam ram_block1a59.clk1_input_clock_enable = "ena3";
defparam ram_block1a59.clk1_output_clock_enable = "ena1";
defparam ram_block1a59.clock_duty_cycle_dependence = "on";
defparam ram_block1a59.data_interleave_offset_in_bits = 1;
defparam ram_block1a59.data_interleave_width_in_bits = 1;
defparam ram_block1a59.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a59.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a59.operation_mode = "dual_port";
defparam ram_block1a59.port_a_address_clear = "none";
defparam ram_block1a59.port_a_address_width = 8;
defparam ram_block1a59.port_a_data_out_clear = "none";
defparam ram_block1a59.port_a_data_out_clock = "none";
defparam ram_block1a59.port_a_data_width = 1;
defparam ram_block1a59.port_a_first_address = 0;
defparam ram_block1a59.port_a_first_bit_number = 59;
defparam ram_block1a59.port_a_last_address = 255;
defparam ram_block1a59.port_a_logical_ram_depth = 256;
defparam ram_block1a59.port_a_logical_ram_width = 144;
defparam ram_block1a59.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a59.port_b_address_clear = "none";
defparam ram_block1a59.port_b_address_clock = "clock1";
defparam ram_block1a59.port_b_address_width = 8;
defparam ram_block1a59.port_b_data_out_clear = "none";
defparam ram_block1a59.port_b_data_out_clock = "clock1";
defparam ram_block1a59.port_b_data_width = 1;
defparam ram_block1a59.port_b_first_address = 0;
defparam ram_block1a59.port_b_first_bit_number = 59;
defparam ram_block1a59.port_b_last_address = 255;
defparam ram_block1a59.port_b_logical_ram_depth = 256;
defparam ram_block1a59.port_b_logical_ram_width = 144;
defparam ram_block1a59.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a59.port_b_read_enable_clock = "clock1";
defparam ram_block1a59.ram_block_type = "auto";

arriaii_ram_block ram_block1a91(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[91]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a91_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a91.clk0_core_clock_enable = "ena0";
defparam ram_block1a91.clk0_input_clock_enable = "ena2";
defparam ram_block1a91.clk1_core_clock_enable = "ena3";
defparam ram_block1a91.clk1_input_clock_enable = "ena3";
defparam ram_block1a91.clk1_output_clock_enable = "ena1";
defparam ram_block1a91.clock_duty_cycle_dependence = "on";
defparam ram_block1a91.data_interleave_offset_in_bits = 1;
defparam ram_block1a91.data_interleave_width_in_bits = 1;
defparam ram_block1a91.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a91.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a91.operation_mode = "dual_port";
defparam ram_block1a91.port_a_address_clear = "none";
defparam ram_block1a91.port_a_address_width = 8;
defparam ram_block1a91.port_a_data_out_clear = "none";
defparam ram_block1a91.port_a_data_out_clock = "none";
defparam ram_block1a91.port_a_data_width = 1;
defparam ram_block1a91.port_a_first_address = 0;
defparam ram_block1a91.port_a_first_bit_number = 91;
defparam ram_block1a91.port_a_last_address = 255;
defparam ram_block1a91.port_a_logical_ram_depth = 256;
defparam ram_block1a91.port_a_logical_ram_width = 144;
defparam ram_block1a91.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a91.port_b_address_clear = "none";
defparam ram_block1a91.port_b_address_clock = "clock1";
defparam ram_block1a91.port_b_address_width = 8;
defparam ram_block1a91.port_b_data_out_clear = "none";
defparam ram_block1a91.port_b_data_out_clock = "clock1";
defparam ram_block1a91.port_b_data_width = 1;
defparam ram_block1a91.port_b_first_address = 0;
defparam ram_block1a91.port_b_first_bit_number = 91;
defparam ram_block1a91.port_b_last_address = 255;
defparam ram_block1a91.port_b_logical_ram_depth = 256;
defparam ram_block1a91.port_b_logical_ram_width = 144;
defparam ram_block1a91.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a91.port_b_read_enable_clock = "clock1";
defparam ram_block1a91.ram_block_type = "auto";

arriaii_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk0_input_clock_enable = "ena2";
defparam ram_block1a27.clk1_core_clock_enable = "ena3";
defparam ram_block1a27.clk1_input_clock_enable = "ena3";
defparam ram_block1a27.clk1_output_clock_enable = "ena1";
defparam ram_block1a27.clock_duty_cycle_dependence = "on";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 8;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 255;
defparam ram_block1a27.port_a_logical_ram_depth = 256;
defparam ram_block1a27.port_a_logical_ram_width = 144;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock1";
defparam ram_block1a27.port_b_address_width = 8;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "clock1";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 255;
defparam ram_block1a27.port_b_logical_ram_depth = 256;
defparam ram_block1a27.port_b_logical_ram_width = 144;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock1";
defparam ram_block1a27.ram_block_type = "auto";

arriaii_ram_block ram_block1a124(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[124]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a124_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a124.clk0_core_clock_enable = "ena0";
defparam ram_block1a124.clk0_input_clock_enable = "ena2";
defparam ram_block1a124.clk1_core_clock_enable = "ena3";
defparam ram_block1a124.clk1_input_clock_enable = "ena3";
defparam ram_block1a124.clk1_output_clock_enable = "ena1";
defparam ram_block1a124.clock_duty_cycle_dependence = "on";
defparam ram_block1a124.data_interleave_offset_in_bits = 1;
defparam ram_block1a124.data_interleave_width_in_bits = 1;
defparam ram_block1a124.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a124.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a124.operation_mode = "dual_port";
defparam ram_block1a124.port_a_address_clear = "none";
defparam ram_block1a124.port_a_address_width = 8;
defparam ram_block1a124.port_a_data_out_clear = "none";
defparam ram_block1a124.port_a_data_out_clock = "none";
defparam ram_block1a124.port_a_data_width = 1;
defparam ram_block1a124.port_a_first_address = 0;
defparam ram_block1a124.port_a_first_bit_number = 124;
defparam ram_block1a124.port_a_last_address = 255;
defparam ram_block1a124.port_a_logical_ram_depth = 256;
defparam ram_block1a124.port_a_logical_ram_width = 144;
defparam ram_block1a124.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a124.port_b_address_clear = "none";
defparam ram_block1a124.port_b_address_clock = "clock1";
defparam ram_block1a124.port_b_address_width = 8;
defparam ram_block1a124.port_b_data_out_clear = "none";
defparam ram_block1a124.port_b_data_out_clock = "clock1";
defparam ram_block1a124.port_b_data_width = 1;
defparam ram_block1a124.port_b_first_address = 0;
defparam ram_block1a124.port_b_first_bit_number = 124;
defparam ram_block1a124.port_b_last_address = 255;
defparam ram_block1a124.port_b_logical_ram_depth = 256;
defparam ram_block1a124.port_b_logical_ram_width = 144;
defparam ram_block1a124.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a124.port_b_read_enable_clock = "clock1";
defparam ram_block1a124.ram_block_type = "auto";

arriaii_ram_block ram_block1a60(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[60]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a60_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a60.clk0_core_clock_enable = "ena0";
defparam ram_block1a60.clk0_input_clock_enable = "ena2";
defparam ram_block1a60.clk1_core_clock_enable = "ena3";
defparam ram_block1a60.clk1_input_clock_enable = "ena3";
defparam ram_block1a60.clk1_output_clock_enable = "ena1";
defparam ram_block1a60.clock_duty_cycle_dependence = "on";
defparam ram_block1a60.data_interleave_offset_in_bits = 1;
defparam ram_block1a60.data_interleave_width_in_bits = 1;
defparam ram_block1a60.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a60.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a60.operation_mode = "dual_port";
defparam ram_block1a60.port_a_address_clear = "none";
defparam ram_block1a60.port_a_address_width = 8;
defparam ram_block1a60.port_a_data_out_clear = "none";
defparam ram_block1a60.port_a_data_out_clock = "none";
defparam ram_block1a60.port_a_data_width = 1;
defparam ram_block1a60.port_a_first_address = 0;
defparam ram_block1a60.port_a_first_bit_number = 60;
defparam ram_block1a60.port_a_last_address = 255;
defparam ram_block1a60.port_a_logical_ram_depth = 256;
defparam ram_block1a60.port_a_logical_ram_width = 144;
defparam ram_block1a60.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a60.port_b_address_clear = "none";
defparam ram_block1a60.port_b_address_clock = "clock1";
defparam ram_block1a60.port_b_address_width = 8;
defparam ram_block1a60.port_b_data_out_clear = "none";
defparam ram_block1a60.port_b_data_out_clock = "clock1";
defparam ram_block1a60.port_b_data_width = 1;
defparam ram_block1a60.port_b_first_address = 0;
defparam ram_block1a60.port_b_first_bit_number = 60;
defparam ram_block1a60.port_b_last_address = 255;
defparam ram_block1a60.port_b_logical_ram_depth = 256;
defparam ram_block1a60.port_b_logical_ram_width = 144;
defparam ram_block1a60.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a60.port_b_read_enable_clock = "clock1";
defparam ram_block1a60.ram_block_type = "auto";

arriaii_ram_block ram_block1a92(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[92]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a92_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a92.clk0_core_clock_enable = "ena0";
defparam ram_block1a92.clk0_input_clock_enable = "ena2";
defparam ram_block1a92.clk1_core_clock_enable = "ena3";
defparam ram_block1a92.clk1_input_clock_enable = "ena3";
defparam ram_block1a92.clk1_output_clock_enable = "ena1";
defparam ram_block1a92.clock_duty_cycle_dependence = "on";
defparam ram_block1a92.data_interleave_offset_in_bits = 1;
defparam ram_block1a92.data_interleave_width_in_bits = 1;
defparam ram_block1a92.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a92.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a92.operation_mode = "dual_port";
defparam ram_block1a92.port_a_address_clear = "none";
defparam ram_block1a92.port_a_address_width = 8;
defparam ram_block1a92.port_a_data_out_clear = "none";
defparam ram_block1a92.port_a_data_out_clock = "none";
defparam ram_block1a92.port_a_data_width = 1;
defparam ram_block1a92.port_a_first_address = 0;
defparam ram_block1a92.port_a_first_bit_number = 92;
defparam ram_block1a92.port_a_last_address = 255;
defparam ram_block1a92.port_a_logical_ram_depth = 256;
defparam ram_block1a92.port_a_logical_ram_width = 144;
defparam ram_block1a92.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a92.port_b_address_clear = "none";
defparam ram_block1a92.port_b_address_clock = "clock1";
defparam ram_block1a92.port_b_address_width = 8;
defparam ram_block1a92.port_b_data_out_clear = "none";
defparam ram_block1a92.port_b_data_out_clock = "clock1";
defparam ram_block1a92.port_b_data_width = 1;
defparam ram_block1a92.port_b_first_address = 0;
defparam ram_block1a92.port_b_first_bit_number = 92;
defparam ram_block1a92.port_b_last_address = 255;
defparam ram_block1a92.port_b_logical_ram_depth = 256;
defparam ram_block1a92.port_b_logical_ram_width = 144;
defparam ram_block1a92.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a92.port_b_read_enable_clock = "clock1";
defparam ram_block1a92.ram_block_type = "auto";

arriaii_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk0_input_clock_enable = "ena2";
defparam ram_block1a28.clk1_core_clock_enable = "ena3";
defparam ram_block1a28.clk1_input_clock_enable = "ena3";
defparam ram_block1a28.clk1_output_clock_enable = "ena1";
defparam ram_block1a28.clock_duty_cycle_dependence = "on";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 8;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 255;
defparam ram_block1a28.port_a_logical_ram_depth = 256;
defparam ram_block1a28.port_a_logical_ram_width = 144;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock1";
defparam ram_block1a28.port_b_address_width = 8;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "clock1";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 255;
defparam ram_block1a28.port_b_logical_ram_depth = 256;
defparam ram_block1a28.port_b_logical_ram_width = 144;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock1";
defparam ram_block1a28.ram_block_type = "auto";

arriaii_ram_block ram_block1a125(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[125]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a125_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a125.clk0_core_clock_enable = "ena0";
defparam ram_block1a125.clk0_input_clock_enable = "ena2";
defparam ram_block1a125.clk1_core_clock_enable = "ena3";
defparam ram_block1a125.clk1_input_clock_enable = "ena3";
defparam ram_block1a125.clk1_output_clock_enable = "ena1";
defparam ram_block1a125.clock_duty_cycle_dependence = "on";
defparam ram_block1a125.data_interleave_offset_in_bits = 1;
defparam ram_block1a125.data_interleave_width_in_bits = 1;
defparam ram_block1a125.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a125.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a125.operation_mode = "dual_port";
defparam ram_block1a125.port_a_address_clear = "none";
defparam ram_block1a125.port_a_address_width = 8;
defparam ram_block1a125.port_a_data_out_clear = "none";
defparam ram_block1a125.port_a_data_out_clock = "none";
defparam ram_block1a125.port_a_data_width = 1;
defparam ram_block1a125.port_a_first_address = 0;
defparam ram_block1a125.port_a_first_bit_number = 125;
defparam ram_block1a125.port_a_last_address = 255;
defparam ram_block1a125.port_a_logical_ram_depth = 256;
defparam ram_block1a125.port_a_logical_ram_width = 144;
defparam ram_block1a125.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a125.port_b_address_clear = "none";
defparam ram_block1a125.port_b_address_clock = "clock1";
defparam ram_block1a125.port_b_address_width = 8;
defparam ram_block1a125.port_b_data_out_clear = "none";
defparam ram_block1a125.port_b_data_out_clock = "clock1";
defparam ram_block1a125.port_b_data_width = 1;
defparam ram_block1a125.port_b_first_address = 0;
defparam ram_block1a125.port_b_first_bit_number = 125;
defparam ram_block1a125.port_b_last_address = 255;
defparam ram_block1a125.port_b_logical_ram_depth = 256;
defparam ram_block1a125.port_b_logical_ram_width = 144;
defparam ram_block1a125.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a125.port_b_read_enable_clock = "clock1";
defparam ram_block1a125.ram_block_type = "auto";

arriaii_ram_block ram_block1a61(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[61]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a61_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a61.clk0_core_clock_enable = "ena0";
defparam ram_block1a61.clk0_input_clock_enable = "ena2";
defparam ram_block1a61.clk1_core_clock_enable = "ena3";
defparam ram_block1a61.clk1_input_clock_enable = "ena3";
defparam ram_block1a61.clk1_output_clock_enable = "ena1";
defparam ram_block1a61.clock_duty_cycle_dependence = "on";
defparam ram_block1a61.data_interleave_offset_in_bits = 1;
defparam ram_block1a61.data_interleave_width_in_bits = 1;
defparam ram_block1a61.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a61.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a61.operation_mode = "dual_port";
defparam ram_block1a61.port_a_address_clear = "none";
defparam ram_block1a61.port_a_address_width = 8;
defparam ram_block1a61.port_a_data_out_clear = "none";
defparam ram_block1a61.port_a_data_out_clock = "none";
defparam ram_block1a61.port_a_data_width = 1;
defparam ram_block1a61.port_a_first_address = 0;
defparam ram_block1a61.port_a_first_bit_number = 61;
defparam ram_block1a61.port_a_last_address = 255;
defparam ram_block1a61.port_a_logical_ram_depth = 256;
defparam ram_block1a61.port_a_logical_ram_width = 144;
defparam ram_block1a61.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a61.port_b_address_clear = "none";
defparam ram_block1a61.port_b_address_clock = "clock1";
defparam ram_block1a61.port_b_address_width = 8;
defparam ram_block1a61.port_b_data_out_clear = "none";
defparam ram_block1a61.port_b_data_out_clock = "clock1";
defparam ram_block1a61.port_b_data_width = 1;
defparam ram_block1a61.port_b_first_address = 0;
defparam ram_block1a61.port_b_first_bit_number = 61;
defparam ram_block1a61.port_b_last_address = 255;
defparam ram_block1a61.port_b_logical_ram_depth = 256;
defparam ram_block1a61.port_b_logical_ram_width = 144;
defparam ram_block1a61.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a61.port_b_read_enable_clock = "clock1";
defparam ram_block1a61.ram_block_type = "auto";

arriaii_ram_block ram_block1a93(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[93]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a93_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a93.clk0_core_clock_enable = "ena0";
defparam ram_block1a93.clk0_input_clock_enable = "ena2";
defparam ram_block1a93.clk1_core_clock_enable = "ena3";
defparam ram_block1a93.clk1_input_clock_enable = "ena3";
defparam ram_block1a93.clk1_output_clock_enable = "ena1";
defparam ram_block1a93.clock_duty_cycle_dependence = "on";
defparam ram_block1a93.data_interleave_offset_in_bits = 1;
defparam ram_block1a93.data_interleave_width_in_bits = 1;
defparam ram_block1a93.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a93.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a93.operation_mode = "dual_port";
defparam ram_block1a93.port_a_address_clear = "none";
defparam ram_block1a93.port_a_address_width = 8;
defparam ram_block1a93.port_a_data_out_clear = "none";
defparam ram_block1a93.port_a_data_out_clock = "none";
defparam ram_block1a93.port_a_data_width = 1;
defparam ram_block1a93.port_a_first_address = 0;
defparam ram_block1a93.port_a_first_bit_number = 93;
defparam ram_block1a93.port_a_last_address = 255;
defparam ram_block1a93.port_a_logical_ram_depth = 256;
defparam ram_block1a93.port_a_logical_ram_width = 144;
defparam ram_block1a93.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a93.port_b_address_clear = "none";
defparam ram_block1a93.port_b_address_clock = "clock1";
defparam ram_block1a93.port_b_address_width = 8;
defparam ram_block1a93.port_b_data_out_clear = "none";
defparam ram_block1a93.port_b_data_out_clock = "clock1";
defparam ram_block1a93.port_b_data_width = 1;
defparam ram_block1a93.port_b_first_address = 0;
defparam ram_block1a93.port_b_first_bit_number = 93;
defparam ram_block1a93.port_b_last_address = 255;
defparam ram_block1a93.port_b_logical_ram_depth = 256;
defparam ram_block1a93.port_b_logical_ram_width = 144;
defparam ram_block1a93.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a93.port_b_read_enable_clock = "clock1";
defparam ram_block1a93.ram_block_type = "auto";

arriaii_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk0_input_clock_enable = "ena2";
defparam ram_block1a29.clk1_core_clock_enable = "ena3";
defparam ram_block1a29.clk1_input_clock_enable = "ena3";
defparam ram_block1a29.clk1_output_clock_enable = "ena1";
defparam ram_block1a29.clock_duty_cycle_dependence = "on";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 8;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 255;
defparam ram_block1a29.port_a_logical_ram_depth = 256;
defparam ram_block1a29.port_a_logical_ram_width = 144;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock1";
defparam ram_block1a29.port_b_address_width = 8;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "clock1";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 255;
defparam ram_block1a29.port_b_logical_ram_depth = 256;
defparam ram_block1a29.port_b_logical_ram_width = 144;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock1";
defparam ram_block1a29.ram_block_type = "auto";

arriaii_ram_block ram_block1a126(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[126]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a126_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a126.clk0_core_clock_enable = "ena0";
defparam ram_block1a126.clk0_input_clock_enable = "ena2";
defparam ram_block1a126.clk1_core_clock_enable = "ena3";
defparam ram_block1a126.clk1_input_clock_enable = "ena3";
defparam ram_block1a126.clk1_output_clock_enable = "ena1";
defparam ram_block1a126.clock_duty_cycle_dependence = "on";
defparam ram_block1a126.data_interleave_offset_in_bits = 1;
defparam ram_block1a126.data_interleave_width_in_bits = 1;
defparam ram_block1a126.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a126.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a126.operation_mode = "dual_port";
defparam ram_block1a126.port_a_address_clear = "none";
defparam ram_block1a126.port_a_address_width = 8;
defparam ram_block1a126.port_a_data_out_clear = "none";
defparam ram_block1a126.port_a_data_out_clock = "none";
defparam ram_block1a126.port_a_data_width = 1;
defparam ram_block1a126.port_a_first_address = 0;
defparam ram_block1a126.port_a_first_bit_number = 126;
defparam ram_block1a126.port_a_last_address = 255;
defparam ram_block1a126.port_a_logical_ram_depth = 256;
defparam ram_block1a126.port_a_logical_ram_width = 144;
defparam ram_block1a126.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a126.port_b_address_clear = "none";
defparam ram_block1a126.port_b_address_clock = "clock1";
defparam ram_block1a126.port_b_address_width = 8;
defparam ram_block1a126.port_b_data_out_clear = "none";
defparam ram_block1a126.port_b_data_out_clock = "clock1";
defparam ram_block1a126.port_b_data_width = 1;
defparam ram_block1a126.port_b_first_address = 0;
defparam ram_block1a126.port_b_first_bit_number = 126;
defparam ram_block1a126.port_b_last_address = 255;
defparam ram_block1a126.port_b_logical_ram_depth = 256;
defparam ram_block1a126.port_b_logical_ram_width = 144;
defparam ram_block1a126.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a126.port_b_read_enable_clock = "clock1";
defparam ram_block1a126.ram_block_type = "auto";

arriaii_ram_block ram_block1a62(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[62]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a62_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a62.clk0_core_clock_enable = "ena0";
defparam ram_block1a62.clk0_input_clock_enable = "ena2";
defparam ram_block1a62.clk1_core_clock_enable = "ena3";
defparam ram_block1a62.clk1_input_clock_enable = "ena3";
defparam ram_block1a62.clk1_output_clock_enable = "ena1";
defparam ram_block1a62.clock_duty_cycle_dependence = "on";
defparam ram_block1a62.data_interleave_offset_in_bits = 1;
defparam ram_block1a62.data_interleave_width_in_bits = 1;
defparam ram_block1a62.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a62.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a62.operation_mode = "dual_port";
defparam ram_block1a62.port_a_address_clear = "none";
defparam ram_block1a62.port_a_address_width = 8;
defparam ram_block1a62.port_a_data_out_clear = "none";
defparam ram_block1a62.port_a_data_out_clock = "none";
defparam ram_block1a62.port_a_data_width = 1;
defparam ram_block1a62.port_a_first_address = 0;
defparam ram_block1a62.port_a_first_bit_number = 62;
defparam ram_block1a62.port_a_last_address = 255;
defparam ram_block1a62.port_a_logical_ram_depth = 256;
defparam ram_block1a62.port_a_logical_ram_width = 144;
defparam ram_block1a62.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a62.port_b_address_clear = "none";
defparam ram_block1a62.port_b_address_clock = "clock1";
defparam ram_block1a62.port_b_address_width = 8;
defparam ram_block1a62.port_b_data_out_clear = "none";
defparam ram_block1a62.port_b_data_out_clock = "clock1";
defparam ram_block1a62.port_b_data_width = 1;
defparam ram_block1a62.port_b_first_address = 0;
defparam ram_block1a62.port_b_first_bit_number = 62;
defparam ram_block1a62.port_b_last_address = 255;
defparam ram_block1a62.port_b_logical_ram_depth = 256;
defparam ram_block1a62.port_b_logical_ram_width = 144;
defparam ram_block1a62.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a62.port_b_read_enable_clock = "clock1";
defparam ram_block1a62.ram_block_type = "auto";

arriaii_ram_block ram_block1a94(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[94]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a94_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a94.clk0_core_clock_enable = "ena0";
defparam ram_block1a94.clk0_input_clock_enable = "ena2";
defparam ram_block1a94.clk1_core_clock_enable = "ena3";
defparam ram_block1a94.clk1_input_clock_enable = "ena3";
defparam ram_block1a94.clk1_output_clock_enable = "ena1";
defparam ram_block1a94.clock_duty_cycle_dependence = "on";
defparam ram_block1a94.data_interleave_offset_in_bits = 1;
defparam ram_block1a94.data_interleave_width_in_bits = 1;
defparam ram_block1a94.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a94.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a94.operation_mode = "dual_port";
defparam ram_block1a94.port_a_address_clear = "none";
defparam ram_block1a94.port_a_address_width = 8;
defparam ram_block1a94.port_a_data_out_clear = "none";
defparam ram_block1a94.port_a_data_out_clock = "none";
defparam ram_block1a94.port_a_data_width = 1;
defparam ram_block1a94.port_a_first_address = 0;
defparam ram_block1a94.port_a_first_bit_number = 94;
defparam ram_block1a94.port_a_last_address = 255;
defparam ram_block1a94.port_a_logical_ram_depth = 256;
defparam ram_block1a94.port_a_logical_ram_width = 144;
defparam ram_block1a94.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a94.port_b_address_clear = "none";
defparam ram_block1a94.port_b_address_clock = "clock1";
defparam ram_block1a94.port_b_address_width = 8;
defparam ram_block1a94.port_b_data_out_clear = "none";
defparam ram_block1a94.port_b_data_out_clock = "clock1";
defparam ram_block1a94.port_b_data_width = 1;
defparam ram_block1a94.port_b_first_address = 0;
defparam ram_block1a94.port_b_first_bit_number = 94;
defparam ram_block1a94.port_b_last_address = 255;
defparam ram_block1a94.port_b_logical_ram_depth = 256;
defparam ram_block1a94.port_b_logical_ram_width = 144;
defparam ram_block1a94.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a94.port_b_read_enable_clock = "clock1";
defparam ram_block1a94.ram_block_type = "auto";

arriaii_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk0_input_clock_enable = "ena2";
defparam ram_block1a30.clk1_core_clock_enable = "ena3";
defparam ram_block1a30.clk1_input_clock_enable = "ena3";
defparam ram_block1a30.clk1_output_clock_enable = "ena1";
defparam ram_block1a30.clock_duty_cycle_dependence = "on";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 8;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 255;
defparam ram_block1a30.port_a_logical_ram_depth = 256;
defparam ram_block1a30.port_a_logical_ram_width = 144;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock1";
defparam ram_block1a30.port_b_address_width = 8;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "clock1";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 255;
defparam ram_block1a30.port_b_logical_ram_depth = 256;
defparam ram_block1a30.port_b_logical_ram_width = 144;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock1";
defparam ram_block1a30.ram_block_type = "auto";

arriaii_ram_block ram_block1a127(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[127]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a127_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a127.clk0_core_clock_enable = "ena0";
defparam ram_block1a127.clk0_input_clock_enable = "ena2";
defparam ram_block1a127.clk1_core_clock_enable = "ena3";
defparam ram_block1a127.clk1_input_clock_enable = "ena3";
defparam ram_block1a127.clk1_output_clock_enable = "ena1";
defparam ram_block1a127.clock_duty_cycle_dependence = "on";
defparam ram_block1a127.data_interleave_offset_in_bits = 1;
defparam ram_block1a127.data_interleave_width_in_bits = 1;
defparam ram_block1a127.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a127.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a127.operation_mode = "dual_port";
defparam ram_block1a127.port_a_address_clear = "none";
defparam ram_block1a127.port_a_address_width = 8;
defparam ram_block1a127.port_a_data_out_clear = "none";
defparam ram_block1a127.port_a_data_out_clock = "none";
defparam ram_block1a127.port_a_data_width = 1;
defparam ram_block1a127.port_a_first_address = 0;
defparam ram_block1a127.port_a_first_bit_number = 127;
defparam ram_block1a127.port_a_last_address = 255;
defparam ram_block1a127.port_a_logical_ram_depth = 256;
defparam ram_block1a127.port_a_logical_ram_width = 144;
defparam ram_block1a127.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a127.port_b_address_clear = "none";
defparam ram_block1a127.port_b_address_clock = "clock1";
defparam ram_block1a127.port_b_address_width = 8;
defparam ram_block1a127.port_b_data_out_clear = "none";
defparam ram_block1a127.port_b_data_out_clock = "clock1";
defparam ram_block1a127.port_b_data_width = 1;
defparam ram_block1a127.port_b_first_address = 0;
defparam ram_block1a127.port_b_first_bit_number = 127;
defparam ram_block1a127.port_b_last_address = 255;
defparam ram_block1a127.port_b_logical_ram_depth = 256;
defparam ram_block1a127.port_b_logical_ram_width = 144;
defparam ram_block1a127.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a127.port_b_read_enable_clock = "clock1";
defparam ram_block1a127.ram_block_type = "auto";

arriaii_ram_block ram_block1a63(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[63]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a63_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a63.clk0_core_clock_enable = "ena0";
defparam ram_block1a63.clk0_input_clock_enable = "ena2";
defparam ram_block1a63.clk1_core_clock_enable = "ena3";
defparam ram_block1a63.clk1_input_clock_enable = "ena3";
defparam ram_block1a63.clk1_output_clock_enable = "ena1";
defparam ram_block1a63.clock_duty_cycle_dependence = "on";
defparam ram_block1a63.data_interleave_offset_in_bits = 1;
defparam ram_block1a63.data_interleave_width_in_bits = 1;
defparam ram_block1a63.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a63.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a63.operation_mode = "dual_port";
defparam ram_block1a63.port_a_address_clear = "none";
defparam ram_block1a63.port_a_address_width = 8;
defparam ram_block1a63.port_a_data_out_clear = "none";
defparam ram_block1a63.port_a_data_out_clock = "none";
defparam ram_block1a63.port_a_data_width = 1;
defparam ram_block1a63.port_a_first_address = 0;
defparam ram_block1a63.port_a_first_bit_number = 63;
defparam ram_block1a63.port_a_last_address = 255;
defparam ram_block1a63.port_a_logical_ram_depth = 256;
defparam ram_block1a63.port_a_logical_ram_width = 144;
defparam ram_block1a63.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a63.port_b_address_clear = "none";
defparam ram_block1a63.port_b_address_clock = "clock1";
defparam ram_block1a63.port_b_address_width = 8;
defparam ram_block1a63.port_b_data_out_clear = "none";
defparam ram_block1a63.port_b_data_out_clock = "clock1";
defparam ram_block1a63.port_b_data_width = 1;
defparam ram_block1a63.port_b_first_address = 0;
defparam ram_block1a63.port_b_first_bit_number = 63;
defparam ram_block1a63.port_b_last_address = 255;
defparam ram_block1a63.port_b_logical_ram_depth = 256;
defparam ram_block1a63.port_b_logical_ram_width = 144;
defparam ram_block1a63.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a63.port_b_read_enable_clock = "clock1";
defparam ram_block1a63.ram_block_type = "auto";

arriaii_ram_block ram_block1a95(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[95]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a95_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a95.clk0_core_clock_enable = "ena0";
defparam ram_block1a95.clk0_input_clock_enable = "ena2";
defparam ram_block1a95.clk1_core_clock_enable = "ena3";
defparam ram_block1a95.clk1_input_clock_enable = "ena3";
defparam ram_block1a95.clk1_output_clock_enable = "ena1";
defparam ram_block1a95.clock_duty_cycle_dependence = "on";
defparam ram_block1a95.data_interleave_offset_in_bits = 1;
defparam ram_block1a95.data_interleave_width_in_bits = 1;
defparam ram_block1a95.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a95.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a95.operation_mode = "dual_port";
defparam ram_block1a95.port_a_address_clear = "none";
defparam ram_block1a95.port_a_address_width = 8;
defparam ram_block1a95.port_a_data_out_clear = "none";
defparam ram_block1a95.port_a_data_out_clock = "none";
defparam ram_block1a95.port_a_data_width = 1;
defparam ram_block1a95.port_a_first_address = 0;
defparam ram_block1a95.port_a_first_bit_number = 95;
defparam ram_block1a95.port_a_last_address = 255;
defparam ram_block1a95.port_a_logical_ram_depth = 256;
defparam ram_block1a95.port_a_logical_ram_width = 144;
defparam ram_block1a95.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a95.port_b_address_clear = "none";
defparam ram_block1a95.port_b_address_clock = "clock1";
defparam ram_block1a95.port_b_address_width = 8;
defparam ram_block1a95.port_b_data_out_clear = "none";
defparam ram_block1a95.port_b_data_out_clock = "clock1";
defparam ram_block1a95.port_b_data_width = 1;
defparam ram_block1a95.port_b_first_address = 0;
defparam ram_block1a95.port_b_first_bit_number = 95;
defparam ram_block1a95.port_b_last_address = 255;
defparam ram_block1a95.port_b_logical_ram_depth = 256;
defparam ram_block1a95.port_b_logical_ram_width = 144;
defparam ram_block1a95.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a95.port_b_read_enable_clock = "clock1";
defparam ram_block1a95.ram_block_type = "auto";

arriaii_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk0_input_clock_enable = "ena2";
defparam ram_block1a31.clk1_core_clock_enable = "ena3";
defparam ram_block1a31.clk1_input_clock_enable = "ena3";
defparam ram_block1a31.clk1_output_clock_enable = "ena1";
defparam ram_block1a31.clock_duty_cycle_dependence = "on";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_alt_ddrx_controller_wrapper:ddr3_int_alt_ddrx_controller_wrapper_inst|alt_ddrx_controller:alt_ddrx_controller_inst|alt_ddrx_input_if:input_if_inst|alt_ddrx_wdata_fifo:wdata_fifo_inst|scfifo:wdata_fifo|scfifo_2a61:auto_generated|a_dpfifo_0131:dpfifo|altsyncram_u1e1:FIFOram|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 8;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 255;
defparam ram_block1a31.port_a_logical_ram_depth = 256;
defparam ram_block1a31.port_a_logical_ram_width = 144;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock1";
defparam ram_block1a31.port_b_address_width = 8;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "clock1";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 255;
defparam ram_block1a31.port_b_logical_ram_depth = 256;
defparam ram_block1a31.port_b_logical_ram_width = 144;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock1";
defparam ram_block1a31.ram_block_type = "auto";

endmodule

module ddr3_int_cntr_hkb (
	clock,
	reset_reg_3,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	counter_reg_bit_6,
	_)/* synthesis synthesis_greybox=0 */;
input 	clock;
input 	reset_reg_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
output 	counter_reg_bit_6;
input 	_;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;
wire \counter_comb_bita5~COUT ;
wire \counter_comb_bita6~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[6] (
	.clk(clock),
	.d(\counter_comb_bita6~sumout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_6),
	.prn(vcc));
defparam \counter_reg_bit[6] .is_wysiwyg = "true";
defparam \counter_reg_bit[6] .power_up = "low";

arriaii_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

arriaii_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h0000FFFF000000FF;
defparam counter_comb_bita1.shared_arith = "off";

arriaii_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h0000FFFF000000FF;
defparam counter_comb_bita2.shared_arith = "off";

arriaii_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h0000FFFF000000FF;
defparam counter_comb_bita3.shared_arith = "off";

arriaii_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h0000FFFF000000FF;
defparam counter_comb_bita4.shared_arith = "off";

arriaii_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(\counter_comb_bita5~COUT ),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h0000FFFF000000FF;
defparam counter_comb_bita5.shared_arith = "off";

arriaii_lcell_comb counter_comb_bita6(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita5~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita6~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita6.extended_lut = "off";
defparam counter_comb_bita6.lut_mask = 64'h0000FFFF000000FF;
defparam counter_comb_bita6.shared_arith = "off";

endmodule

module ddr3_int_cntr_ikb (
	clock,
	avalon_write_req,
	reset_reg_3,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	counter_reg_bit_6,
	counter_reg_bit_7)/* synthesis synthesis_greybox=0 */;
input 	clock;
input 	avalon_write_req;
input 	reset_reg_3;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
output 	counter_reg_bit_6;
output 	counter_reg_bit_7;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;
wire \counter_comb_bita5~COUT ;
wire \counter_comb_bita6~sumout ;
wire \counter_comb_bita6~COUT ;
wire \counter_comb_bita7~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(avalon_write_req),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(avalon_write_req),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(avalon_write_req),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(avalon_write_req),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(avalon_write_req),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(avalon_write_req),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[6] (
	.clk(clock),
	.d(\counter_comb_bita6~sumout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(avalon_write_req),
	.q(counter_reg_bit_6),
	.prn(vcc));
defparam \counter_reg_bit[6] .is_wysiwyg = "true";
defparam \counter_reg_bit[6] .power_up = "low";

dffeas \counter_reg_bit[7] (
	.clk(clock),
	.d(\counter_comb_bita7~sumout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(avalon_write_req),
	.q(counter_reg_bit_7),
	.prn(vcc));
defparam \counter_reg_bit[7] .is_wysiwyg = "true";
defparam \counter_reg_bit[7] .power_up = "low";

arriaii_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

arriaii_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h0000FFFF000000FF;
defparam counter_comb_bita1.shared_arith = "off";

arriaii_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h0000FFFF000000FF;
defparam counter_comb_bita2.shared_arith = "off";

arriaii_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h0000FFFF000000FF;
defparam counter_comb_bita3.shared_arith = "off";

arriaii_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h0000FFFF000000FF;
defparam counter_comb_bita4.shared_arith = "off";

arriaii_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(\counter_comb_bita5~COUT ),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h0000FFFF000000FF;
defparam counter_comb_bita5.shared_arith = "off";

arriaii_lcell_comb counter_comb_bita6(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita5~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita6~sumout ),
	.cout(\counter_comb_bita6~COUT ),
	.shareout());
defparam counter_comb_bita6.extended_lut = "off";
defparam counter_comb_bita6.lut_mask = 64'h0000FFFF000000FF;
defparam counter_comb_bita6.shared_arith = "off";

arriaii_lcell_comb counter_comb_bita7(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita6~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita7~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita7.extended_lut = "off";
defparam counter_comb_bita7.lut_mask = 64'h0000FFFF000000FF;
defparam counter_comb_bita7.shared_arith = "off";

endmodule

module ddr3_int_cntr_uk7 (
	clock,
	avalon_write_req,
	counter_reg_bit_5,
	counter_reg_bit_7,
	counter_reg_bit_6,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_4,
	counter_reg_bit_3,
	reset_reg_3,
	_)/* synthesis synthesis_greybox=0 */;
input 	clock;
input 	avalon_write_req;
output 	counter_reg_bit_5;
output 	counter_reg_bit_7;
output 	counter_reg_bit_6;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
input 	reset_reg_3;
input 	_;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;
wire \counter_comb_bita5~COUT ;
wire \counter_comb_bita6~COUT ;
wire \counter_comb_bita7~sumout ;
wire \counter_comb_bita6~sumout ;
wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita3~sumout ;


dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[7] (
	.clk(clock),
	.d(\counter_comb_bita7~sumout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_7),
	.prn(vcc));
defparam \counter_reg_bit[7] .is_wysiwyg = "true";
defparam \counter_reg_bit[7] .power_up = "low";

dffeas \counter_reg_bit[6] (
	.clk(clock),
	.d(\counter_comb_bita6~sumout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_6),
	.prn(vcc));
defparam \counter_reg_bit[6] .is_wysiwyg = "true";
defparam \counter_reg_bit[6] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(reset_reg_3),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

arriaii_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

arriaii_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(!avalon_write_req),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita1.shared_arith = "off";

arriaii_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(!avalon_write_req),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita2.shared_arith = "off";

arriaii_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(!avalon_write_req),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita3.shared_arith = "off";

arriaii_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(!avalon_write_req),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita4.shared_arith = "off";

arriaii_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(!avalon_write_req),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(\counter_comb_bita5~COUT ),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita5.shared_arith = "off";

arriaii_lcell_comb counter_comb_bita6(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_6),
	.datae(gnd),
	.dataf(!avalon_write_req),
	.datag(gnd),
	.cin(\counter_comb_bita5~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita6~sumout ),
	.cout(\counter_comb_bita6~COUT ),
	.shareout());
defparam counter_comb_bita6.extended_lut = "off";
defparam counter_comb_bita6.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita6.shared_arith = "off";

arriaii_lcell_comb counter_comb_bita7(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_7),
	.datae(gnd),
	.dataf(!avalon_write_req),
	.datag(gnd),
	.cin(\counter_comb_bita6~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita7~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita7.extended_lut = "off";
defparam counter_comb_bita7.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita7.shared_arith = "off";

endmodule

module ddr3_int_alt_ddrx_state_machine (
	ctl_clk,
	auto_refresh_logic_per_chip0int_refresh_req,
	out_cmd_info_valid_0,
	do_read_r1,
	do_auto_precharge_r1,
	do_write_r1,
	out_cmd_info_valid_2,
	out_cmd_info_valid_3,
	out_cmd_info_valid_4,
	out_cmd_info_valid_1,
	pipe_10_0,
	pipe_12_0,
	pipe_11_0,
	pipe_32_0,
	pipe_12_2,
	pipe_12_3,
	pipe_12_1,
	pipe_10_2,
	pipe_10_3,
	pipe_10_1,
	pipe_11_2,
	pipe_11_3,
	pipe_11_1,
	pipe_29_0,
	pipe_28_0,
	pipe_33_0,
	do_burst_chop_r1,
	pipe_12_4,
	pipe_11_4,
	pipe_10_4,
	pipe_25_5,
	pipe_25_0,
	pipe_26_5,
	pipe_26_0,
	pipe_24_5,
	pipe_24_0,
	pipe_22_5,
	pipe_22_0,
	pipe_23_5,
	pipe_23_0,
	pipe_21_5,
	pipe_21_0,
	pipe_19_5,
	pipe_19_0,
	pipe_20_5,
	pipe_20_0,
	pipe_15_5,
	pipe_15_0,
	pipe_13_5,
	pipe_13_0,
	pipe_14_5,
	pipe_14_0,
	pipe_18_5,
	pipe_18_0,
	pipe_16_5,
	pipe_16_0,
	pipe_17_5,
	pipe_17_0,
	pipe_12_5,
	pipe_11_5,
	pipe_10_5,
	pipe_25_3,
	pipe_26_3,
	pipe_24_3,
	pipe_22_3,
	pipe_23_3,
	pipe_21_3,
	pipe_19_3,
	pipe_20_3,
	pipe_15_3,
	pipe_13_3,
	pipe_14_3,
	pipe_18_3,
	pipe_16_3,
	pipe_17_3,
	pipe_25_4,
	pipe_26_4,
	pipe_24_4,
	pipe_22_4,
	pipe_23_4,
	pipe_21_4,
	pipe_19_4,
	pipe_20_4,
	pipe_15_4,
	pipe_13_4,
	pipe_14_4,
	pipe_18_4,
	pipe_16_4,
	pipe_17_4,
	pipe_12_6,
	pipe_11_6,
	pipe_10_6,
	pipe_25_6,
	pipe_26_6,
	pipe_24_6,
	pipe_22_6,
	pipe_23_6,
	pipe_21_6,
	pipe_19_6,
	pipe_20_6,
	pipe_15_6,
	pipe_13_6,
	pipe_14_6,
	pipe_18_6,
	pipe_16_6,
	pipe_17_6,
	pipe_26_7,
	pipe_24_7,
	pipe_25_7,
	pipe_23_7,
	pipe_21_7,
	pipe_22_7,
	pipe_20_7,
	pipe_18_7,
	pipe_19_7,
	pipe_17_7,
	pipe_15_7,
	pipe_16_7,
	pipe_11_7,
	pipe_10_7,
	pipe_14_7,
	pipe_12_7,
	pipe_13_7,
	pipe_25_2,
	pipe_26_2,
	pipe_24_2,
	pipe_22_2,
	pipe_23_2,
	pipe_21_2,
	pipe_19_2,
	pipe_20_2,
	pipe_15_2,
	pipe_13_2,
	pipe_14_2,
	pipe_18_2,
	pipe_16_2,
	pipe_17_2,
	pipe_25_1,
	pipe_26_1,
	pipe_24_1,
	pipe_22_1,
	pipe_23_1,
	pipe_21_1,
	pipe_19_1,
	pipe_20_1,
	pipe_15_1,
	pipe_13_1,
	pipe_14_1,
	pipe_18_1,
	pipe_16_1,
	pipe_17_1,
	pipe_2_0,
	to_row_addr_r_0,
	to_row_addr_r_1,
	to_col_addr_r_2,
	to_row_addr_r_2,
	to_col_addr_r_3,
	to_row_addr_r_3,
	to_col_addr_r_4,
	to_row_addr_r_4,
	to_col_addr_r_5,
	to_row_addr_r_5,
	to_col_addr_r_6,
	to_row_addr_r_6,
	to_col_addr_r_7,
	to_row_addr_r_7,
	to_col_addr_r_8,
	to_row_addr_r_8,
	to_col_addr_r_9,
	to_row_addr_r_9,
	to_row_addr_r_10,
	to_row_addr_r_11,
	to_row_addr_r_12,
	to_row_addr_r_13,
	pipe_3_0,
	pipe_4_0,
	pipe_5_0,
	pipe_6_0,
	pipe_7_0,
	pipe_8_0,
	pipe_9_0,
	hold_ready,
	pipefull_7,
	int_refresh_ack1,
	ctl_init_success,
	internal_ready,
	avalon_write_req,
	fetch1,
	read_req,
	write_req,
	pipefull_6,
	do_precharge_all_r1,
	out_cs_can_refresh_0,
	ctl_reset_n,
	always38,
	pipefull_0,
	do_refresh_r1,
	add_lat_on,
	out_cmd_can_activate_0,
	out_cmd_bank_is_open_0,
	can_al_activate_write,
	to_chip_r_0,
	always381,
	to_bank_addr_r_2,
	current_bank_2,
	to_bank_addr_r_0,
	current_bank_0,
	to_bank_addr_r_1,
	current_bank_1,
	always382,
	out_cmd_can_write_0,
	can_al_activate_read,
	out_cmd_can_read_0,
	pipefull_5,
	rdwr_data_valid_r1,
	out_cs_all_banks_closed_0,
	out_cs_can_precharge_all_0,
	do_activate_r1,
	pipefull_1,
	out_cmd_can_activate_2,
	out_cmd_bank_is_open_2,
	out_cmd_can_activate_3,
	out_cmd_bank_is_open_3,
	out_cmd_can_activate_4,
	out_cmd_bank_is_open_4,
	out_cmd_can_activate_1,
	out_cmd_bank_is_open_1,
	pipefull_4,
	pipefull_2,
	pipefull_3,
	local_write_req)/* synthesis synthesis_greybox=0 */;
input 	ctl_clk;
input 	auto_refresh_logic_per_chip0int_refresh_req;
input 	out_cmd_info_valid_0;
output 	do_read_r1;
output 	do_auto_precharge_r1;
output 	do_write_r1;
input 	out_cmd_info_valid_2;
input 	out_cmd_info_valid_3;
input 	out_cmd_info_valid_4;
input 	out_cmd_info_valid_1;
input 	pipe_10_0;
input 	pipe_12_0;
input 	pipe_11_0;
input 	pipe_32_0;
input 	pipe_12_2;
input 	pipe_12_3;
input 	pipe_12_1;
input 	pipe_10_2;
input 	pipe_10_3;
input 	pipe_10_1;
input 	pipe_11_2;
input 	pipe_11_3;
input 	pipe_11_1;
input 	pipe_29_0;
input 	pipe_28_0;
input 	pipe_33_0;
output 	do_burst_chop_r1;
input 	pipe_12_4;
input 	pipe_11_4;
input 	pipe_10_4;
input 	pipe_25_5;
input 	pipe_25_0;
input 	pipe_26_5;
input 	pipe_26_0;
input 	pipe_24_5;
input 	pipe_24_0;
input 	pipe_22_5;
input 	pipe_22_0;
input 	pipe_23_5;
input 	pipe_23_0;
input 	pipe_21_5;
input 	pipe_21_0;
input 	pipe_19_5;
input 	pipe_19_0;
input 	pipe_20_5;
input 	pipe_20_0;
input 	pipe_15_5;
input 	pipe_15_0;
input 	pipe_13_5;
input 	pipe_13_0;
input 	pipe_14_5;
input 	pipe_14_0;
input 	pipe_18_5;
input 	pipe_18_0;
input 	pipe_16_5;
input 	pipe_16_0;
input 	pipe_17_5;
input 	pipe_17_0;
input 	pipe_12_5;
input 	pipe_11_5;
input 	pipe_10_5;
input 	pipe_25_3;
input 	pipe_26_3;
input 	pipe_24_3;
input 	pipe_22_3;
input 	pipe_23_3;
input 	pipe_21_3;
input 	pipe_19_3;
input 	pipe_20_3;
input 	pipe_15_3;
input 	pipe_13_3;
input 	pipe_14_3;
input 	pipe_18_3;
input 	pipe_16_3;
input 	pipe_17_3;
input 	pipe_25_4;
input 	pipe_26_4;
input 	pipe_24_4;
input 	pipe_22_4;
input 	pipe_23_4;
input 	pipe_21_4;
input 	pipe_19_4;
input 	pipe_20_4;
input 	pipe_15_4;
input 	pipe_13_4;
input 	pipe_14_4;
input 	pipe_18_4;
input 	pipe_16_4;
input 	pipe_17_4;
input 	pipe_12_6;
input 	pipe_11_6;
input 	pipe_10_6;
input 	pipe_25_6;
input 	pipe_26_6;
input 	pipe_24_6;
input 	pipe_22_6;
input 	pipe_23_6;
input 	pipe_21_6;
input 	pipe_19_6;
input 	pipe_20_6;
input 	pipe_15_6;
input 	pipe_13_6;
input 	pipe_14_6;
input 	pipe_18_6;
input 	pipe_16_6;
input 	pipe_17_6;
input 	pipe_26_7;
input 	pipe_24_7;
input 	pipe_25_7;
input 	pipe_23_7;
input 	pipe_21_7;
input 	pipe_22_7;
input 	pipe_20_7;
input 	pipe_18_7;
input 	pipe_19_7;
input 	pipe_17_7;
input 	pipe_15_7;
input 	pipe_16_7;
input 	pipe_11_7;
input 	pipe_10_7;
input 	pipe_14_7;
input 	pipe_12_7;
input 	pipe_13_7;
input 	pipe_25_2;
input 	pipe_26_2;
input 	pipe_24_2;
input 	pipe_22_2;
input 	pipe_23_2;
input 	pipe_21_2;
input 	pipe_19_2;
input 	pipe_20_2;
input 	pipe_15_2;
input 	pipe_13_2;
input 	pipe_14_2;
input 	pipe_18_2;
input 	pipe_16_2;
input 	pipe_17_2;
input 	pipe_25_1;
input 	pipe_26_1;
input 	pipe_24_1;
input 	pipe_22_1;
input 	pipe_23_1;
input 	pipe_21_1;
input 	pipe_19_1;
input 	pipe_20_1;
input 	pipe_15_1;
input 	pipe_13_1;
input 	pipe_14_1;
input 	pipe_18_1;
input 	pipe_16_1;
input 	pipe_17_1;
input 	pipe_2_0;
output 	to_row_addr_r_0;
output 	to_row_addr_r_1;
output 	to_col_addr_r_2;
output 	to_row_addr_r_2;
output 	to_col_addr_r_3;
output 	to_row_addr_r_3;
output 	to_col_addr_r_4;
output 	to_row_addr_r_4;
output 	to_col_addr_r_5;
output 	to_row_addr_r_5;
output 	to_col_addr_r_6;
output 	to_row_addr_r_6;
output 	to_col_addr_r_7;
output 	to_row_addr_r_7;
output 	to_col_addr_r_8;
output 	to_row_addr_r_8;
output 	to_col_addr_r_9;
output 	to_row_addr_r_9;
output 	to_row_addr_r_10;
output 	to_row_addr_r_11;
output 	to_row_addr_r_12;
output 	to_row_addr_r_13;
input 	pipe_3_0;
input 	pipe_4_0;
input 	pipe_5_0;
input 	pipe_6_0;
input 	pipe_7_0;
input 	pipe_8_0;
input 	pipe_9_0;
input 	hold_ready;
input 	pipefull_7;
output 	int_refresh_ack1;
input 	ctl_init_success;
input 	internal_ready;
input 	avalon_write_req;
output 	fetch1;
input 	read_req;
input 	write_req;
input 	pipefull_6;
output 	do_precharge_all_r1;
input 	out_cs_can_refresh_0;
input 	ctl_reset_n;
output 	always38;
input 	pipefull_0;
output 	do_refresh_r1;
input 	add_lat_on;
input 	out_cmd_can_activate_0;
input 	out_cmd_bank_is_open_0;
input 	can_al_activate_write;
output 	to_chip_r_0;
output 	always381;
output 	to_bank_addr_r_2;
output 	current_bank_2;
output 	to_bank_addr_r_0;
output 	current_bank_0;
output 	to_bank_addr_r_1;
output 	current_bank_1;
output 	always382;
input 	out_cmd_can_write_0;
input 	can_al_activate_read;
input 	out_cmd_can_read_0;
input 	pipefull_5;
output 	rdwr_data_valid_r1;
input 	out_cs_all_banks_closed_0;
input 	out_cs_can_precharge_all_0;
output 	do_activate_r1;
input 	pipefull_1;
input 	out_cmd_can_activate_2;
input 	out_cmd_bank_is_open_2;
input 	out_cmd_can_activate_3;
input 	out_cmd_bank_is_open_3;
input 	out_cmd_can_activate_4;
input 	out_cmd_bank_is_open_4;
input 	out_cmd_can_activate_1;
input 	out_cmd_bank_is_open_1;
input 	pipefull_4;
input 	pipefull_2;
input 	pipefull_3;
input 	local_write_req;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always38~2_combout ;
wire \always38~7_combout ;
wire \Equal47~0_combout ;
wire \Equal47~1_combout ;
wire \Equal47~2_combout ;
wire \Equal47~3_combout ;
wire \Equal47~4_combout ;
wire \Equal47~5_combout ;
wire \Equal41~0_combout ;
wire \Equal44~0_combout ;
wire \auto_autopch_req_0~2_combout ;
wire \auto_autopch_req_c~0_combout ;
wire \auto_autopch_req_c~1_combout ;
wire \auto_autopch_req_c~2_combout ;
wire \auto_autopch_req_c~3_combout ;
wire \auto_autopch_req_c~4_combout ;
wire \auto_autopch_req_c~5_combout ;
wire \auto_autopch_req_c~6_combout ;
wire \always14~2_combout ;
wire \always14~3_combout ;
wire \always14~4_combout ;
wire \always14~5_combout ;
wire \Equal29~0_combout ;
wire \Equal29~1_combout ;
wire \Equal29~2_combout ;
wire \Equal29~3_combout ;
wire \Equal29~4_combout ;
wire \Equal29~5_combout ;
wire \Equal32~0_combout ;
wire \Equal32~1_combout ;
wire \Equal32~2_combout ;
wire \Equal32~3_combout ;
wire \Equal32~4_combout ;
wire \Equal32~5_combout ;
wire \auto_autopch_req_c~7_combout ;
wire \always14~6_combout ;
wire \Equal22~0_combout ;
wire \Equal20~0_combout ;
wire \Equal21~0_combout ;
wire \Equal23~1_combout ;
wire \current_read~q ;
wire \always38~5_combout ;
wire \always38~6_combout ;
wire \current_burstcount_counter_temp[0]~q ;
wire \Selector19~0_combout ;
wire \start_burst~q ;
wire \start_burst_r~q ;
wire \current_col[2]~q ;
wire \burst_delay~0_combout ;
wire \burst_delay~q ;
wire \always29~0_combout ;
wire \current_burstcount_counter[0]~0_combout ;
wire \current_burstcount_counter[0]~q ;
wire \write_burst_length~0_combout ;
wire \start_write_burst_r~q ;
wire \current_write~q ;
wire \always17~0_combout ;
wire \Add0~2_sumout ;
wire \proper_beats_in_fifo[9]~0_combout ;
wire \proper_beats_in_fifo[0]~q ;
wire \Add0~3 ;
wire \Add0~6_sumout ;
wire \proper_beats_in_fifo[1]~q ;
wire \always38~8_combout ;
wire \Add0~7 ;
wire \Add0~10_sumout ;
wire \proper_beats_in_fifo[2]~q ;
wire \Add0~11 ;
wire \Add0~14_sumout ;
wire \proper_beats_in_fifo[3]~q ;
wire \Add0~15 ;
wire \Add0~18_sumout ;
wire \proper_beats_in_fifo[4]~q ;
wire \Add0~19 ;
wire \Add0~22_sumout ;
wire \proper_beats_in_fifo[5]~q ;
wire \Add0~23 ;
wire \Add0~26_sumout ;
wire \proper_beats_in_fifo[6]~q ;
wire \Add0~27 ;
wire \Add0~30_sumout ;
wire \proper_beats_in_fifo[7]~q ;
wire \Add0~31 ;
wire \Add0~34_sumout ;
wire \proper_beats_in_fifo[8]~q ;
wire \Add0~35 ;
wire \Add0~38_sumout ;
wire \proper_beats_in_fifo[9]~q ;
wire \always38~9_combout ;
wire \current_burstcount_counter_temp[1]~q ;
wire \always38~10_combout ;
wire \always38~11_combout ;
wire \always38~1_combout ;
wire \Selector20~0_combout ;
wire \always14~0_combout ;
wire \Equal4~0_combout ;
wire \always11~0_combout ;
wire \always12~0_combout ;
wire \Equal8~0_combout ;
wire \Equal6~0_combout ;
wire \always12~1_combout ;
wire \always12~2_combout ;
wire \Equal18~0_combout ;
wire \Equal16~0_combout ;
wire \Equal14~0_combout ;
wire \Equal12~0_combout ;
wire \always13~0_combout ;
wire \always13~1_combout ;
wire \lookahead_allowed_to_cmd[3]~q ;
wire \lookahead_allowed_to_cmd[2]~q ;
wire \lookahead_allowed_to_cmd[1]~q ;
wire \always39~0_combout ;
wire \always39~1_combout ;
wire \always14~1_combout ;
wire \always10~0_combout ;
wire \lookahead_allowed_to_cmd[0]~q ;
wire \always39~2_combout ;
wire \to_bank_addr_r[2]~0_combout ;
wire \Selector20~1_combout ;
wire \Selector20~2_combout ;
wire \just_did_activate~q ;
wire \always38~12_combout ;
wire \always38~13_combout ;
wire \always38~14_combout ;
wire \always38~15_combout ;
wire \Selector6~0_combout ;
wire \state.READWRITE~q ;
wire \always15~1_combout ;
wire \always15~2_combout ;
wire \Equal50~0_combout ;
wire \Equal50~1_combout ;
wire \Equal50~2_combout ;
wire \Equal50~3_combout ;
wire \Equal50~4_combout ;
wire \Equal50~5_combout ;
wire \Equal50~6_combout ;
wire \always15~0_combout ;
wire \always15~5_combout ;
wire \always15~6_combout ;
wire \always15~3_combout ;
wire \always15~4_combout ;
wire \Equal41~1_combout ;
wire \Equal41~2_combout ;
wire \Equal41~3_combout ;
wire \Equal41~4_combout ;
wire \Equal41~5_combout ;
wire \Equal44~1_combout ;
wire \Equal44~2_combout ;
wire \Equal44~3_combout ;
wire \Equal44~4_combout ;
wire \Equal44~5_combout ;
wire \auto_autopch_req~0_combout ;
wire \auto_autopch_req_0~0_combout ;
wire \auto_autopch_req_0~1_combout ;
wire \auto_autopch_req_0~3_combout ;
wire \auto_autopch_req_0~4_combout ;
wire \auto_autopch_req_0~5_combout ;
wire \auto_autopch_req_0~6_combout ;
wire \auto_autopch_req_0~7_combout ;
wire \auto_autopch_req~4_combout ;
wire \auto_autopch_req~1_combout ;
wire \always14~7_combout ;
wire \always14~8_combout ;
wire \always14~9_combout ;
wire \auto_autopch_req_c~8_combout ;
wire \always14~10_combout ;
wire \always14~11_combout ;
wire \current_row[10]~q ;
wire \current_row[9]~q ;
wire \Equal22~1_combout ;
wire \current_row[7]~q ;
wire \current_row[6]~q ;
wire \Equal22~2_combout ;
wire \current_row[1]~q ;
wire \current_row[0]~q ;
wire \Equal22~3_combout ;
wire \current_row[4]~q ;
wire \current_row[3]~q ;
wire \Equal22~4_combout ;
wire \Equal22~5_combout ;
wire \current_row[11]~q ;
wire \Equal20~1_combout ;
wire \current_row[8]~q ;
wire \Equal20~2_combout ;
wire \current_row[2]~q ;
wire \Equal20~3_combout ;
wire \current_row[5]~q ;
wire \Equal20~4_combout ;
wire \Equal20~5_combout ;
wire \Equal21~1_combout ;
wire \Equal21~2_combout ;
wire \Equal21~3_combout ;
wire \Equal21~4_combout ;
wire \Equal21~5_combout ;
wire \auto_autopch_req_c~9_combout ;
wire \current_row[13]~q ;
wire \current_row[12]~q ;
wire \Equal23~0_combout ;
wire \Equal23~2_combout ;
wire \Equal23~3_combout ;
wire \Equal23~4_combout ;
wire \Equal23~5_combout ;
wire \auto_autopch_req_c~10_combout ;
wire \Equal26~0_combout ;
wire \Equal26~1_combout ;
wire \Equal26~2_combout ;
wire \Equal26~3_combout ;
wire \Equal26~4_combout ;
wire \Equal26~5_combout ;
wire \Equal26~6_combout ;
wire \auto_autopch_req_c~11_combout ;
wire \always15~7_combout ;
wire \Equal37~0_combout ;
wire \Equal37~1_combout ;
wire \Equal37~2_combout ;
wire \Equal37~3_combout ;
wire \Equal37~4_combout ;
wire \Equal37~5_combout ;
wire \Equal37~6_combout ;
wire \Equal39~0_combout ;
wire \Equal39~1_combout ;
wire \Equal39~2_combout ;
wire \Equal39~3_combout ;
wire \Equal39~4_combout ;
wire \Equal39~5_combout ;
wire \Equal39~6_combout ;
wire \auto_autopch_req~2_combout ;
wire \auto_autopch_req~3_combout ;
wire \auto_autopch_req~q ;
wire \do_auto_precharge~0_combout ;
wire \current_read~_wirecell_combout ;
wire \fetch_r~q ;
wire \current_burstcount_counter[1]~1_combout ;
wire \current_burstcount_counter[1]~q ;
wire \always39~3_combout ;
wire \to_row_addr_r[5]~0_combout ;
wire \to_row_addr_r[5]~1_combout ;
wire \Selector39~0_combout ;
wire \to_bank_addr_r[2]~1_combout ;
wire \state.INIT~0_combout ;
wire \state.INIT~q ;
wire \to_bank_addr_r[2]~2_combout ;
wire \to_row_addr_r[5]~2_combout ;
wire \Selector38~0_combout ;
wire \to_addr~0_combout ;
wire \Selector37~0_combout ;
wire \current_col[3]~q ;
wire \Selector36~0_combout ;
wire \current_col[4]~q ;
wire \Selector35~0_combout ;
wire \current_col[5]~q ;
wire \Selector34~0_combout ;
wire \current_col[6]~q ;
wire \Selector33~0_combout ;
wire \current_col[7]~q ;
wire \Selector32~0_combout ;
wire \current_col[8]~q ;
wire \Selector31~0_combout ;
wire \current_col[9]~q ;
wire \Selector30~0_combout ;
wire \Selector29~0_combout ;
wire \Selector28~0_combout ;
wire \Selector27~0_combout ;
wire \Selector26~0_combout ;
wire \Selector2~0_combout ;
wire \Selector15~0_combout ;
wire \for_chip_refresh_req~q ;
wire \Selector2~1_combout ;
wire \Selector2~2_combout ;
wire \state.FETCH~q ;
wire \Selector7~0_combout ;
wire \Selector4~1_combout ;
wire \state.PCHALL~q ;
wire \Selector4~0_combout ;
wire \Selector7~1_combout ;
wire \state.REFRESH~q ;
wire \Selector0~0_combout ;
wire \Selector0~1_combout ;
wire \state.DO2~q ;
wire \Selector11~1_combout ;
wire \Selector14~0_combout ;
wire \Selector14~1_combout ;
wire \for_chip_saved[0]~0_combout ;
wire \for_chip_saved[0]~q ;
wire \Selector14~2_combout ;
wire \Selector14~3_combout ;
wire \for_chip[0]~q ;
wire \Selector10~0_combout ;
wire \Selector10~1_combout ;
wire \Selector11~0_combout ;
wire \Selector11~2_combout ;
wire \do_precharge_all~0_combout ;
wire \Selector22~0_combout ;
wire \Selector23~0_combout ;
wire \Selector23~1_combout ;
wire \Selector25~0_combout ;
wire \Selector25~1_combout ;
wire \Selector24~0_combout ;
wire \Selector24~1_combout ;
wire \new_gen_rdwr_data_valid~0_combout ;


arriaii_lcell_comb \always38~2 (
	.dataa(!add_lat_on),
	.datab(!\always38~1_combout ),
	.datac(!can_al_activate_write),
	.datad(!\current_write~q ),
	.datae(!do_read_r1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always38~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always38~2 .extended_lut = "off";
defparam \always38~2 .lut_mask = 64'h0001000000010000;
defparam \always38~2 .shared_arith = "off";

arriaii_lcell_comb \always38~7 (
	.dataa(!\fetch_r~q ),
	.datab(!\current_burstcount_counter[1]~q ),
	.datac(!\current_burstcount_counter[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always38~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always38~7 .extended_lut = "off";
defparam \always38~7 .lut_mask = 64'h0808080808080808;
defparam \always38~7 .shared_arith = "off";

arriaii_lcell_comb \Equal47~0 (
	.dataa(!pipe_25_5),
	.datab(!pipe_25_0),
	.datac(!pipe_26_5),
	.datad(!pipe_26_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal47~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal47~0 .extended_lut = "off";
defparam \Equal47~0 .lut_mask = 64'h9009900990099009;
defparam \Equal47~0 .shared_arith = "off";

arriaii_lcell_comb \Equal47~1 (
	.dataa(!pipe_24_5),
	.datab(!pipe_24_0),
	.datac(!pipe_22_5),
	.datad(!pipe_22_0),
	.datae(!pipe_23_5),
	.dataf(!pipe_23_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal47~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal47~1 .extended_lut = "off";
defparam \Equal47~1 .lut_mask = 64'h9009000000009009;
defparam \Equal47~1 .shared_arith = "off";

arriaii_lcell_comb \Equal47~2 (
	.dataa(!pipe_21_5),
	.datab(!pipe_21_0),
	.datac(!pipe_19_5),
	.datad(!pipe_19_0),
	.datae(!pipe_20_5),
	.dataf(!pipe_20_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal47~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal47~2 .extended_lut = "off";
defparam \Equal47~2 .lut_mask = 64'h9009000000009009;
defparam \Equal47~2 .shared_arith = "off";

arriaii_lcell_comb \Equal47~3 (
	.dataa(!pipe_15_5),
	.datab(!pipe_15_0),
	.datac(!pipe_13_5),
	.datad(!pipe_13_0),
	.datae(!pipe_14_5),
	.dataf(!pipe_14_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal47~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal47~3 .extended_lut = "off";
defparam \Equal47~3 .lut_mask = 64'h9009000000009009;
defparam \Equal47~3 .shared_arith = "off";

arriaii_lcell_comb \Equal47~4 (
	.dataa(!pipe_18_5),
	.datab(!pipe_18_0),
	.datac(!pipe_16_5),
	.datad(!pipe_16_0),
	.datae(!pipe_17_5),
	.dataf(!pipe_17_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal47~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal47~4 .extended_lut = "off";
defparam \Equal47~4 .lut_mask = 64'h9009000000009009;
defparam \Equal47~4 .shared_arith = "off";

arriaii_lcell_comb \Equal47~5 (
	.dataa(!\Equal47~0_combout ),
	.datab(!\Equal47~1_combout ),
	.datac(!\Equal47~2_combout ),
	.datad(!\Equal47~3_combout ),
	.datae(!\Equal47~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal47~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal47~5 .extended_lut = "off";
defparam \Equal47~5 .lut_mask = 64'h0000000100000001;
defparam \Equal47~5 .shared_arith = "off";

arriaii_lcell_comb \Equal41~0 (
	.dataa(!pipe_25_0),
	.datab(!pipe_26_0),
	.datac(!pipe_25_3),
	.datad(!pipe_26_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal41~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal41~0 .extended_lut = "off";
defparam \Equal41~0 .lut_mask = 64'h8421842184218421;
defparam \Equal41~0 .shared_arith = "off";

arriaii_lcell_comb \Equal44~0 (
	.dataa(!pipe_25_0),
	.datab(!pipe_26_0),
	.datac(!pipe_25_4),
	.datad(!pipe_26_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal44~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal44~0 .extended_lut = "off";
defparam \Equal44~0 .lut_mask = 64'h8421842184218421;
defparam \Equal44~0 .shared_arith = "off";

arriaii_lcell_comb \auto_autopch_req_0~2 (
	.dataa(!pipe_19_0),
	.datab(!pipe_20_0),
	.datac(!pipe_18_0),
	.datad(!pipe_20_7),
	.datae(!pipe_18_7),
	.dataf(!pipe_19_7),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_autopch_req_0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_autopch_req_0~2 .extended_lut = "off";
defparam \auto_autopch_req_0~2 .lut_mask = 64'h8020080240100401;
defparam \auto_autopch_req_0~2 .shared_arith = "off";

arriaii_lcell_comb \auto_autopch_req_c~0 (
	.dataa(!pipe_26_7),
	.datab(!pipe_24_7),
	.datac(!pipe_25_7),
	.datad(!\current_row[13]~q ),
	.datae(!\current_row[11]~q ),
	.dataf(!\current_row[12]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_autopch_req_c~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_autopch_req_c~0 .extended_lut = "off";
defparam \auto_autopch_req_c~0 .lut_mask = 64'h8040201008040201;
defparam \auto_autopch_req_c~0 .shared_arith = "off";

arriaii_lcell_comb \auto_autopch_req_c~1 (
	.dataa(!pipe_23_7),
	.datab(!pipe_21_7),
	.datac(!pipe_22_7),
	.datad(!\current_row[10]~q ),
	.datae(!\current_row[8]~q ),
	.dataf(!\current_row[9]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_autopch_req_c~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_autopch_req_c~1 .extended_lut = "off";
defparam \auto_autopch_req_c~1 .lut_mask = 64'h8040201008040201;
defparam \auto_autopch_req_c~1 .shared_arith = "off";

arriaii_lcell_comb \auto_autopch_req_c~2 (
	.dataa(!pipe_20_7),
	.datab(!pipe_18_7),
	.datac(!pipe_19_7),
	.datad(!\current_row[7]~q ),
	.datae(!\current_row[5]~q ),
	.dataf(!\current_row[6]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_autopch_req_c~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_autopch_req_c~2 .extended_lut = "off";
defparam \auto_autopch_req_c~2 .lut_mask = 64'h8040201008040201;
defparam \auto_autopch_req_c~2 .shared_arith = "off";

arriaii_lcell_comb \auto_autopch_req_c~3 (
	.dataa(!pipe_17_7),
	.datab(!pipe_15_7),
	.datac(!pipe_16_7),
	.datad(!\current_row[4]~q ),
	.datae(!\current_row[2]~q ),
	.dataf(!\current_row[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_autopch_req_c~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_autopch_req_c~3 .extended_lut = "off";
defparam \auto_autopch_req_c~3 .lut_mask = 64'h8040201008040201;
defparam \auto_autopch_req_c~3 .shared_arith = "off";

arriaii_lcell_comb \auto_autopch_req_c~4 (
	.dataa(!pipefull_7),
	.datab(!current_bank_0),
	.datac(!current_bank_1),
	.datad(!pipe_11_7),
	.datae(!pipe_10_7),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_autopch_req_c~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_autopch_req_c~4 .extended_lut = "off";
defparam \auto_autopch_req_c~4 .lut_mask = 64'h4004100140041001;
defparam \auto_autopch_req_c~4 .shared_arith = "off";

arriaii_lcell_comb \auto_autopch_req_c~5 (
	.dataa(!current_bank_2),
	.datab(!pipe_14_7),
	.datac(!pipe_12_7),
	.datad(!pipe_13_7),
	.datae(!\current_row[1]~q ),
	.dataf(!\current_row[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_autopch_req_c~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_autopch_req_c~5 .extended_lut = "off";
defparam \auto_autopch_req_c~5 .lut_mask = 64'h8400210000840021;
defparam \auto_autopch_req_c~5 .shared_arith = "off";

arriaii_lcell_comb \auto_autopch_req_c~6 (
	.dataa(!\auto_autopch_req_c~0_combout ),
	.datab(!\auto_autopch_req_c~1_combout ),
	.datac(!\auto_autopch_req_c~2_combout ),
	.datad(!\auto_autopch_req_c~3_combout ),
	.datae(!\auto_autopch_req_c~4_combout ),
	.dataf(!\auto_autopch_req_c~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_autopch_req_c~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_autopch_req_c~6 .extended_lut = "off";
defparam \auto_autopch_req_c~6 .lut_mask = 64'h0000000000000001;
defparam \auto_autopch_req_c~6 .shared_arith = "off";

arriaii_lcell_comb \always14~2 (
	.dataa(!current_bank_0),
	.datab(!pipefull_5),
	.datac(!pipe_10_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always14~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always14~2 .extended_lut = "off";
defparam \always14~2 .lut_mask = 64'h2121212121212121;
defparam \always14~2 .shared_arith = "off";

arriaii_lcell_comb \always14~3 (
	.dataa(!current_bank_2),
	.datab(!current_bank_1),
	.datac(!pipe_12_5),
	.datad(!pipe_11_5),
	.datae(!\always14~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always14~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always14~3 .extended_lut = "off";
defparam \always14~3 .lut_mask = 64'h0000842100008421;
defparam \always14~3 .shared_arith = "off";

arriaii_lcell_comb \always14~4 (
	.dataa(!pipefull_6),
	.datab(!current_bank_0),
	.datac(!pipe_10_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always14~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always14~4 .extended_lut = "off";
defparam \always14~4 .lut_mask = 64'h4141414141414141;
defparam \always14~4 .shared_arith = "off";

arriaii_lcell_comb \always14~5 (
	.dataa(!current_bank_2),
	.datab(!current_bank_1),
	.datac(!pipe_12_6),
	.datad(!pipe_11_6),
	.datae(!\always14~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always14~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always14~5 .extended_lut = "off";
defparam \always14~5 .lut_mask = 64'h0000842100008421;
defparam \always14~5 .shared_arith = "off";

arriaii_lcell_comb \Equal29~0 (
	.dataa(!pipe_25_5),
	.datab(!pipe_26_5),
	.datac(!\current_row[13]~q ),
	.datad(!\current_row[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal29~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal29~0 .extended_lut = "off";
defparam \Equal29~0 .lut_mask = 64'h8241824182418241;
defparam \Equal29~0 .shared_arith = "off";

arriaii_lcell_comb \Equal29~1 (
	.dataa(!pipe_24_5),
	.datab(!pipe_22_5),
	.datac(!pipe_23_5),
	.datad(!\current_row[11]~q ),
	.datae(!\current_row[10]~q ),
	.dataf(!\current_row[9]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal29~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal29~1 .extended_lut = "off";
defparam \Equal29~1 .lut_mask = 64'h8040080420100201;
defparam \Equal29~1 .shared_arith = "off";

arriaii_lcell_comb \Equal29~2 (
	.dataa(!pipe_21_5),
	.datab(!pipe_19_5),
	.datac(!pipe_20_5),
	.datad(!\current_row[8]~q ),
	.datae(!\current_row[7]~q ),
	.dataf(!\current_row[6]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal29~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal29~2 .extended_lut = "off";
defparam \Equal29~2 .lut_mask = 64'h8040080420100201;
defparam \Equal29~2 .shared_arith = "off";

arriaii_lcell_comb \Equal29~3 (
	.dataa(!pipe_15_5),
	.datab(!pipe_13_5),
	.datac(!pipe_14_5),
	.datad(!\current_row[2]~q ),
	.datae(!\current_row[1]~q ),
	.dataf(!\current_row[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal29~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal29~3 .extended_lut = "off";
defparam \Equal29~3 .lut_mask = 64'h8040080420100201;
defparam \Equal29~3 .shared_arith = "off";

arriaii_lcell_comb \Equal29~4 (
	.dataa(!pipe_18_5),
	.datab(!pipe_16_5),
	.datac(!pipe_17_5),
	.datad(!\current_row[5]~q ),
	.datae(!\current_row[4]~q ),
	.dataf(!\current_row[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal29~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal29~4 .extended_lut = "off";
defparam \Equal29~4 .lut_mask = 64'h8040080420100201;
defparam \Equal29~4 .shared_arith = "off";

arriaii_lcell_comb \Equal29~5 (
	.dataa(!\Equal29~0_combout ),
	.datab(!\Equal29~1_combout ),
	.datac(!\Equal29~2_combout ),
	.datad(!\Equal29~3_combout ),
	.datae(!\Equal29~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal29~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal29~5 .extended_lut = "off";
defparam \Equal29~5 .lut_mask = 64'h0000000100000001;
defparam \Equal29~5 .shared_arith = "off";

arriaii_lcell_comb \Equal32~0 (
	.dataa(!pipe_25_6),
	.datab(!pipe_26_6),
	.datac(!\current_row[13]~q ),
	.datad(!\current_row[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal32~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal32~0 .extended_lut = "off";
defparam \Equal32~0 .lut_mask = 64'h8241824182418241;
defparam \Equal32~0 .shared_arith = "off";

arriaii_lcell_comb \Equal32~1 (
	.dataa(!pipe_24_6),
	.datab(!pipe_22_6),
	.datac(!pipe_23_6),
	.datad(!\current_row[11]~q ),
	.datae(!\current_row[10]~q ),
	.dataf(!\current_row[9]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal32~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal32~1 .extended_lut = "off";
defparam \Equal32~1 .lut_mask = 64'h8040080420100201;
defparam \Equal32~1 .shared_arith = "off";

arriaii_lcell_comb \Equal32~2 (
	.dataa(!pipe_21_6),
	.datab(!pipe_19_6),
	.datac(!pipe_20_6),
	.datad(!\current_row[8]~q ),
	.datae(!\current_row[7]~q ),
	.dataf(!\current_row[6]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal32~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal32~2 .extended_lut = "off";
defparam \Equal32~2 .lut_mask = 64'h8040080420100201;
defparam \Equal32~2 .shared_arith = "off";

arriaii_lcell_comb \Equal32~3 (
	.dataa(!pipe_15_6),
	.datab(!pipe_13_6),
	.datac(!pipe_14_6),
	.datad(!\current_row[2]~q ),
	.datae(!\current_row[1]~q ),
	.dataf(!\current_row[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal32~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal32~3 .extended_lut = "off";
defparam \Equal32~3 .lut_mask = 64'h8040080420100201;
defparam \Equal32~3 .shared_arith = "off";

arriaii_lcell_comb \Equal32~4 (
	.dataa(!pipe_18_6),
	.datab(!pipe_16_6),
	.datac(!pipe_17_6),
	.datad(!\current_row[5]~q ),
	.datae(!\current_row[4]~q ),
	.dataf(!\current_row[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal32~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal32~4 .extended_lut = "off";
defparam \Equal32~4 .lut_mask = 64'h8040080420100201;
defparam \Equal32~4 .shared_arith = "off";

arriaii_lcell_comb \Equal32~5 (
	.dataa(!\Equal32~0_combout ),
	.datab(!\Equal32~1_combout ),
	.datac(!\Equal32~2_combout ),
	.datad(!\Equal32~3_combout ),
	.datae(!\Equal32~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal32~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal32~5 .extended_lut = "off";
defparam \Equal32~5 .lut_mask = 64'h0000000100000001;
defparam \Equal32~5 .shared_arith = "off";

arriaii_lcell_comb \auto_autopch_req_c~7 (
	.dataa(!\auto_autopch_req_c~6_combout ),
	.datab(!\always14~3_combout ),
	.datac(!\always14~5_combout ),
	.datad(!\Equal29~5_combout ),
	.datae(!\Equal32~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_autopch_req_c~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_autopch_req_c~7 .extended_lut = "off";
defparam \auto_autopch_req_c~7 .lut_mask = 64'hBF8CB380BF8CB380;
defparam \auto_autopch_req_c~7 .shared_arith = "off";

arriaii_lcell_comb \always14~6 (
	.dataa(!pipefull_3),
	.datab(!\Equal12~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always14~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always14~6 .extended_lut = "off";
defparam \always14~6 .lut_mask = 64'h1111111111111111;
defparam \always14~6 .shared_arith = "off";

arriaii_lcell_comb \Equal22~0 (
	.dataa(!\current_row[13]~q ),
	.datab(!\current_row[12]~q ),
	.datac(!pipe_25_2),
	.datad(!pipe_26_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal22~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal22~0 .extended_lut = "off";
defparam \Equal22~0 .lut_mask = 64'h8241824182418241;
defparam \Equal22~0 .shared_arith = "off";

arriaii_lcell_comb \Equal20~0 (
	.dataa(!pipe_25_0),
	.datab(!pipe_26_0),
	.datac(!\current_row[13]~q ),
	.datad(!\current_row[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal20~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal20~0 .extended_lut = "off";
defparam \Equal20~0 .lut_mask = 64'h8241824182418241;
defparam \Equal20~0 .shared_arith = "off";

arriaii_lcell_comb \Equal21~0 (
	.dataa(!\current_row[13]~q ),
	.datab(!\current_row[12]~q ),
	.datac(!pipe_25_1),
	.datad(!pipe_26_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal21~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal21~0 .extended_lut = "off";
defparam \Equal21~0 .lut_mask = 64'h8241824182418241;
defparam \Equal21~0 .shared_arith = "off";

arriaii_lcell_comb \Equal23~1 (
	.dataa(!pipe_24_3),
	.datab(!pipe_22_3),
	.datac(!pipe_23_3),
	.datad(!\current_row[11]~q ),
	.datae(!\current_row[10]~q ),
	.dataf(!\current_row[9]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal23~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal23~1 .extended_lut = "off";
defparam \Equal23~1 .lut_mask = 64'h8040080420100201;
defparam \Equal23~1 .shared_arith = "off";

dffeas do_read_r(
	.clk(ctl_clk),
	.d(\current_read~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(!\state.READWRITE~q ),
	.sload(gnd),
	.ena(vcc),
	.q(do_read_r1),
	.prn(vcc));
defparam do_read_r.is_wysiwyg = "true";
defparam do_read_r.power_up = "low";

dffeas do_auto_precharge_r(
	.clk(ctl_clk),
	.d(\do_auto_precharge~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(!\state.READWRITE~q ),
	.sload(gnd),
	.ena(vcc),
	.q(do_auto_precharge_r1),
	.prn(vcc));
defparam do_auto_precharge_r.is_wysiwyg = "true";
defparam do_auto_precharge_r.power_up = "low";

dffeas do_write_r(
	.clk(ctl_clk),
	.d(\current_read~_wirecell_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(!\state.READWRITE~q ),
	.sload(gnd),
	.ena(vcc),
	.q(do_write_r1),
	.prn(vcc));
defparam do_write_r.is_wysiwyg = "true";
defparam do_write_r.power_up = "low";

dffeas do_burst_chop_r(
	.clk(ctl_clk),
	.d(\always39~3_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(!\state.READWRITE~q ),
	.sload(gnd),
	.ena(vcc),
	.q(do_burst_chop_r1),
	.prn(vcc));
defparam do_burst_chop_r.is_wysiwyg = "true";
defparam do_burst_chop_r.power_up = "low";

dffeas \to_row_addr_r[0] (
	.clk(ctl_clk),
	.d(\Selector39~0_combout ),
	.asdata(\current_row[0]~q ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\to_row_addr_r[5]~2_combout ),
	.sload(\to_bank_addr_r[2]~1_combout ),
	.ena(vcc),
	.q(to_row_addr_r_0),
	.prn(vcc));
defparam \to_row_addr_r[0] .is_wysiwyg = "true";
defparam \to_row_addr_r[0] .power_up = "low";

dffeas \to_row_addr_r[1] (
	.clk(ctl_clk),
	.d(\Selector38~0_combout ),
	.asdata(\current_row[1]~q ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\to_row_addr_r[5]~2_combout ),
	.sload(\to_bank_addr_r[2]~1_combout ),
	.ena(vcc),
	.q(to_row_addr_r_1),
	.prn(vcc));
defparam \to_row_addr_r[1] .is_wysiwyg = "true";
defparam \to_row_addr_r[1] .power_up = "low";

dffeas \to_col_addr_r[2] (
	.clk(ctl_clk),
	.d(\to_addr~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(!\state.READWRITE~q ),
	.sload(gnd),
	.ena(vcc),
	.q(to_col_addr_r_2),
	.prn(vcc));
defparam \to_col_addr_r[2] .is_wysiwyg = "true";
defparam \to_col_addr_r[2] .power_up = "low";

dffeas \to_row_addr_r[2] (
	.clk(ctl_clk),
	.d(\Selector37~0_combout ),
	.asdata(\current_row[2]~q ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\to_row_addr_r[5]~2_combout ),
	.sload(\to_bank_addr_r[2]~1_combout ),
	.ena(vcc),
	.q(to_row_addr_r_2),
	.prn(vcc));
defparam \to_row_addr_r[2] .is_wysiwyg = "true";
defparam \to_row_addr_r[2] .power_up = "low";

dffeas \to_col_addr_r[3] (
	.clk(ctl_clk),
	.d(\current_col[3]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(!\state.READWRITE~q ),
	.sload(gnd),
	.ena(vcc),
	.q(to_col_addr_r_3),
	.prn(vcc));
defparam \to_col_addr_r[3] .is_wysiwyg = "true";
defparam \to_col_addr_r[3] .power_up = "low";

dffeas \to_row_addr_r[3] (
	.clk(ctl_clk),
	.d(\Selector36~0_combout ),
	.asdata(\current_row[3]~q ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\to_row_addr_r[5]~2_combout ),
	.sload(\to_bank_addr_r[2]~1_combout ),
	.ena(vcc),
	.q(to_row_addr_r_3),
	.prn(vcc));
defparam \to_row_addr_r[3] .is_wysiwyg = "true";
defparam \to_row_addr_r[3] .power_up = "low";

dffeas \to_col_addr_r[4] (
	.clk(ctl_clk),
	.d(\current_col[4]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(!\state.READWRITE~q ),
	.sload(gnd),
	.ena(vcc),
	.q(to_col_addr_r_4),
	.prn(vcc));
defparam \to_col_addr_r[4] .is_wysiwyg = "true";
defparam \to_col_addr_r[4] .power_up = "low";

dffeas \to_row_addr_r[4] (
	.clk(ctl_clk),
	.d(\Selector35~0_combout ),
	.asdata(\current_row[4]~q ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\to_row_addr_r[5]~2_combout ),
	.sload(\to_bank_addr_r[2]~1_combout ),
	.ena(vcc),
	.q(to_row_addr_r_4),
	.prn(vcc));
defparam \to_row_addr_r[4] .is_wysiwyg = "true";
defparam \to_row_addr_r[4] .power_up = "low";

dffeas \to_col_addr_r[5] (
	.clk(ctl_clk),
	.d(\current_col[5]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(!\state.READWRITE~q ),
	.sload(gnd),
	.ena(vcc),
	.q(to_col_addr_r_5),
	.prn(vcc));
defparam \to_col_addr_r[5] .is_wysiwyg = "true";
defparam \to_col_addr_r[5] .power_up = "low";

dffeas \to_row_addr_r[5] (
	.clk(ctl_clk),
	.d(\Selector34~0_combout ),
	.asdata(\current_row[5]~q ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\to_row_addr_r[5]~2_combout ),
	.sload(\to_bank_addr_r[2]~1_combout ),
	.ena(vcc),
	.q(to_row_addr_r_5),
	.prn(vcc));
defparam \to_row_addr_r[5] .is_wysiwyg = "true";
defparam \to_row_addr_r[5] .power_up = "low";

dffeas \to_col_addr_r[6] (
	.clk(ctl_clk),
	.d(\current_col[6]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(!\state.READWRITE~q ),
	.sload(gnd),
	.ena(vcc),
	.q(to_col_addr_r_6),
	.prn(vcc));
defparam \to_col_addr_r[6] .is_wysiwyg = "true";
defparam \to_col_addr_r[6] .power_up = "low";

dffeas \to_row_addr_r[6] (
	.clk(ctl_clk),
	.d(\Selector33~0_combout ),
	.asdata(\current_row[6]~q ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\to_row_addr_r[5]~2_combout ),
	.sload(\to_bank_addr_r[2]~1_combout ),
	.ena(vcc),
	.q(to_row_addr_r_6),
	.prn(vcc));
defparam \to_row_addr_r[6] .is_wysiwyg = "true";
defparam \to_row_addr_r[6] .power_up = "low";

dffeas \to_col_addr_r[7] (
	.clk(ctl_clk),
	.d(\current_col[7]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(!\state.READWRITE~q ),
	.sload(gnd),
	.ena(vcc),
	.q(to_col_addr_r_7),
	.prn(vcc));
defparam \to_col_addr_r[7] .is_wysiwyg = "true";
defparam \to_col_addr_r[7] .power_up = "low";

dffeas \to_row_addr_r[7] (
	.clk(ctl_clk),
	.d(\Selector32~0_combout ),
	.asdata(\current_row[7]~q ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\to_row_addr_r[5]~2_combout ),
	.sload(\to_bank_addr_r[2]~1_combout ),
	.ena(vcc),
	.q(to_row_addr_r_7),
	.prn(vcc));
defparam \to_row_addr_r[7] .is_wysiwyg = "true";
defparam \to_row_addr_r[7] .power_up = "low";

dffeas \to_col_addr_r[8] (
	.clk(ctl_clk),
	.d(\current_col[8]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(!\state.READWRITE~q ),
	.sload(gnd),
	.ena(vcc),
	.q(to_col_addr_r_8),
	.prn(vcc));
defparam \to_col_addr_r[8] .is_wysiwyg = "true";
defparam \to_col_addr_r[8] .power_up = "low";

dffeas \to_row_addr_r[8] (
	.clk(ctl_clk),
	.d(\Selector31~0_combout ),
	.asdata(\current_row[8]~q ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\to_row_addr_r[5]~2_combout ),
	.sload(\to_bank_addr_r[2]~1_combout ),
	.ena(vcc),
	.q(to_row_addr_r_8),
	.prn(vcc));
defparam \to_row_addr_r[8] .is_wysiwyg = "true";
defparam \to_row_addr_r[8] .power_up = "low";

dffeas \to_col_addr_r[9] (
	.clk(ctl_clk),
	.d(\current_col[9]~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(!\state.READWRITE~q ),
	.sload(gnd),
	.ena(vcc),
	.q(to_col_addr_r_9),
	.prn(vcc));
defparam \to_col_addr_r[9] .is_wysiwyg = "true";
defparam \to_col_addr_r[9] .power_up = "low";

dffeas \to_row_addr_r[9] (
	.clk(ctl_clk),
	.d(\Selector30~0_combout ),
	.asdata(\current_row[9]~q ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\to_row_addr_r[5]~2_combout ),
	.sload(\to_bank_addr_r[2]~1_combout ),
	.ena(vcc),
	.q(to_row_addr_r_9),
	.prn(vcc));
defparam \to_row_addr_r[9] .is_wysiwyg = "true";
defparam \to_row_addr_r[9] .power_up = "low";

dffeas \to_row_addr_r[10] (
	.clk(ctl_clk),
	.d(\Selector29~0_combout ),
	.asdata(\current_row[10]~q ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\to_row_addr_r[5]~2_combout ),
	.sload(\to_bank_addr_r[2]~1_combout ),
	.ena(vcc),
	.q(to_row_addr_r_10),
	.prn(vcc));
defparam \to_row_addr_r[10] .is_wysiwyg = "true";
defparam \to_row_addr_r[10] .power_up = "low";

dffeas \to_row_addr_r[11] (
	.clk(ctl_clk),
	.d(\Selector28~0_combout ),
	.asdata(\current_row[11]~q ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\to_row_addr_r[5]~2_combout ),
	.sload(\to_bank_addr_r[2]~1_combout ),
	.ena(vcc),
	.q(to_row_addr_r_11),
	.prn(vcc));
defparam \to_row_addr_r[11] .is_wysiwyg = "true";
defparam \to_row_addr_r[11] .power_up = "low";

dffeas \to_row_addr_r[12] (
	.clk(ctl_clk),
	.d(\Selector27~0_combout ),
	.asdata(\current_row[12]~q ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\to_row_addr_r[5]~2_combout ),
	.sload(\to_bank_addr_r[2]~1_combout ),
	.ena(vcc),
	.q(to_row_addr_r_12),
	.prn(vcc));
defparam \to_row_addr_r[12] .is_wysiwyg = "true";
defparam \to_row_addr_r[12] .power_up = "low";

dffeas \to_row_addr_r[13] (
	.clk(ctl_clk),
	.d(\Selector26~0_combout ),
	.asdata(\current_row[13]~q ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(\to_row_addr_r[5]~2_combout ),
	.sload(\to_bank_addr_r[2]~1_combout ),
	.ena(vcc),
	.q(to_row_addr_r_13),
	.prn(vcc));
defparam \to_row_addr_r[13] .is_wysiwyg = "true";
defparam \to_row_addr_r[13] .power_up = "low";

dffeas int_refresh_ack(
	.clk(ctl_clk),
	.d(\Selector10~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(int_refresh_ack1),
	.prn(vcc));
defparam int_refresh_ack.is_wysiwyg = "true";
defparam int_refresh_ack.power_up = "low";

dffeas fetch(
	.clk(ctl_clk),
	.d(\Selector11~2_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(fetch1),
	.prn(vcc));
defparam fetch.is_wysiwyg = "true";
defparam fetch.power_up = "low";

dffeas do_precharge_all_r(
	.clk(ctl_clk),
	.d(\do_precharge_all~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(do_precharge_all_r1),
	.prn(vcc));
defparam do_precharge_all_r.is_wysiwyg = "true";
defparam do_precharge_all_r.power_up = "low";

arriaii_lcell_comb \always38~0 (
	.dataa(!read_req),
	.datab(!write_req),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always38),
	.sumout(),
	.cout(),
	.shareout());
defparam \always38~0 .extended_lut = "off";
defparam \always38~0 .lut_mask = 64'h8888888888888888;
defparam \always38~0 .shared_arith = "off";

dffeas do_refresh_r(
	.clk(ctl_clk),
	.d(\Selector10~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(do_refresh_r1),
	.prn(vcc));
defparam do_refresh_r.is_wysiwyg = "true";
defparam do_refresh_r.power_up = "low";

dffeas \to_chip_r[0] (
	.clk(ctl_clk),
	.d(\Selector22~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(to_chip_r_0),
	.prn(vcc));
defparam \to_chip_r[0] .is_wysiwyg = "true";
defparam \to_chip_r[0] .power_up = "low";

arriaii_lcell_comb \always38~3 (
	.dataa(!to_chip_r_0),
	.datab(!do_auto_precharge_r1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always381),
	.sumout(),
	.cout(),
	.shareout());
defparam \always38~3 .extended_lut = "off";
defparam \always38~3 .lut_mask = 64'h1111111111111111;
defparam \always38~3 .shared_arith = "off";

dffeas \to_bank_addr_r[2] (
	.clk(ctl_clk),
	.d(\Selector23~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(to_bank_addr_r_2),
	.prn(vcc));
defparam \to_bank_addr_r[2] .is_wysiwyg = "true";
defparam \to_bank_addr_r[2] .power_up = "low";

dffeas \current_bank[2] (
	.clk(ctl_clk),
	.d(pipe_12_0),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fetch1),
	.q(current_bank_2),
	.prn(vcc));
defparam \current_bank[2] .is_wysiwyg = "true";
defparam \current_bank[2] .power_up = "low";

dffeas \to_bank_addr_r[0] (
	.clk(ctl_clk),
	.d(\Selector25~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(to_bank_addr_r_0),
	.prn(vcc));
defparam \to_bank_addr_r[0] .is_wysiwyg = "true";
defparam \to_bank_addr_r[0] .power_up = "low";

dffeas \current_bank[0] (
	.clk(ctl_clk),
	.d(pipe_10_0),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fetch1),
	.q(current_bank_0),
	.prn(vcc));
defparam \current_bank[0] .is_wysiwyg = "true";
defparam \current_bank[0] .power_up = "low";

dffeas \to_bank_addr_r[1] (
	.clk(ctl_clk),
	.d(\Selector24~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(to_bank_addr_r_1),
	.prn(vcc));
defparam \to_bank_addr_r[1] .is_wysiwyg = "true";
defparam \to_bank_addr_r[1] .power_up = "low";

dffeas \current_bank[1] (
	.clk(ctl_clk),
	.d(pipe_11_0),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fetch1),
	.q(current_bank_1),
	.prn(vcc));
defparam \current_bank[1] .is_wysiwyg = "true";
defparam \current_bank[1] .power_up = "low";

arriaii_lcell_comb \always38~4 (
	.dataa(!to_bank_addr_r_2),
	.datab(!current_bank_2),
	.datac(!to_bank_addr_r_0),
	.datad(!current_bank_0),
	.datae(!to_bank_addr_r_1),
	.dataf(!current_bank_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always382),
	.sumout(),
	.cout(),
	.shareout());
defparam \always38~4 .extended_lut = "off";
defparam \always38~4 .lut_mask = 64'h9009000000009009;
defparam \always38~4 .shared_arith = "off";

dffeas rdwr_data_valid_r(
	.clk(ctl_clk),
	.d(\new_gen_rdwr_data_valid~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rdwr_data_valid_r1),
	.prn(vcc));
defparam rdwr_data_valid_r.is_wysiwyg = "true";
defparam rdwr_data_valid_r.power_up = "low";

dffeas do_activate_r(
	.clk(ctl_clk),
	.d(\Selector20~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(do_activate_r1),
	.prn(vcc));
defparam do_activate_r.is_wysiwyg = "true";
defparam do_activate_r.power_up = "low";

dffeas current_read(
	.clk(ctl_clk),
	.d(pipe_33_0),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fetch1),
	.q(\current_read~q ),
	.prn(vcc));
defparam current_read.is_wysiwyg = "true";
defparam current_read.power_up = "low";

arriaii_lcell_comb \always38~5 (
	.dataa(!out_cmd_info_valid_0),
	.datab(!out_cmd_bank_is_open_0),
	.datac(!always381),
	.datad(!always382),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always38~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always38~5 .extended_lut = "off";
defparam \always38~5 .lut_mask = 64'h1110111011101110;
defparam \always38~5 .shared_arith = "off";

arriaii_lcell_comb \always38~6 (
	.dataa(!\current_write~q ),
	.datab(!do_read_r1),
	.datac(!out_cmd_can_write_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always38~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always38~6 .extended_lut = "off";
defparam \always38~6 .lut_mask = 64'h0404040404040404;
defparam \always38~6 .shared_arith = "off";

dffeas \current_burstcount_counter_temp[0] (
	.clk(ctl_clk),
	.d(pipe_28_0),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fetch1),
	.q(\current_burstcount_counter_temp[0]~q ),
	.prn(vcc));
defparam \current_burstcount_counter_temp[0] .is_wysiwyg = "true";
defparam \current_burstcount_counter_temp[0] .power_up = "low";

arriaii_lcell_comb \Selector19~0 (
	.dataa(!\state.DO2~q ),
	.datab(!\start_burst~q ),
	.datac(!\always38~15_combout ),
	.datad(!\state.READWRITE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector19~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector19~0 .extended_lut = "off";
defparam \Selector19~0 .lut_mask = 64'h3715371537153715;
defparam \Selector19~0 .shared_arith = "off";

dffeas start_burst(
	.clk(ctl_clk),
	.d(\Selector19~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\start_burst~q ),
	.prn(vcc));
defparam start_burst.is_wysiwyg = "true";
defparam start_burst.power_up = "low";

dffeas start_burst_r(
	.clk(ctl_clk),
	.d(\start_burst~q ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\start_burst_r~q ),
	.prn(vcc));
defparam start_burst_r.is_wysiwyg = "true";
defparam start_burst_r.power_up = "low";

dffeas \current_col[2] (
	.clk(ctl_clk),
	.d(pipe_2_0),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fetch1),
	.q(\current_col[2]~q ),
	.prn(vcc));
defparam \current_col[2] .is_wysiwyg = "true";
defparam \current_col[2] .power_up = "low";

arriaii_lcell_comb \burst_delay~0 (
	.dataa(!\fetch_r~q ),
	.datab(!\start_burst~q ),
	.datac(!\start_burst_r~q ),
	.datad(!\burst_delay~q ),
	.datae(!\current_col[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\burst_delay~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \burst_delay~0 .extended_lut = "off";
defparam \burst_delay~0 .lut_mask = 64'h008055D5008055D5;
defparam \burst_delay~0 .shared_arith = "off";

dffeas burst_delay(
	.clk(ctl_clk),
	.d(\burst_delay~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\burst_delay~q ),
	.prn(vcc));
defparam burst_delay.is_wysiwyg = "true";
defparam burst_delay.power_up = "low";

arriaii_lcell_comb \always29~0 (
	.dataa(!\current_burstcount_counter[1]~q ),
	.datab(!\current_burstcount_counter[0]~q ),
	.datac(!\start_burst~q ),
	.datad(!\start_burst_r~q ),
	.datae(!\burst_delay~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always29~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always29~0 .extended_lut = "off";
defparam \always29~0 .lut_mask = 64'h0777000007770000;
defparam \always29~0 .shared_arith = "off";

arriaii_lcell_comb \current_burstcount_counter[0]~0 (
	.dataa(!\fetch_r~q ),
	.datab(!\current_burstcount_counter[0]~q ),
	.datac(!\current_burstcount_counter_temp[0]~q ),
	.datad(!\always29~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\current_burstcount_counter[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \current_burstcount_counter[0]~0 .extended_lut = "off";
defparam \current_burstcount_counter[0]~0 .lut_mask = 64'h278D278D278D278D;
defparam \current_burstcount_counter[0]~0 .shared_arith = "off";

dffeas \current_burstcount_counter[0] (
	.clk(ctl_clk),
	.d(\current_burstcount_counter[0]~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\current_burstcount_counter[0]~q ),
	.prn(vcc));
defparam \current_burstcount_counter[0] .is_wysiwyg = "true";
defparam \current_burstcount_counter[0] .power_up = "low";

arriaii_lcell_comb \write_burst_length~0 (
	.dataa(!\current_write~q ),
	.datab(!\start_burst~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write_burst_length~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_burst_length~0 .extended_lut = "off";
defparam \write_burst_length~0 .lut_mask = 64'h1111111111111111;
defparam \write_burst_length~0 .shared_arith = "off";

dffeas start_write_burst_r(
	.clk(ctl_clk),
	.d(\write_burst_length~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\start_write_burst_r~q ),
	.prn(vcc));
defparam start_write_burst_r.is_wysiwyg = "true";
defparam start_write_burst_r.power_up = "low";

dffeas current_write(
	.clk(ctl_clk),
	.d(pipe_32_0),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fetch1),
	.q(\current_write~q ),
	.prn(vcc));
defparam current_write.is_wysiwyg = "true";
defparam current_write.power_up = "low";

arriaii_lcell_comb \always17~0 (
	.dataa(!\current_burstcount_counter[1]~q ),
	.datab(!\current_burstcount_counter[0]~q ),
	.datac(!\start_write_burst_r~q ),
	.datad(!\burst_delay~q ),
	.datae(!\current_write~q ),
	.dataf(!\start_burst~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always17~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always17~0 .extended_lut = "off";
defparam \always17~0 .lut_mask = 64'hF8FFF8FFF8FF88FF;
defparam \always17~0 .shared_arith = "off";

arriaii_lcell_comb \Add0~2 (
	.dataa(!internal_ready),
	.datab(!hold_ready),
	.datac(!local_write_req),
	.datad(!\always17~0_combout ),
	.datae(gnd),
	.dataf(!\proper_beats_in_fifo[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~2_sumout ),
	.cout(\Add0~3 ),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h0000FF000000FBFF;
defparam \Add0~2 .shared_arith = "off";

arriaii_lcell_comb \proper_beats_in_fifo[9]~0 (
	.dataa(!avalon_write_req),
	.datab(!\always17~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\proper_beats_in_fifo[9]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \proper_beats_in_fifo[9]~0 .extended_lut = "off";
defparam \proper_beats_in_fifo[9]~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \proper_beats_in_fifo[9]~0 .shared_arith = "off";

dffeas \proper_beats_in_fifo[0] (
	.clk(ctl_clk),
	.d(\Add0~2_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\proper_beats_in_fifo[9]~0_combout ),
	.q(\proper_beats_in_fifo[0]~q ),
	.prn(vcc));
defparam \proper_beats_in_fifo[0] .is_wysiwyg = "true";
defparam \proper_beats_in_fifo[0] .power_up = "low";

arriaii_lcell_comb \Add0~6 (
	.dataa(!internal_ready),
	.datab(!hold_ready),
	.datac(gnd),
	.datad(!\proper_beats_in_fifo[1]~q ),
	.datae(gnd),
	.dataf(!local_write_req),
	.datag(gnd),
	.cin(\Add0~3 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~6_sumout ),
	.cout(\Add0~7 ),
	.shareout());
defparam \Add0~6 .extended_lut = "off";
defparam \Add0~6 .lut_mask = 64'h00000044000000FF;
defparam \Add0~6 .shared_arith = "off";

dffeas \proper_beats_in_fifo[1] (
	.clk(ctl_clk),
	.d(\Add0~6_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\proper_beats_in_fifo[9]~0_combout ),
	.q(\proper_beats_in_fifo[1]~q ),
	.prn(vcc));
defparam \proper_beats_in_fifo[1] .is_wysiwyg = "true";
defparam \proper_beats_in_fifo[1] .power_up = "low";

arriaii_lcell_comb \always38~8 (
	.dataa(!\current_write~q ),
	.datab(!\proper_beats_in_fifo[1]~q ),
	.datac(!\proper_beats_in_fifo[0]~q ),
	.datad(!\start_write_burst_r~q ),
	.datae(!\start_burst~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always38~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always38~8 .extended_lut = "off";
defparam \always38~8 .lut_mask = 64'h3303230333032303;
defparam \always38~8 .shared_arith = "off";

arriaii_lcell_comb \Add0~10 (
	.dataa(!local_write_req),
	.datab(!hold_ready),
	.datac(gnd),
	.datad(!\proper_beats_in_fifo[2]~q ),
	.datae(gnd),
	.dataf(!internal_ready),
	.datag(gnd),
	.cin(\Add0~7 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~10_sumout ),
	.cout(\Add0~11 ),
	.shareout());
defparam \Add0~10 .extended_lut = "off";
defparam \Add0~10 .lut_mask = 64'h00000044000000FF;
defparam \Add0~10 .shared_arith = "off";

dffeas \proper_beats_in_fifo[2] (
	.clk(ctl_clk),
	.d(\Add0~10_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\proper_beats_in_fifo[9]~0_combout ),
	.q(\proper_beats_in_fifo[2]~q ),
	.prn(vcc));
defparam \proper_beats_in_fifo[2] .is_wysiwyg = "true";
defparam \proper_beats_in_fifo[2] .power_up = "low";

arriaii_lcell_comb \Add0~14 (
	.dataa(!local_write_req),
	.datab(!hold_ready),
	.datac(gnd),
	.datad(!\proper_beats_in_fifo[3]~q ),
	.datae(gnd),
	.dataf(!internal_ready),
	.datag(gnd),
	.cin(\Add0~11 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~14_sumout ),
	.cout(\Add0~15 ),
	.shareout());
defparam \Add0~14 .extended_lut = "off";
defparam \Add0~14 .lut_mask = 64'h00000044000000FF;
defparam \Add0~14 .shared_arith = "off";

dffeas \proper_beats_in_fifo[3] (
	.clk(ctl_clk),
	.d(\Add0~14_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\proper_beats_in_fifo[9]~0_combout ),
	.q(\proper_beats_in_fifo[3]~q ),
	.prn(vcc));
defparam \proper_beats_in_fifo[3] .is_wysiwyg = "true";
defparam \proper_beats_in_fifo[3] .power_up = "low";

arriaii_lcell_comb \Add0~18 (
	.dataa(!local_write_req),
	.datab(!hold_ready),
	.datac(gnd),
	.datad(!\proper_beats_in_fifo[4]~q ),
	.datae(gnd),
	.dataf(!internal_ready),
	.datag(gnd),
	.cin(\Add0~15 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~18_sumout ),
	.cout(\Add0~19 ),
	.shareout());
defparam \Add0~18 .extended_lut = "off";
defparam \Add0~18 .lut_mask = 64'h00000044000000FF;
defparam \Add0~18 .shared_arith = "off";

dffeas \proper_beats_in_fifo[4] (
	.clk(ctl_clk),
	.d(\Add0~18_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\proper_beats_in_fifo[9]~0_combout ),
	.q(\proper_beats_in_fifo[4]~q ),
	.prn(vcc));
defparam \proper_beats_in_fifo[4] .is_wysiwyg = "true";
defparam \proper_beats_in_fifo[4] .power_up = "low";

arriaii_lcell_comb \Add0~22 (
	.dataa(!local_write_req),
	.datab(!hold_ready),
	.datac(gnd),
	.datad(!\proper_beats_in_fifo[5]~q ),
	.datae(gnd),
	.dataf(!internal_ready),
	.datag(gnd),
	.cin(\Add0~19 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~22_sumout ),
	.cout(\Add0~23 ),
	.shareout());
defparam \Add0~22 .extended_lut = "off";
defparam \Add0~22 .lut_mask = 64'h00000044000000FF;
defparam \Add0~22 .shared_arith = "off";

dffeas \proper_beats_in_fifo[5] (
	.clk(ctl_clk),
	.d(\Add0~22_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\proper_beats_in_fifo[9]~0_combout ),
	.q(\proper_beats_in_fifo[5]~q ),
	.prn(vcc));
defparam \proper_beats_in_fifo[5] .is_wysiwyg = "true";
defparam \proper_beats_in_fifo[5] .power_up = "low";

arriaii_lcell_comb \Add0~26 (
	.dataa(!local_write_req),
	.datab(!hold_ready),
	.datac(gnd),
	.datad(!\proper_beats_in_fifo[6]~q ),
	.datae(gnd),
	.dataf(!internal_ready),
	.datag(gnd),
	.cin(\Add0~23 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~26_sumout ),
	.cout(\Add0~27 ),
	.shareout());
defparam \Add0~26 .extended_lut = "off";
defparam \Add0~26 .lut_mask = 64'h00000044000000FF;
defparam \Add0~26 .shared_arith = "off";

dffeas \proper_beats_in_fifo[6] (
	.clk(ctl_clk),
	.d(\Add0~26_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\proper_beats_in_fifo[9]~0_combout ),
	.q(\proper_beats_in_fifo[6]~q ),
	.prn(vcc));
defparam \proper_beats_in_fifo[6] .is_wysiwyg = "true";
defparam \proper_beats_in_fifo[6] .power_up = "low";

arriaii_lcell_comb \Add0~30 (
	.dataa(!local_write_req),
	.datab(!hold_ready),
	.datac(gnd),
	.datad(!\proper_beats_in_fifo[7]~q ),
	.datae(gnd),
	.dataf(!internal_ready),
	.datag(gnd),
	.cin(\Add0~27 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~30_sumout ),
	.cout(\Add0~31 ),
	.shareout());
defparam \Add0~30 .extended_lut = "off";
defparam \Add0~30 .lut_mask = 64'h00000044000000FF;
defparam \Add0~30 .shared_arith = "off";

dffeas \proper_beats_in_fifo[7] (
	.clk(ctl_clk),
	.d(\Add0~30_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\proper_beats_in_fifo[9]~0_combout ),
	.q(\proper_beats_in_fifo[7]~q ),
	.prn(vcc));
defparam \proper_beats_in_fifo[7] .is_wysiwyg = "true";
defparam \proper_beats_in_fifo[7] .power_up = "low";

arriaii_lcell_comb \Add0~34 (
	.dataa(!local_write_req),
	.datab(!hold_ready),
	.datac(gnd),
	.datad(!\proper_beats_in_fifo[8]~q ),
	.datae(gnd),
	.dataf(!internal_ready),
	.datag(gnd),
	.cin(\Add0~31 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~34_sumout ),
	.cout(\Add0~35 ),
	.shareout());
defparam \Add0~34 .extended_lut = "off";
defparam \Add0~34 .lut_mask = 64'h00000044000000FF;
defparam \Add0~34 .shared_arith = "off";

dffeas \proper_beats_in_fifo[8] (
	.clk(ctl_clk),
	.d(\Add0~34_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\proper_beats_in_fifo[9]~0_combout ),
	.q(\proper_beats_in_fifo[8]~q ),
	.prn(vcc));
defparam \proper_beats_in_fifo[8] .is_wysiwyg = "true";
defparam \proper_beats_in_fifo[8] .power_up = "low";

arriaii_lcell_comb \Add0~38 (
	.dataa(!local_write_req),
	.datab(!hold_ready),
	.datac(gnd),
	.datad(!\proper_beats_in_fifo[9]~q ),
	.datae(gnd),
	.dataf(!internal_ready),
	.datag(gnd),
	.cin(\Add0~35 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~38_sumout ),
	.cout(),
	.shareout());
defparam \Add0~38 .extended_lut = "off";
defparam \Add0~38 .lut_mask = 64'h00000044000000FF;
defparam \Add0~38 .shared_arith = "off";

dffeas \proper_beats_in_fifo[9] (
	.clk(ctl_clk),
	.d(\Add0~38_sumout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\proper_beats_in_fifo[9]~0_combout ),
	.q(\proper_beats_in_fifo[9]~q ),
	.prn(vcc));
defparam \proper_beats_in_fifo[9] .is_wysiwyg = "true";
defparam \proper_beats_in_fifo[9] .power_up = "low";

arriaii_lcell_comb \always38~9 (
	.dataa(!\proper_beats_in_fifo[5]~q ),
	.datab(!\proper_beats_in_fifo[6]~q ),
	.datac(!\proper_beats_in_fifo[7]~q ),
	.datad(!\proper_beats_in_fifo[9]~q ),
	.datae(!\proper_beats_in_fifo[8]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always38~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always38~9 .extended_lut = "off";
defparam \always38~9 .lut_mask = 64'h8000000080000000;
defparam \always38~9 .shared_arith = "off";

dffeas \current_burstcount_counter_temp[1] (
	.clk(ctl_clk),
	.d(pipe_29_0),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fetch1),
	.q(\current_burstcount_counter_temp[1]~q ),
	.prn(vcc));
defparam \current_burstcount_counter_temp[1] .is_wysiwyg = "true";
defparam \current_burstcount_counter_temp[1] .power_up = "low";

arriaii_lcell_comb \always38~10 (
	.dataa(!\fetch_r~q ),
	.datab(!\current_burstcount_counter_temp[1]~q ),
	.datac(!\current_burstcount_counter_temp[0]~q ),
	.datad(!\proper_beats_in_fifo[3]~q ),
	.datae(!\proper_beats_in_fifo[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always38~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always38~10 .extended_lut = "off";
defparam \always38~10 .lut_mask = 64'hFB000000FB000000;
defparam \always38~10 .shared_arith = "off";

arriaii_lcell_comb \always38~11 (
	.dataa(!\always38~7_combout ),
	.datab(!\always38~8_combout ),
	.datac(!\proper_beats_in_fifo[4]~q ),
	.datad(!\always38~9_combout ),
	.datae(!\always38~10_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always38~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always38~11 .extended_lut = "off";
defparam \always38~11 .lut_mask = 64'h0000008000000080;
defparam \always38~11 .shared_arith = "off";

arriaii_lcell_comb \always38~1 (
	.dataa(!out_cmd_info_valid_0),
	.datab(!\just_did_activate~q ),
	.datac(!out_cmd_can_activate_0),
	.datad(!out_cmd_bank_is_open_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always38~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always38~1 .extended_lut = "off";
defparam \always38~1 .lut_mask = 64'h0400040004000400;
defparam \always38~1 .shared_arith = "off";

arriaii_lcell_comb \Selector20~0 (
	.dataa(!add_lat_on),
	.datab(!\always38~1_combout ),
	.datac(!can_al_activate_write),
	.datad(!can_al_activate_read),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector20~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector20~0 .extended_lut = "off";
defparam \Selector20~0 .lut_mask = 64'h2333233323332333;
defparam \Selector20~0 .shared_arith = "off";

arriaii_lcell_comb \always14~0 (
	.dataa(!current_bank_0),
	.datab(!current_bank_1),
	.datac(!pipe_10_1),
	.datad(!pipe_11_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always14~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always14~0 .extended_lut = "off";
defparam \always14~0 .lut_mask = 64'h8421842184218421;
defparam \always14~0 .shared_arith = "off";

arriaii_lcell_comb \Equal4~0 (
	.dataa(!pipe_10_0),
	.datab(!pipe_12_0),
	.datac(!pipe_11_0),
	.datad(!pipe_12_1),
	.datae(!pipe_10_1),
	.dataf(!pipe_11_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~0 .extended_lut = "off";
defparam \Equal4~0 .lut_mask = 64'h8020401008020401;
defparam \Equal4~0 .shared_arith = "off";

arriaii_lcell_comb \always11~0 (
	.dataa(!current_bank_2),
	.datab(!pipefull_1),
	.datac(!pipe_12_1),
	.datad(!\always14~0_combout ),
	.datae(!\Equal4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always11~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always11~0 .extended_lut = "off";
defparam \always11~0 .lut_mask = 64'h3312000033120000;
defparam \always11~0 .shared_arith = "off";

arriaii_lcell_comb \always12~0 (
	.dataa(!pipe_10_2),
	.datab(!pipe_10_1),
	.datac(!pipe_11_2),
	.datad(!pipe_11_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always12~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always12~0 .extended_lut = "off";
defparam \always12~0 .lut_mask = 64'h9009900990099009;
defparam \always12~0 .shared_arith = "off";

arriaii_lcell_comb \Equal8~0 (
	.dataa(!pipe_10_0),
	.datab(!pipe_12_0),
	.datac(!pipe_11_0),
	.datad(!pipe_12_2),
	.datae(!pipe_10_2),
	.dataf(!pipe_11_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal8~0 .extended_lut = "off";
defparam \Equal8~0 .lut_mask = 64'h8020401008020401;
defparam \Equal8~0 .shared_arith = "off";

arriaii_lcell_comb \Equal6~0 (
	.dataa(!current_bank_0),
	.datab(!current_bank_1),
	.datac(!pipe_10_2),
	.datad(!pipe_11_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal6~0 .extended_lut = "off";
defparam \Equal6~0 .lut_mask = 64'h8421842184218421;
defparam \Equal6~0 .shared_arith = "off";

arriaii_lcell_comb \always12~1 (
	.dataa(!current_bank_2),
	.datab(!pipe_12_2),
	.datac(!pipefull_2),
	.datad(!\Equal6~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always12~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always12~1 .extended_lut = "off";
defparam \always12~1 .lut_mask = 64'h0F060F060F060F06;
defparam \always12~1 .shared_arith = "off";

arriaii_lcell_comb \always12~2 (
	.dataa(!pipe_12_2),
	.datab(!pipe_12_1),
	.datac(!\always12~0_combout ),
	.datad(!\Equal8~0_combout ),
	.datae(!\always12~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always12~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always12~2 .extended_lut = "off";
defparam \always12~2 .lut_mask = 64'h0000F6000000F600;
defparam \always12~2 .shared_arith = "off";

arriaii_lcell_comb \Equal18~0 (
	.dataa(!pipe_10_2),
	.datab(!pipe_10_3),
	.datac(!pipe_11_2),
	.datad(!pipe_11_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal18~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal18~0 .extended_lut = "off";
defparam \Equal18~0 .lut_mask = 64'h9009900990099009;
defparam \Equal18~0 .shared_arith = "off";

arriaii_lcell_comb \Equal16~0 (
	.dataa(!pipe_10_3),
	.datab(!pipe_10_1),
	.datac(!pipe_11_3),
	.datad(!pipe_11_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal16~0 .extended_lut = "off";
defparam \Equal16~0 .lut_mask = 64'h9009900990099009;
defparam \Equal16~0 .shared_arith = "off";

arriaii_lcell_comb \Equal14~0 (
	.dataa(!pipe_10_0),
	.datab(!pipe_11_0),
	.datac(!pipe_10_3),
	.datad(!pipe_11_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal14~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal14~0 .extended_lut = "off";
defparam \Equal14~0 .lut_mask = 64'h8421842184218421;
defparam \Equal14~0 .shared_arith = "off";

arriaii_lcell_comb \Equal12~0 (
	.dataa(!current_bank_2),
	.datab(!current_bank_0),
	.datac(!current_bank_1),
	.datad(!pipe_12_3),
	.datae(!pipe_10_3),
	.dataf(!pipe_11_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal12~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal12~0 .extended_lut = "off";
defparam \Equal12~0 .lut_mask = 64'h8040201008040201;
defparam \Equal12~0 .shared_arith = "off";

arriaii_lcell_comb \always13~0 (
	.dataa(!pipe_12_0),
	.datab(!pipe_12_3),
	.datac(!pipefull_3),
	.datad(!\Equal14~0_combout ),
	.datae(!\Equal12~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always13~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always13~0 .extended_lut = "off";
defparam \always13~0 .lut_mask = 64'h0F0600000F060000;
defparam \always13~0 .shared_arith = "off";

arriaii_lcell_comb \always13~1 (
	.dataa(!pipe_12_2),
	.datab(!pipe_12_3),
	.datac(!pipe_12_1),
	.datad(!\Equal18~0_combout ),
	.datae(!\Equal16~0_combout ),
	.dataf(!\always13~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always13~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always13~1 .extended_lut = "off";
defparam \always13~1 .lut_mask = 64'h00000000FF663C24;
defparam \always13~1 .shared_arith = "off";

dffeas \lookahead_allowed_to_cmd[3] (
	.clk(ctl_clk),
	.d(\always13~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(fetch1),
	.sload(gnd),
	.ena(vcc),
	.q(\lookahead_allowed_to_cmd[3]~q ),
	.prn(vcc));
defparam \lookahead_allowed_to_cmd[3] .is_wysiwyg = "true";
defparam \lookahead_allowed_to_cmd[3] .power_up = "low";

dffeas \lookahead_allowed_to_cmd[2] (
	.clk(ctl_clk),
	.d(\always12~2_combout ),
	.asdata(\lookahead_allowed_to_cmd[3]~q ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(fetch1),
	.ena(vcc),
	.q(\lookahead_allowed_to_cmd[2]~q ),
	.prn(vcc));
defparam \lookahead_allowed_to_cmd[2] .is_wysiwyg = "true";
defparam \lookahead_allowed_to_cmd[2] .power_up = "low";

dffeas \lookahead_allowed_to_cmd[1] (
	.clk(ctl_clk),
	.d(\always11~0_combout ),
	.asdata(\lookahead_allowed_to_cmd[2]~q ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(fetch1),
	.ena(vcc),
	.q(\lookahead_allowed_to_cmd[1]~q ),
	.prn(vcc));
defparam \lookahead_allowed_to_cmd[1] .is_wysiwyg = "true";
defparam \lookahead_allowed_to_cmd[1] .power_up = "low";

arriaii_lcell_comb \always39~0 (
	.dataa(!\just_did_activate~q ),
	.datab(!out_cmd_info_valid_2),
	.datac(!\lookahead_allowed_to_cmd[1]~q ),
	.datad(!out_cmd_can_activate_2),
	.datae(!out_cmd_bank_is_open_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always39~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always39~0 .extended_lut = "off";
defparam \always39~0 .lut_mask = 64'h0002000000020000;
defparam \always39~0 .shared_arith = "off";

arriaii_lcell_comb \always39~1 (
	.dataa(!\just_did_activate~q ),
	.datab(!out_cmd_info_valid_3),
	.datac(!\lookahead_allowed_to_cmd[2]~q ),
	.datad(!out_cmd_can_activate_3),
	.datae(!out_cmd_bank_is_open_3),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always39~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always39~1 .extended_lut = "off";
defparam \always39~1 .lut_mask = 64'h0002000000020000;
defparam \always39~1 .shared_arith = "off";

arriaii_lcell_comb \always14~1 (
	.dataa(!current_bank_0),
	.datab(!current_bank_1),
	.datac(!pipe_10_0),
	.datad(!pipe_11_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always14~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always14~1 .extended_lut = "off";
defparam \always14~1 .lut_mask = 64'h8421842184218421;
defparam \always14~1 .shared_arith = "off";

arriaii_lcell_comb \always10~0 (
	.dataa(!pipefull_0),
	.datab(!current_bank_2),
	.datac(!pipe_12_0),
	.datad(!\always14~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~0 .extended_lut = "off";
defparam \always10~0 .lut_mask = 64'h5514551455145514;
defparam \always10~0 .shared_arith = "off";

dffeas \lookahead_allowed_to_cmd[0] (
	.clk(ctl_clk),
	.d(\always10~0_combout ),
	.asdata(\lookahead_allowed_to_cmd[1]~q ),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(fetch1),
	.ena(vcc),
	.q(\lookahead_allowed_to_cmd[0]~q ),
	.prn(vcc));
defparam \lookahead_allowed_to_cmd[0] .is_wysiwyg = "true";
defparam \lookahead_allowed_to_cmd[0] .power_up = "low";

arriaii_lcell_comb \always39~2 (
	.dataa(!\just_did_activate~q ),
	.datab(!\lookahead_allowed_to_cmd[0]~q ),
	.datac(!out_cmd_info_valid_1),
	.datad(!out_cmd_can_activate_1),
	.datae(!out_cmd_bank_is_open_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always39~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always39~2 .extended_lut = "off";
defparam \always39~2 .lut_mask = 64'h0002000000020000;
defparam \always39~2 .shared_arith = "off";

arriaii_lcell_comb \to_bank_addr_r[2]~0 (
	.dataa(!\just_did_activate~q ),
	.datab(!\lookahead_allowed_to_cmd[3]~q ),
	.datac(!out_cmd_info_valid_4),
	.datad(!out_cmd_can_activate_4),
	.datae(!out_cmd_bank_is_open_4),
	.dataf(!\always39~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\to_bank_addr_r[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \to_bank_addr_r[2]~0 .extended_lut = "off";
defparam \to_bank_addr_r[2]~0 .lut_mask = 64'hFFFDFFFF00000000;
defparam \to_bank_addr_r[2]~0 .shared_arith = "off";

arriaii_lcell_comb \Selector20~1 (
	.dataa(!\state.DO2~q ),
	.datab(!\Selector20~0_combout ),
	.datac(!\always39~0_combout ),
	.datad(!\always39~1_combout ),
	.datae(!\to_bank_addr_r[2]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector20~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector20~1 .extended_lut = "off";
defparam \Selector20~1 .lut_mask = 64'h5555155555551555;
defparam \Selector20~1 .shared_arith = "off";

arriaii_lcell_comb \Selector20~2 (
	.dataa(!\state.DO2~q ),
	.datab(!\just_did_activate~q ),
	.datac(!\state.READWRITE~q ),
	.datad(!\Selector20~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector20~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector20~2 .extended_lut = "off";
defparam \Selector20~2 .lut_mask = 64'h20FF20FF20FF20FF;
defparam \Selector20~2 .shared_arith = "off";

dffeas just_did_activate(
	.clk(ctl_clk),
	.d(\Selector20~2_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\just_did_activate~q ),
	.prn(vcc));
defparam just_did_activate.is_wysiwyg = "true";
defparam just_did_activate.power_up = "low";

arriaii_lcell_comb \always38~12 (
	.dataa(!add_lat_on),
	.datab(!out_cmd_info_valid_0),
	.datac(!\just_did_activate~q ),
	.datad(!out_cmd_can_activate_0),
	.datae(!out_cmd_bank_is_open_0),
	.dataf(!can_al_activate_read),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always38~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always38~12 .extended_lut = "off";
defparam \always38~12 .lut_mask = 64'h0000000000100000;
defparam \always38~12 .shared_arith = "off";

arriaii_lcell_comb \always38~13 (
	.dataa(!out_cmd_info_valid_0),
	.datab(!out_cmd_bank_is_open_0),
	.datac(!always381),
	.datad(!always382),
	.datae(!\always38~12_combout ),
	.dataf(!out_cmd_can_read_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always38~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always38~13 .extended_lut = "off";
defparam \always38~13 .lut_mask = 64'hFFFF0000EEEF0000;
defparam \always38~13 .shared_arith = "off";

arriaii_lcell_comb \always38~14 (
	.dataa(!\current_read~q ),
	.datab(!do_write_r1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always38~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always38~14 .extended_lut = "off";
defparam \always38~14 .lut_mask = 64'h4444444444444444;
defparam \always38~14 .shared_arith = "off";

arriaii_lcell_comb \always38~15 (
	.dataa(!\always38~2_combout ),
	.datab(!\always38~5_combout ),
	.datac(!\always38~6_combout ),
	.datad(!\always38~11_combout ),
	.datae(!\always38~13_combout ),
	.dataf(!\always38~14_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always38~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always38~15 .extended_lut = "off";
defparam \always38~15 .lut_mask = 64'h57005700FFFF5700;
defparam \always38~15 .shared_arith = "off";

arriaii_lcell_comb \Selector6~0 (
	.dataa(!\state.DO2~q ),
	.datab(!\always38~15_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~0 .extended_lut = "off";
defparam \Selector6~0 .lut_mask = 64'h1111111111111111;
defparam \Selector6~0 .shared_arith = "off";

dffeas \state.READWRITE (
	.clk(ctl_clk),
	.d(\Selector6~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.READWRITE~q ),
	.prn(vcc));
defparam \state.READWRITE .is_wysiwyg = "true";
defparam \state.READWRITE .power_up = "low";

arriaii_lcell_comb \always15~1 (
	.dataa(!pipe_10_0),
	.datab(!pipefull_4),
	.datac(!pipe_10_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always15~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always15~1 .extended_lut = "off";
defparam \always15~1 .lut_mask = 64'h2121212121212121;
defparam \always15~1 .shared_arith = "off";

arriaii_lcell_comb \always15~2 (
	.dataa(!pipe_12_0),
	.datab(!pipe_11_0),
	.datac(!pipe_12_4),
	.datad(!pipe_11_4),
	.datae(!\always15~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always15~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always15~2 .extended_lut = "off";
defparam \always15~2 .lut_mask = 64'h0000842100008421;
defparam \always15~2 .shared_arith = "off";

arriaii_lcell_comb \Equal50~0 (
	.dataa(!pipe_25_0),
	.datab(!pipe_26_0),
	.datac(!pipe_25_6),
	.datad(!pipe_26_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal50~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal50~0 .extended_lut = "off";
defparam \Equal50~0 .lut_mask = 64'h8421842184218421;
defparam \Equal50~0 .shared_arith = "off";

arriaii_lcell_comb \Equal50~1 (
	.dataa(!pipe_22_0),
	.datab(!pipe_23_0),
	.datac(!pipe_22_6),
	.datad(!pipe_23_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal50~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal50~1 .extended_lut = "off";
defparam \Equal50~1 .lut_mask = 64'h8421842184218421;
defparam \Equal50~1 .shared_arith = "off";

arriaii_lcell_comb \Equal50~2 (
	.dataa(!pipe_21_0),
	.datab(!pipe_19_0),
	.datac(!pipe_20_0),
	.datad(!pipe_21_6),
	.datae(!pipe_19_6),
	.dataf(!pipe_20_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal50~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal50~2 .extended_lut = "off";
defparam \Equal50~2 .lut_mask = 64'h8040201008040201;
defparam \Equal50~2 .shared_arith = "off";

arriaii_lcell_comb \Equal50~3 (
	.dataa(!pipe_15_0),
	.datab(!pipe_13_0),
	.datac(!pipe_14_0),
	.datad(!pipe_15_6),
	.datae(!pipe_13_6),
	.dataf(!pipe_14_6),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal50~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal50~3 .extended_lut = "off";
defparam \Equal50~3 .lut_mask = 64'h8040201008040201;
defparam \Equal50~3 .shared_arith = "off";

arriaii_lcell_comb \Equal50~4 (
	.dataa(!pipe_16_0),
	.datab(!pipe_17_0),
	.datac(!pipe_16_6),
	.datad(!pipe_17_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal50~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal50~4 .extended_lut = "off";
defparam \Equal50~4 .lut_mask = 64'h8421842184218421;
defparam \Equal50~4 .shared_arith = "off";

arriaii_lcell_comb \Equal50~5 (
	.dataa(!pipe_18_0),
	.datab(!\Equal50~2_combout ),
	.datac(!\Equal50~3_combout ),
	.datad(!pipe_18_6),
	.datae(!\Equal50~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal50~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal50~5 .extended_lut = "off";
defparam \Equal50~5 .lut_mask = 64'h0000020100000201;
defparam \Equal50~5 .shared_arith = "off";

arriaii_lcell_comb \Equal50~6 (
	.dataa(!pipe_24_0),
	.datab(!\Equal50~0_combout ),
	.datac(!pipe_24_6),
	.datad(!\Equal50~1_combout ),
	.datae(!\Equal50~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal50~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal50~6 .extended_lut = "off";
defparam \Equal50~6 .lut_mask = 64'h0000002100000021;
defparam \Equal50~6 .shared_arith = "off";

arriaii_lcell_comb \always15~0 (
	.dataa(!pipe_12_0),
	.datab(!pipe_12_3),
	.datac(!pipefull_3),
	.datad(!\Equal14~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always15~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always15~0 .extended_lut = "off";
defparam \always15~0 .lut_mask = 64'h0009000900090009;
defparam \always15~0 .shared_arith = "off";

arriaii_lcell_comb \always15~5 (
	.dataa(!pipefull_6),
	.datab(!pipe_10_0),
	.datac(!pipe_10_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always15~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always15~5 .extended_lut = "off";
defparam \always15~5 .lut_mask = 64'h4141414141414141;
defparam \always15~5 .shared_arith = "off";

arriaii_lcell_comb \always15~6 (
	.dataa(!pipe_12_0),
	.datab(!pipe_11_0),
	.datac(!pipe_12_6),
	.datad(!pipe_11_6),
	.datae(!\always15~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always15~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always15~6 .extended_lut = "off";
defparam \always15~6 .lut_mask = 64'h0000842100008421;
defparam \always15~6 .shared_arith = "off";

arriaii_lcell_comb \always15~3 (
	.dataa(!pipefull_5),
	.datab(!pipe_10_0),
	.datac(!pipe_10_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always15~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always15~3 .extended_lut = "off";
defparam \always15~3 .lut_mask = 64'h4141414141414141;
defparam \always15~3 .shared_arith = "off";

arriaii_lcell_comb \always15~4 (
	.dataa(!pipe_12_0),
	.datab(!pipe_11_0),
	.datac(!pipe_12_5),
	.datad(!pipe_11_5),
	.datae(!\always15~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always15~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always15~4 .extended_lut = "off";
defparam \always15~4 .lut_mask = 64'h0000842100008421;
defparam \always15~4 .shared_arith = "off";

arriaii_lcell_comb \Equal41~1 (
	.dataa(!pipe_24_0),
	.datab(!pipe_22_0),
	.datac(!pipe_23_0),
	.datad(!pipe_24_3),
	.datae(!pipe_22_3),
	.dataf(!pipe_23_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal41~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal41~1 .extended_lut = "off";
defparam \Equal41~1 .lut_mask = 64'h8040201008040201;
defparam \Equal41~1 .shared_arith = "off";

arriaii_lcell_comb \Equal41~2 (
	.dataa(!pipe_21_0),
	.datab(!pipe_19_0),
	.datac(!pipe_20_0),
	.datad(!pipe_21_3),
	.datae(!pipe_19_3),
	.dataf(!pipe_20_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal41~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal41~2 .extended_lut = "off";
defparam \Equal41~2 .lut_mask = 64'h8040201008040201;
defparam \Equal41~2 .shared_arith = "off";

arriaii_lcell_comb \Equal41~3 (
	.dataa(!pipe_15_0),
	.datab(!pipe_13_0),
	.datac(!pipe_14_0),
	.datad(!pipe_15_3),
	.datae(!pipe_13_3),
	.dataf(!pipe_14_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal41~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal41~3 .extended_lut = "off";
defparam \Equal41~3 .lut_mask = 64'h8040201008040201;
defparam \Equal41~3 .shared_arith = "off";

arriaii_lcell_comb \Equal41~4 (
	.dataa(!pipe_18_0),
	.datab(!pipe_16_0),
	.datac(!pipe_17_0),
	.datad(!pipe_18_3),
	.datae(!pipe_16_3),
	.dataf(!pipe_17_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal41~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal41~4 .extended_lut = "off";
defparam \Equal41~4 .lut_mask = 64'h8040201008040201;
defparam \Equal41~4 .shared_arith = "off";

arriaii_lcell_comb \Equal41~5 (
	.dataa(!\Equal41~0_combout ),
	.datab(!\Equal41~1_combout ),
	.datac(!\Equal41~2_combout ),
	.datad(!\Equal41~3_combout ),
	.datae(!\Equal41~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal41~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal41~5 .extended_lut = "off";
defparam \Equal41~5 .lut_mask = 64'h0000000100000001;
defparam \Equal41~5 .shared_arith = "off";

arriaii_lcell_comb \Equal44~1 (
	.dataa(!pipe_24_0),
	.datab(!pipe_22_0),
	.datac(!pipe_23_0),
	.datad(!pipe_24_4),
	.datae(!pipe_22_4),
	.dataf(!pipe_23_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal44~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal44~1 .extended_lut = "off";
defparam \Equal44~1 .lut_mask = 64'h8040201008040201;
defparam \Equal44~1 .shared_arith = "off";

arriaii_lcell_comb \Equal44~2 (
	.dataa(!pipe_21_0),
	.datab(!pipe_19_0),
	.datac(!pipe_20_0),
	.datad(!pipe_21_4),
	.datae(!pipe_19_4),
	.dataf(!pipe_20_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal44~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal44~2 .extended_lut = "off";
defparam \Equal44~2 .lut_mask = 64'h8040201008040201;
defparam \Equal44~2 .shared_arith = "off";

arriaii_lcell_comb \Equal44~3 (
	.dataa(!pipe_15_0),
	.datab(!pipe_13_0),
	.datac(!pipe_14_0),
	.datad(!pipe_15_4),
	.datae(!pipe_13_4),
	.dataf(!pipe_14_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal44~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal44~3 .extended_lut = "off";
defparam \Equal44~3 .lut_mask = 64'h8040201008040201;
defparam \Equal44~3 .shared_arith = "off";

arriaii_lcell_comb \Equal44~4 (
	.dataa(!pipe_18_0),
	.datab(!pipe_16_0),
	.datac(!pipe_17_0),
	.datad(!pipe_18_4),
	.datae(!pipe_16_4),
	.dataf(!pipe_17_4),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal44~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal44~4 .extended_lut = "off";
defparam \Equal44~4 .lut_mask = 64'h8040201008040201;
defparam \Equal44~4 .shared_arith = "off";

arriaii_lcell_comb \Equal44~5 (
	.dataa(!\Equal44~0_combout ),
	.datab(!\Equal44~1_combout ),
	.datac(!\Equal44~2_combout ),
	.datad(!\Equal44~3_combout ),
	.datae(!\Equal44~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal44~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal44~5 .extended_lut = "off";
defparam \Equal44~5 .lut_mask = 64'h0000000100000001;
defparam \Equal44~5 .shared_arith = "off";

arriaii_lcell_comb \auto_autopch_req~0 (
	.dataa(!\Equal47~5_combout ),
	.datab(!\always15~0_combout ),
	.datac(!\always15~2_combout ),
	.datad(!\always15~4_combout ),
	.datae(!\Equal41~5_combout ),
	.dataf(!\Equal44~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_autopch_req~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_autopch_req~0 .extended_lut = "off";
defparam \auto_autopch_req~0 .lut_mask = 64'h3FBF0C8C33B30080;
defparam \auto_autopch_req~0 .shared_arith = "off";

arriaii_lcell_comb \auto_autopch_req_0~0 (
	.dataa(!pipe_25_0),
	.datab(!pipe_26_0),
	.datac(!pipe_24_0),
	.datad(!pipe_26_7),
	.datae(!pipe_24_7),
	.dataf(!pipe_25_7),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_autopch_req_0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_autopch_req_0~0 .extended_lut = "off";
defparam \auto_autopch_req_0~0 .lut_mask = 64'h8020080240100401;
defparam \auto_autopch_req_0~0 .shared_arith = "off";

arriaii_lcell_comb \auto_autopch_req_0~1 (
	.dataa(!pipe_22_0),
	.datab(!pipe_21_0),
	.datac(!pipe_21_7),
	.datad(!pipe_22_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_autopch_req_0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_autopch_req_0~1 .extended_lut = "off";
defparam \auto_autopch_req_0~1 .lut_mask = 64'h8241824182418241;
defparam \auto_autopch_req_0~1 .shared_arith = "off";

arriaii_lcell_comb \auto_autopch_req_0~3 (
	.dataa(!pipe_15_0),
	.datab(!pipe_16_0),
	.datac(!pipe_17_0),
	.datad(!pipe_17_7),
	.datae(!pipe_15_7),
	.dataf(!pipe_16_7),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_autopch_req_0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_autopch_req_0~3 .extended_lut = "off";
defparam \auto_autopch_req_0~3 .lut_mask = 64'h8008400420021001;
defparam \auto_autopch_req_0~3 .shared_arith = "off";

arriaii_lcell_comb \auto_autopch_req_0~4 (
	.dataa(!pipefull_7),
	.datab(!pipe_10_0),
	.datac(!pipe_11_0),
	.datad(!pipe_11_7),
	.datae(!pipe_10_7),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_autopch_req_0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_autopch_req_0~4 .extended_lut = "off";
defparam \auto_autopch_req_0~4 .lut_mask = 64'h4004100140041001;
defparam \auto_autopch_req_0~4 .shared_arith = "off";

arriaii_lcell_comb \auto_autopch_req_0~5 (
	.dataa(!pipe_12_0),
	.datab(!pipe_13_0),
	.datac(!pipe_14_0),
	.datad(!pipe_14_7),
	.datae(!pipe_12_7),
	.dataf(!pipe_13_7),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_autopch_req_0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_autopch_req_0~5 .extended_lut = "off";
defparam \auto_autopch_req_0~5 .lut_mask = 64'h8008400420021001;
defparam \auto_autopch_req_0~5 .shared_arith = "off";

arriaii_lcell_comb \auto_autopch_req_0~6 (
	.dataa(!\auto_autopch_req_0~2_combout ),
	.datab(!\auto_autopch_req_0~3_combout ),
	.datac(!\auto_autopch_req_0~4_combout ),
	.datad(!\auto_autopch_req_0~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_autopch_req_0~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_autopch_req_0~6 .extended_lut = "off";
defparam \auto_autopch_req_0~6 .lut_mask = 64'h0001000100010001;
defparam \auto_autopch_req_0~6 .shared_arith = "off";

arriaii_lcell_comb \auto_autopch_req_0~7 (
	.dataa(!pipe_23_0),
	.datab(!\auto_autopch_req_0~0_combout ),
	.datac(!pipe_23_7),
	.datad(!\auto_autopch_req_0~1_combout ),
	.datae(!\auto_autopch_req_0~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_autopch_req_0~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_autopch_req_0~7 .extended_lut = "off";
defparam \auto_autopch_req_0~7 .lut_mask = 64'hFFFFFFDEFFFFFFDE;
defparam \auto_autopch_req_0~7 .shared_arith = "off";

arriaii_lcell_comb \auto_autopch_req~4 (
	.dataa(!\always15~4_combout ),
	.datab(!\always15~2_combout ),
	.datac(!\Equal50~6_combout ),
	.datad(!\always15~0_combout ),
	.datae(!\always15~6_combout ),
	.dataf(!\auto_autopch_req~0_combout ),
	.datag(!\auto_autopch_req_0~7_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_autopch_req~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_autopch_req~4 .extended_lut = "on";
defparam \auto_autopch_req~4 .lut_mask = 64'h08008000FFFFFFFF;
defparam \auto_autopch_req~4 .shared_arith = "off";

arriaii_lcell_comb \auto_autopch_req~1 (
	.dataa(!fetch1),
	.datab(!pipefull_1),
	.datac(!pipefull_2),
	.datad(!\Equal4~0_combout ),
	.datae(!\Equal8~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_autopch_req~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_autopch_req~1 .extended_lut = "off";
defparam \auto_autopch_req~1 .lut_mask = 64'h5544504055445040;
defparam \auto_autopch_req~1 .shared_arith = "off";

arriaii_lcell_comb \always14~7 (
	.dataa(!current_bank_2),
	.datab(!pipe_12_2),
	.datac(!pipefull_2),
	.datad(!\Equal6~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always14~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always14~7 .extended_lut = "off";
defparam \always14~7 .lut_mask = 64'h0009000900090009;
defparam \always14~7 .shared_arith = "off";

arriaii_lcell_comb \always14~8 (
	.dataa(!pipefull_0),
	.datab(!current_bank_2),
	.datac(!pipe_12_0),
	.datad(!\always14~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always14~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always14~8 .extended_lut = "off";
defparam \always14~8 .lut_mask = 64'h0041004100410041;
defparam \always14~8 .shared_arith = "off";

arriaii_lcell_comb \always14~9 (
	.dataa(!current_bank_2),
	.datab(!pipefull_1),
	.datac(!pipe_12_1),
	.datad(!\always14~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always14~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always14~9 .extended_lut = "off";
defparam \always14~9 .lut_mask = 64'h0021002100210021;
defparam \always14~9 .shared_arith = "off";

arriaii_lcell_comb \auto_autopch_req_c~8 (
	.dataa(!\always14~6_combout ),
	.datab(!\always14~7_combout ),
	.datac(!\always14~8_combout ),
	.datad(!\always14~9_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_autopch_req_c~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_autopch_req_c~8 .extended_lut = "off";
defparam \auto_autopch_req_c~8 .lut_mask = 64'h8000800080008000;
defparam \auto_autopch_req_c~8 .shared_arith = "off";

arriaii_lcell_comb \always14~10 (
	.dataa(!current_bank_0),
	.datab(!pipefull_4),
	.datac(!pipe_10_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always14~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always14~10 .extended_lut = "off";
defparam \always14~10 .lut_mask = 64'h2121212121212121;
defparam \always14~10 .shared_arith = "off";

arriaii_lcell_comb \always14~11 (
	.dataa(!current_bank_2),
	.datab(!current_bank_1),
	.datac(!pipe_12_4),
	.datad(!pipe_11_4),
	.datae(!\always14~10_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always14~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always14~11 .extended_lut = "off";
defparam \always14~11 .lut_mask = 64'h0000842100008421;
defparam \always14~11 .shared_arith = "off";

dffeas \current_row[10] (
	.clk(ctl_clk),
	.d(pipe_23_0),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fetch1),
	.q(\current_row[10]~q ),
	.prn(vcc));
defparam \current_row[10] .is_wysiwyg = "true";
defparam \current_row[10] .power_up = "low";

dffeas \current_row[9] (
	.clk(ctl_clk),
	.d(pipe_22_0),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fetch1),
	.q(\current_row[9]~q ),
	.prn(vcc));
defparam \current_row[9] .is_wysiwyg = "true";
defparam \current_row[9] .power_up = "low";

arriaii_lcell_comb \Equal22~1 (
	.dataa(!\current_row[11]~q ),
	.datab(!\current_row[10]~q ),
	.datac(!\current_row[9]~q ),
	.datad(!pipe_24_2),
	.datae(!pipe_22_2),
	.dataf(!pipe_23_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal22~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal22~1 .extended_lut = "off";
defparam \Equal22~1 .lut_mask = 64'h8040080420100201;
defparam \Equal22~1 .shared_arith = "off";

dffeas \current_row[7] (
	.clk(ctl_clk),
	.d(pipe_20_0),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fetch1),
	.q(\current_row[7]~q ),
	.prn(vcc));
defparam \current_row[7] .is_wysiwyg = "true";
defparam \current_row[7] .power_up = "low";

dffeas \current_row[6] (
	.clk(ctl_clk),
	.d(pipe_19_0),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fetch1),
	.q(\current_row[6]~q ),
	.prn(vcc));
defparam \current_row[6] .is_wysiwyg = "true";
defparam \current_row[6] .power_up = "low";

arriaii_lcell_comb \Equal22~2 (
	.dataa(!\current_row[8]~q ),
	.datab(!\current_row[7]~q ),
	.datac(!\current_row[6]~q ),
	.datad(!pipe_21_2),
	.datae(!pipe_19_2),
	.dataf(!pipe_20_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal22~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal22~2 .extended_lut = "off";
defparam \Equal22~2 .lut_mask = 64'h8040080420100201;
defparam \Equal22~2 .shared_arith = "off";

dffeas \current_row[1] (
	.clk(ctl_clk),
	.d(pipe_14_0),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fetch1),
	.q(\current_row[1]~q ),
	.prn(vcc));
defparam \current_row[1] .is_wysiwyg = "true";
defparam \current_row[1] .power_up = "low";

dffeas \current_row[0] (
	.clk(ctl_clk),
	.d(pipe_13_0),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fetch1),
	.q(\current_row[0]~q ),
	.prn(vcc));
defparam \current_row[0] .is_wysiwyg = "true";
defparam \current_row[0] .power_up = "low";

arriaii_lcell_comb \Equal22~3 (
	.dataa(!\current_row[2]~q ),
	.datab(!\current_row[1]~q ),
	.datac(!\current_row[0]~q ),
	.datad(!pipe_15_2),
	.datae(!pipe_13_2),
	.dataf(!pipe_14_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal22~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal22~3 .extended_lut = "off";
defparam \Equal22~3 .lut_mask = 64'h8040080420100201;
defparam \Equal22~3 .shared_arith = "off";

dffeas \current_row[4] (
	.clk(ctl_clk),
	.d(pipe_17_0),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fetch1),
	.q(\current_row[4]~q ),
	.prn(vcc));
defparam \current_row[4] .is_wysiwyg = "true";
defparam \current_row[4] .power_up = "low";

dffeas \current_row[3] (
	.clk(ctl_clk),
	.d(pipe_16_0),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fetch1),
	.q(\current_row[3]~q ),
	.prn(vcc));
defparam \current_row[3] .is_wysiwyg = "true";
defparam \current_row[3] .power_up = "low";

arriaii_lcell_comb \Equal22~4 (
	.dataa(!\current_row[5]~q ),
	.datab(!\current_row[4]~q ),
	.datac(!\current_row[3]~q ),
	.datad(!pipe_18_2),
	.datae(!pipe_16_2),
	.dataf(!pipe_17_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal22~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal22~4 .extended_lut = "off";
defparam \Equal22~4 .lut_mask = 64'h8040080420100201;
defparam \Equal22~4 .shared_arith = "off";

arriaii_lcell_comb \Equal22~5 (
	.dataa(!\Equal22~0_combout ),
	.datab(!\Equal22~1_combout ),
	.datac(!\Equal22~2_combout ),
	.datad(!\Equal22~3_combout ),
	.datae(!\Equal22~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal22~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal22~5 .extended_lut = "off";
defparam \Equal22~5 .lut_mask = 64'h0000000100000001;
defparam \Equal22~5 .shared_arith = "off";

dffeas \current_row[11] (
	.clk(ctl_clk),
	.d(pipe_24_0),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fetch1),
	.q(\current_row[11]~q ),
	.prn(vcc));
defparam \current_row[11] .is_wysiwyg = "true";
defparam \current_row[11] .power_up = "low";

arriaii_lcell_comb \Equal20~1 (
	.dataa(!pipe_24_0),
	.datab(!pipe_22_0),
	.datac(!pipe_23_0),
	.datad(!\current_row[11]~q ),
	.datae(!\current_row[10]~q ),
	.dataf(!\current_row[9]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal20~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal20~1 .extended_lut = "off";
defparam \Equal20~1 .lut_mask = 64'h8040080420100201;
defparam \Equal20~1 .shared_arith = "off";

dffeas \current_row[8] (
	.clk(ctl_clk),
	.d(pipe_21_0),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fetch1),
	.q(\current_row[8]~q ),
	.prn(vcc));
defparam \current_row[8] .is_wysiwyg = "true";
defparam \current_row[8] .power_up = "low";

arriaii_lcell_comb \Equal20~2 (
	.dataa(!pipe_21_0),
	.datab(!pipe_19_0),
	.datac(!pipe_20_0),
	.datad(!\current_row[8]~q ),
	.datae(!\current_row[7]~q ),
	.dataf(!\current_row[6]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal20~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal20~2 .extended_lut = "off";
defparam \Equal20~2 .lut_mask = 64'h8040080420100201;
defparam \Equal20~2 .shared_arith = "off";

dffeas \current_row[2] (
	.clk(ctl_clk),
	.d(pipe_15_0),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fetch1),
	.q(\current_row[2]~q ),
	.prn(vcc));
defparam \current_row[2] .is_wysiwyg = "true";
defparam \current_row[2] .power_up = "low";

arriaii_lcell_comb \Equal20~3 (
	.dataa(!pipe_15_0),
	.datab(!pipe_13_0),
	.datac(!pipe_14_0),
	.datad(!\current_row[2]~q ),
	.datae(!\current_row[1]~q ),
	.dataf(!\current_row[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal20~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal20~3 .extended_lut = "off";
defparam \Equal20~3 .lut_mask = 64'h8040080420100201;
defparam \Equal20~3 .shared_arith = "off";

dffeas \current_row[5] (
	.clk(ctl_clk),
	.d(pipe_18_0),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fetch1),
	.q(\current_row[5]~q ),
	.prn(vcc));
defparam \current_row[5] .is_wysiwyg = "true";
defparam \current_row[5] .power_up = "low";

arriaii_lcell_comb \Equal20~4 (
	.dataa(!pipe_18_0),
	.datab(!pipe_16_0),
	.datac(!pipe_17_0),
	.datad(!\current_row[5]~q ),
	.datae(!\current_row[4]~q ),
	.dataf(!\current_row[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal20~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal20~4 .extended_lut = "off";
defparam \Equal20~4 .lut_mask = 64'h8040080420100201;
defparam \Equal20~4 .shared_arith = "off";

arriaii_lcell_comb \Equal20~5 (
	.dataa(!\Equal20~0_combout ),
	.datab(!\Equal20~1_combout ),
	.datac(!\Equal20~2_combout ),
	.datad(!\Equal20~3_combout ),
	.datae(!\Equal20~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal20~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal20~5 .extended_lut = "off";
defparam \Equal20~5 .lut_mask = 64'h0000000100000001;
defparam \Equal20~5 .shared_arith = "off";

arriaii_lcell_comb \Equal21~1 (
	.dataa(!\current_row[11]~q ),
	.datab(!\current_row[10]~q ),
	.datac(!\current_row[9]~q ),
	.datad(!pipe_24_1),
	.datae(!pipe_22_1),
	.dataf(!pipe_23_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal21~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal21~1 .extended_lut = "off";
defparam \Equal21~1 .lut_mask = 64'h8040080420100201;
defparam \Equal21~1 .shared_arith = "off";

arriaii_lcell_comb \Equal21~2 (
	.dataa(!\current_row[8]~q ),
	.datab(!\current_row[7]~q ),
	.datac(!\current_row[6]~q ),
	.datad(!pipe_21_1),
	.datae(!pipe_19_1),
	.dataf(!pipe_20_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal21~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal21~2 .extended_lut = "off";
defparam \Equal21~2 .lut_mask = 64'h8040080420100201;
defparam \Equal21~2 .shared_arith = "off";

arriaii_lcell_comb \Equal21~3 (
	.dataa(!\current_row[2]~q ),
	.datab(!\current_row[1]~q ),
	.datac(!\current_row[0]~q ),
	.datad(!pipe_15_1),
	.datae(!pipe_13_1),
	.dataf(!pipe_14_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal21~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal21~3 .extended_lut = "off";
defparam \Equal21~3 .lut_mask = 64'h8040080420100201;
defparam \Equal21~3 .shared_arith = "off";

arriaii_lcell_comb \Equal21~4 (
	.dataa(!\current_row[5]~q ),
	.datab(!\current_row[4]~q ),
	.datac(!\current_row[3]~q ),
	.datad(!pipe_18_1),
	.datae(!pipe_16_1),
	.dataf(!pipe_17_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal21~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal21~4 .extended_lut = "off";
defparam \Equal21~4 .lut_mask = 64'h8040080420100201;
defparam \Equal21~4 .shared_arith = "off";

arriaii_lcell_comb \Equal21~5 (
	.dataa(!\Equal21~0_combout ),
	.datab(!\Equal21~1_combout ),
	.datac(!\Equal21~2_combout ),
	.datad(!\Equal21~3_combout ),
	.datae(!\Equal21~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal21~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal21~5 .extended_lut = "off";
defparam \Equal21~5 .lut_mask = 64'h0000000100000001;
defparam \Equal21~5 .shared_arith = "off";

arriaii_lcell_comb \auto_autopch_req_c~9 (
	.dataa(!\always14~7_combout ),
	.datab(!\always14~8_combout ),
	.datac(!\always14~9_combout ),
	.datad(!\Equal22~5_combout ),
	.datae(!\Equal20~5_combout ),
	.dataf(!\Equal21~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_autopch_req_c~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_autopch_req_c~9 .extended_lut = "off";
defparam \auto_autopch_req_c~9 .lut_mask = 64'h7F3F4C0C73334000;
defparam \auto_autopch_req_c~9 .shared_arith = "off";

dffeas \current_row[13] (
	.clk(ctl_clk),
	.d(pipe_26_0),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fetch1),
	.q(\current_row[13]~q ),
	.prn(vcc));
defparam \current_row[13] .is_wysiwyg = "true";
defparam \current_row[13] .power_up = "low";

dffeas \current_row[12] (
	.clk(ctl_clk),
	.d(pipe_25_0),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fetch1),
	.q(\current_row[12]~q ),
	.prn(vcc));
defparam \current_row[12] .is_wysiwyg = "true";
defparam \current_row[12] .power_up = "low";

arriaii_lcell_comb \Equal23~0 (
	.dataa(!pipe_25_3),
	.datab(!pipe_26_3),
	.datac(!\current_row[13]~q ),
	.datad(!\current_row[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal23~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal23~0 .extended_lut = "off";
defparam \Equal23~0 .lut_mask = 64'h8241824182418241;
defparam \Equal23~0 .shared_arith = "off";

arriaii_lcell_comb \Equal23~2 (
	.dataa(!pipe_21_3),
	.datab(!pipe_19_3),
	.datac(!pipe_20_3),
	.datad(!\current_row[8]~q ),
	.datae(!\current_row[7]~q ),
	.dataf(!\current_row[6]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal23~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal23~2 .extended_lut = "off";
defparam \Equal23~2 .lut_mask = 64'h8040080420100201;
defparam \Equal23~2 .shared_arith = "off";

arriaii_lcell_comb \Equal23~3 (
	.dataa(!pipe_15_3),
	.datab(!pipe_13_3),
	.datac(!pipe_14_3),
	.datad(!\current_row[2]~q ),
	.datae(!\current_row[1]~q ),
	.dataf(!\current_row[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal23~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal23~3 .extended_lut = "off";
defparam \Equal23~3 .lut_mask = 64'h8040080420100201;
defparam \Equal23~3 .shared_arith = "off";

arriaii_lcell_comb \Equal23~4 (
	.dataa(!pipe_18_3),
	.datab(!pipe_16_3),
	.datac(!pipe_17_3),
	.datad(!\current_row[5]~q ),
	.datae(!\current_row[4]~q ),
	.dataf(!\current_row[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal23~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal23~4 .extended_lut = "off";
defparam \Equal23~4 .lut_mask = 64'h8040080420100201;
defparam \Equal23~4 .shared_arith = "off";

arriaii_lcell_comb \Equal23~5 (
	.dataa(!\Equal23~1_combout ),
	.datab(!\Equal23~2_combout ),
	.datac(!\Equal23~3_combout ),
	.datad(!\Equal23~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal23~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal23~5 .extended_lut = "off";
defparam \Equal23~5 .lut_mask = 64'h0001000100010001;
defparam \Equal23~5 .shared_arith = "off";

arriaii_lcell_comb \auto_autopch_req_c~10 (
	.dataa(!\always14~6_combout ),
	.datab(!\always14~7_combout ),
	.datac(!\always14~8_combout ),
	.datad(!\always14~9_combout ),
	.datae(!\Equal23~0_combout ),
	.dataf(!\Equal23~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_autopch_req_c~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_autopch_req_c~10 .extended_lut = "off";
defparam \auto_autopch_req_c~10 .lut_mask = 64'h4000400040000000;
defparam \auto_autopch_req_c~10 .shared_arith = "off";

arriaii_lcell_comb \Equal26~0 (
	.dataa(!pipe_25_4),
	.datab(!pipe_26_4),
	.datac(!\current_row[13]~q ),
	.datad(!\current_row[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal26~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal26~0 .extended_lut = "off";
defparam \Equal26~0 .lut_mask = 64'h8241824182418241;
defparam \Equal26~0 .shared_arith = "off";

arriaii_lcell_comb \Equal26~1 (
	.dataa(!pipe_22_4),
	.datab(!pipe_23_4),
	.datac(!\current_row[10]~q ),
	.datad(!\current_row[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal26~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal26~1 .extended_lut = "off";
defparam \Equal26~1 .lut_mask = 64'h8241824182418241;
defparam \Equal26~1 .shared_arith = "off";

arriaii_lcell_comb \Equal26~2 (
	.dataa(!pipe_21_4),
	.datab(!pipe_19_4),
	.datac(!pipe_20_4),
	.datad(!\current_row[8]~q ),
	.datae(!\current_row[7]~q ),
	.dataf(!\current_row[6]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal26~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal26~2 .extended_lut = "off";
defparam \Equal26~2 .lut_mask = 64'h8040080420100201;
defparam \Equal26~2 .shared_arith = "off";

arriaii_lcell_comb \Equal26~3 (
	.dataa(!pipe_15_4),
	.datab(!pipe_13_4),
	.datac(!pipe_14_4),
	.datad(!\current_row[2]~q ),
	.datae(!\current_row[1]~q ),
	.dataf(!\current_row[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal26~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal26~3 .extended_lut = "off";
defparam \Equal26~3 .lut_mask = 64'h8040080420100201;
defparam \Equal26~3 .shared_arith = "off";

arriaii_lcell_comb \Equal26~4 (
	.dataa(!pipe_16_4),
	.datab(!pipe_17_4),
	.datac(!\current_row[4]~q ),
	.datad(!\current_row[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal26~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal26~4 .extended_lut = "off";
defparam \Equal26~4 .lut_mask = 64'h8241824182418241;
defparam \Equal26~4 .shared_arith = "off";

arriaii_lcell_comb \Equal26~5 (
	.dataa(!pipe_18_4),
	.datab(!\current_row[5]~q ),
	.datac(!\Equal26~2_combout ),
	.datad(!\Equal26~3_combout ),
	.datae(!\Equal26~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal26~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal26~5 .extended_lut = "off";
defparam \Equal26~5 .lut_mask = 64'h0000000900000009;
defparam \Equal26~5 .shared_arith = "off";

arriaii_lcell_comb \Equal26~6 (
	.dataa(!pipe_24_4),
	.datab(!\current_row[11]~q ),
	.datac(!\Equal26~0_combout ),
	.datad(!\Equal26~1_combout ),
	.datae(!\Equal26~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal26~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal26~6 .extended_lut = "off";
defparam \Equal26~6 .lut_mask = 64'h0000000900000009;
defparam \Equal26~6 .shared_arith = "off";

arriaii_lcell_comb \auto_autopch_req_c~11 (
	.dataa(!\auto_autopch_req_c~7_combout ),
	.datab(!\auto_autopch_req_c~8_combout ),
	.datac(!\always14~11_combout ),
	.datad(!\auto_autopch_req_c~9_combout ),
	.datae(!\auto_autopch_req_c~10_combout ),
	.dataf(!\Equal26~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_autopch_req_c~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_autopch_req_c~11 .extended_lut = "off";
defparam \auto_autopch_req_c~11 .lut_mask = 64'hEC000000EF000000;
defparam \auto_autopch_req_c~11 .shared_arith = "off";

arriaii_lcell_comb \always15~7 (
	.dataa(!pipefull_1),
	.datab(!\Equal4~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always15~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always15~7 .extended_lut = "off";
defparam \always15~7 .lut_mask = 64'h1111111111111111;
defparam \always15~7 .shared_arith = "off";

arriaii_lcell_comb \Equal37~0 (
	.dataa(!pipe_25_0),
	.datab(!pipe_26_0),
	.datac(!pipe_25_1),
	.datad(!pipe_26_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal37~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal37~0 .extended_lut = "off";
defparam \Equal37~0 .lut_mask = 64'h8421842184218421;
defparam \Equal37~0 .shared_arith = "off";

arriaii_lcell_comb \Equal37~1 (
	.dataa(!pipe_22_0),
	.datab(!pipe_23_0),
	.datac(!pipe_22_1),
	.datad(!pipe_23_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal37~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal37~1 .extended_lut = "off";
defparam \Equal37~1 .lut_mask = 64'h8421842184218421;
defparam \Equal37~1 .shared_arith = "off";

arriaii_lcell_comb \Equal37~2 (
	.dataa(!pipe_21_0),
	.datab(!pipe_19_0),
	.datac(!pipe_20_0),
	.datad(!pipe_21_1),
	.datae(!pipe_19_1),
	.dataf(!pipe_20_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal37~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal37~2 .extended_lut = "off";
defparam \Equal37~2 .lut_mask = 64'h8040201008040201;
defparam \Equal37~2 .shared_arith = "off";

arriaii_lcell_comb \Equal37~3 (
	.dataa(!pipe_15_0),
	.datab(!pipe_13_0),
	.datac(!pipe_14_0),
	.datad(!pipe_15_1),
	.datae(!pipe_13_1),
	.dataf(!pipe_14_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal37~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal37~3 .extended_lut = "off";
defparam \Equal37~3 .lut_mask = 64'h8040201008040201;
defparam \Equal37~3 .shared_arith = "off";

arriaii_lcell_comb \Equal37~4 (
	.dataa(!pipe_16_0),
	.datab(!pipe_17_0),
	.datac(!pipe_16_1),
	.datad(!pipe_17_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal37~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal37~4 .extended_lut = "off";
defparam \Equal37~4 .lut_mask = 64'h8421842184218421;
defparam \Equal37~4 .shared_arith = "off";

arriaii_lcell_comb \Equal37~5 (
	.dataa(!pipe_18_0),
	.datab(!pipe_18_1),
	.datac(!\Equal37~2_combout ),
	.datad(!\Equal37~3_combout ),
	.datae(!\Equal37~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal37~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal37~5 .extended_lut = "off";
defparam \Equal37~5 .lut_mask = 64'h0000000900000009;
defparam \Equal37~5 .shared_arith = "off";

arriaii_lcell_comb \Equal37~6 (
	.dataa(!pipe_24_0),
	.datab(!pipe_24_1),
	.datac(!\Equal37~0_combout ),
	.datad(!\Equal37~1_combout ),
	.datae(!\Equal37~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal37~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal37~6 .extended_lut = "off";
defparam \Equal37~6 .lut_mask = 64'h0000000900000009;
defparam \Equal37~6 .shared_arith = "off";

arriaii_lcell_comb \Equal39~0 (
	.dataa(!pipe_25_0),
	.datab(!pipe_26_0),
	.datac(!pipe_25_2),
	.datad(!pipe_26_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal39~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal39~0 .extended_lut = "off";
defparam \Equal39~0 .lut_mask = 64'h8421842184218421;
defparam \Equal39~0 .shared_arith = "off";

arriaii_lcell_comb \Equal39~1 (
	.dataa(!pipe_22_0),
	.datab(!pipe_23_0),
	.datac(!pipe_22_2),
	.datad(!pipe_23_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal39~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal39~1 .extended_lut = "off";
defparam \Equal39~1 .lut_mask = 64'h8421842184218421;
defparam \Equal39~1 .shared_arith = "off";

arriaii_lcell_comb \Equal39~2 (
	.dataa(!pipe_21_0),
	.datab(!pipe_19_0),
	.datac(!pipe_20_0),
	.datad(!pipe_21_2),
	.datae(!pipe_19_2),
	.dataf(!pipe_20_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal39~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal39~2 .extended_lut = "off";
defparam \Equal39~2 .lut_mask = 64'h8040201008040201;
defparam \Equal39~2 .shared_arith = "off";

arriaii_lcell_comb \Equal39~3 (
	.dataa(!pipe_15_0),
	.datab(!pipe_13_0),
	.datac(!pipe_14_0),
	.datad(!pipe_15_2),
	.datae(!pipe_13_2),
	.dataf(!pipe_14_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal39~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal39~3 .extended_lut = "off";
defparam \Equal39~3 .lut_mask = 64'h8040201008040201;
defparam \Equal39~3 .shared_arith = "off";

arriaii_lcell_comb \Equal39~4 (
	.dataa(!pipe_16_0),
	.datab(!pipe_17_0),
	.datac(!pipe_16_2),
	.datad(!pipe_17_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal39~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal39~4 .extended_lut = "off";
defparam \Equal39~4 .lut_mask = 64'h8421842184218421;
defparam \Equal39~4 .shared_arith = "off";

arriaii_lcell_comb \Equal39~5 (
	.dataa(!pipe_18_0),
	.datab(!pipe_18_2),
	.datac(!\Equal39~2_combout ),
	.datad(!\Equal39~3_combout ),
	.datae(!\Equal39~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal39~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal39~5 .extended_lut = "off";
defparam \Equal39~5 .lut_mask = 64'h0000000900000009;
defparam \Equal39~5 .shared_arith = "off";

arriaii_lcell_comb \Equal39~6 (
	.dataa(!pipe_24_0),
	.datab(!pipe_24_2),
	.datac(!\Equal39~0_combout ),
	.datad(!\Equal39~1_combout ),
	.datae(!\Equal39~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal39~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal39~6 .extended_lut = "off";
defparam \Equal39~6 .lut_mask = 64'h0000000900000009;
defparam \Equal39~6 .shared_arith = "off";

arriaii_lcell_comb \auto_autopch_req~2 (
	.dataa(!fetch1),
	.datab(!pipefull_2),
	.datac(!\Equal8~0_combout ),
	.datad(!\always15~7_combout ),
	.datae(!\Equal37~6_combout ),
	.dataf(!\Equal39~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_autopch_req~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_autopch_req~2 .extended_lut = "off";
defparam \auto_autopch_req~2 .lut_mask = 64'h0155010000550000;
defparam \auto_autopch_req~2 .shared_arith = "off";

arriaii_lcell_comb \auto_autopch_req~3 (
	.dataa(!fetch1),
	.datab(!\auto_autopch_req~4_combout ),
	.datac(!\auto_autopch_req~1_combout ),
	.datad(!\auto_autopch_req_c~11_combout ),
	.datae(!\auto_autopch_req~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_autopch_req~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_autopch_req~3 .extended_lut = "off";
defparam \auto_autopch_req~3 .lut_mask = 64'hAB03FFFFAB03FFFF;
defparam \auto_autopch_req~3 .shared_arith = "off";

dffeas auto_autopch_req(
	.clk(ctl_clk),
	.d(\auto_autopch_req~3_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_autopch_req~q ),
	.prn(vcc));
defparam auto_autopch_req.is_wysiwyg = "true";
defparam auto_autopch_req.power_up = "low";

arriaii_lcell_comb \do_auto_precharge~0 (
	.dataa(!fetch1),
	.datab(!auto_refresh_logic_per_chip0int_refresh_req),
	.datac(!\auto_autopch_req~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\do_auto_precharge~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \do_auto_precharge~0 .extended_lut = "off";
defparam \do_auto_precharge~0 .lut_mask = 64'h2F2F2F2F2F2F2F2F;
defparam \do_auto_precharge~0 .shared_arith = "off";

arriaii_lcell_comb \current_read~_wirecell (
	.dataa(!\current_read~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\current_read~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \current_read~_wirecell .extended_lut = "off";
defparam \current_read~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \current_read~_wirecell .shared_arith = "off";

dffeas fetch_r(
	.clk(ctl_clk),
	.d(fetch1),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fetch_r~q ),
	.prn(vcc));
defparam fetch_r.is_wysiwyg = "true";
defparam fetch_r.power_up = "low";

arriaii_lcell_comb \current_burstcount_counter[1]~1 (
	.dataa(!\start_burst_r~q ),
	.datab(!\start_burst~q ),
	.datac(!\current_burstcount_counter_temp[1]~q ),
	.datad(!\current_burstcount_counter[0]~q ),
	.datae(!\fetch_r~q ),
	.dataf(!\current_burstcount_counter[1]~q ),
	.datag(!\burst_delay~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\current_burstcount_counter[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \current_burstcount_counter[1]~1 .extended_lut = "on";
defparam \current_burstcount_counter[1]~1 .lut_mask = 64'h00000F0F8FFF0F0F;
defparam \current_burstcount_counter[1]~1 .shared_arith = "off";

dffeas \current_burstcount_counter[1] (
	.clk(ctl_clk),
	.d(\current_burstcount_counter[1]~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\current_burstcount_counter[1]~q ),
	.prn(vcc));
defparam \current_burstcount_counter[1] .is_wysiwyg = "true";
defparam \current_burstcount_counter[1] .power_up = "low";

arriaii_lcell_comb \always39~3 (
	.dataa(!\current_burstcount_counter[1]~q ),
	.datab(!\current_burstcount_counter[0]~q ),
	.datac(!\burst_delay~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always39~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always39~3 .extended_lut = "off";
defparam \always39~3 .lut_mask = 64'h2F2F2F2F2F2F2F2F;
defparam \always39~3 .shared_arith = "off";

arriaii_lcell_comb \to_row_addr_r[5]~0 (
	.dataa(!\always39~0_combout ),
	.datab(!\always39~1_combout ),
	.datac(!\always39~2_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\to_row_addr_r[5]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \to_row_addr_r[5]~0 .extended_lut = "off";
defparam \to_row_addr_r[5]~0 .lut_mask = 64'h7070707070707070;
defparam \to_row_addr_r[5]~0 .shared_arith = "off";

arriaii_lcell_comb \to_row_addr_r[5]~1 (
	.dataa(!\always39~0_combout ),
	.datab(!\always39~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\to_row_addr_r[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \to_row_addr_r[5]~1 .extended_lut = "off";
defparam \to_row_addr_r[5]~1 .lut_mask = 64'h8888888888888888;
defparam \to_row_addr_r[5]~1 .shared_arith = "off";

arriaii_lcell_comb \Selector39~0 (
	.dataa(!pipe_13_0),
	.datab(!pipe_13_1),
	.datac(!pipe_13_3),
	.datad(!pipe_13_2),
	.datae(!\to_row_addr_r[5]~0_combout ),
	.dataf(!\to_row_addr_r[5]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector39~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector39~0 .extended_lut = "off";
defparam \Selector39~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Selector39~0 .shared_arith = "off";

arriaii_lcell_comb \to_bank_addr_r[2]~1 (
	.dataa(!\state.DO2~q ),
	.datab(!add_lat_on),
	.datac(!\always38~1_combout ),
	.datad(!can_al_activate_write),
	.datae(!can_al_activate_read),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\to_bank_addr_r[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \to_bank_addr_r[2]~1 .extended_lut = "off";
defparam \to_bank_addr_r[2]~1 .lut_mask = 64'hAEAFAFAFAEAFAFAF;
defparam \to_bank_addr_r[2]~1 .shared_arith = "off";

arriaii_lcell_comb \state.INIT~0 (
	.dataa(!ctl_init_success),
	.datab(!\state.INIT~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state.INIT~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state.INIT~0 .extended_lut = "off";
defparam \state.INIT~0 .lut_mask = 64'h7777777777777777;
defparam \state.INIT~0 .shared_arith = "off";

dffeas \state.INIT (
	.clk(ctl_clk),
	.d(\state.INIT~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.INIT~q ),
	.prn(vcc));
defparam \state.INIT .is_wysiwyg = "true";
defparam \state.INIT .power_up = "low";

arriaii_lcell_comb \to_bank_addr_r[2]~2 (
	.dataa(!\state.DO2~q ),
	.datab(!\state.READWRITE~q ),
	.datac(!\state.INIT~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\to_bank_addr_r[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \to_bank_addr_r[2]~2 .extended_lut = "off";
defparam \to_bank_addr_r[2]~2 .lut_mask = 64'h0707070707070707;
defparam \to_bank_addr_r[2]~2 .shared_arith = "off";

arriaii_lcell_comb \to_row_addr_r[5]~2 (
	.dataa(!\always39~0_combout ),
	.datab(!\always39~1_combout ),
	.datac(!\to_bank_addr_r[2]~0_combout ),
	.datad(!\to_bank_addr_r[2]~1_combout ),
	.datae(!\to_bank_addr_r[2]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\to_row_addr_r[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \to_row_addr_r[5]~2 .extended_lut = "off";
defparam \to_row_addr_r[5]~2 .lut_mask = 64'h08FF080008FF0800;
defparam \to_row_addr_r[5]~2 .shared_arith = "off";

arriaii_lcell_comb \Selector38~0 (
	.dataa(!pipe_14_0),
	.datab(!pipe_14_1),
	.datac(!pipe_14_3),
	.datad(!pipe_14_2),
	.datae(!\to_row_addr_r[5]~0_combout ),
	.dataf(!\to_row_addr_r[5]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector38~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector38~0 .extended_lut = "off";
defparam \Selector38~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Selector38~0 .shared_arith = "off";

arriaii_lcell_comb \to_addr~0 (
	.dataa(!\current_burstcount_counter[1]~q ),
	.datab(!\current_burstcount_counter[0]~q ),
	.datac(!\burst_delay~q ),
	.datad(!\current_col[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\to_addr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \to_addr~0 .extended_lut = "off";
defparam \to_addr~0 .lut_mask = 64'h002F002F002F002F;
defparam \to_addr~0 .shared_arith = "off";

arriaii_lcell_comb \Selector37~0 (
	.dataa(!pipe_15_0),
	.datab(!pipe_15_1),
	.datac(!pipe_15_3),
	.datad(!pipe_15_2),
	.datae(!\to_row_addr_r[5]~0_combout ),
	.dataf(!\to_row_addr_r[5]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector37~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector37~0 .extended_lut = "off";
defparam \Selector37~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Selector37~0 .shared_arith = "off";

dffeas \current_col[3] (
	.clk(ctl_clk),
	.d(pipe_3_0),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fetch1),
	.q(\current_col[3]~q ),
	.prn(vcc));
defparam \current_col[3] .is_wysiwyg = "true";
defparam \current_col[3] .power_up = "low";

arriaii_lcell_comb \Selector36~0 (
	.dataa(!pipe_16_0),
	.datab(!pipe_16_1),
	.datac(!pipe_16_3),
	.datad(!pipe_16_2),
	.datae(!\to_row_addr_r[5]~0_combout ),
	.dataf(!\to_row_addr_r[5]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector36~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector36~0 .extended_lut = "off";
defparam \Selector36~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Selector36~0 .shared_arith = "off";

dffeas \current_col[4] (
	.clk(ctl_clk),
	.d(pipe_4_0),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fetch1),
	.q(\current_col[4]~q ),
	.prn(vcc));
defparam \current_col[4] .is_wysiwyg = "true";
defparam \current_col[4] .power_up = "low";

arriaii_lcell_comb \Selector35~0 (
	.dataa(!pipe_17_0),
	.datab(!pipe_17_1),
	.datac(!pipe_17_3),
	.datad(!pipe_17_2),
	.datae(!\to_row_addr_r[5]~0_combout ),
	.dataf(!\to_row_addr_r[5]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector35~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector35~0 .extended_lut = "off";
defparam \Selector35~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Selector35~0 .shared_arith = "off";

dffeas \current_col[5] (
	.clk(ctl_clk),
	.d(pipe_5_0),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fetch1),
	.q(\current_col[5]~q ),
	.prn(vcc));
defparam \current_col[5] .is_wysiwyg = "true";
defparam \current_col[5] .power_up = "low";

arriaii_lcell_comb \Selector34~0 (
	.dataa(!pipe_18_0),
	.datab(!pipe_18_1),
	.datac(!pipe_18_3),
	.datad(!pipe_18_2),
	.datae(!\to_row_addr_r[5]~0_combout ),
	.dataf(!\to_row_addr_r[5]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector34~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector34~0 .extended_lut = "off";
defparam \Selector34~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Selector34~0 .shared_arith = "off";

dffeas \current_col[6] (
	.clk(ctl_clk),
	.d(pipe_6_0),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fetch1),
	.q(\current_col[6]~q ),
	.prn(vcc));
defparam \current_col[6] .is_wysiwyg = "true";
defparam \current_col[6] .power_up = "low";

arriaii_lcell_comb \Selector33~0 (
	.dataa(!pipe_19_0),
	.datab(!pipe_19_1),
	.datac(!pipe_19_3),
	.datad(!pipe_19_2),
	.datae(!\to_row_addr_r[5]~0_combout ),
	.dataf(!\to_row_addr_r[5]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector33~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector33~0 .extended_lut = "off";
defparam \Selector33~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Selector33~0 .shared_arith = "off";

dffeas \current_col[7] (
	.clk(ctl_clk),
	.d(pipe_7_0),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fetch1),
	.q(\current_col[7]~q ),
	.prn(vcc));
defparam \current_col[7] .is_wysiwyg = "true";
defparam \current_col[7] .power_up = "low";

arriaii_lcell_comb \Selector32~0 (
	.dataa(!pipe_20_0),
	.datab(!pipe_20_1),
	.datac(!pipe_20_3),
	.datad(!pipe_20_2),
	.datae(!\to_row_addr_r[5]~0_combout ),
	.dataf(!\to_row_addr_r[5]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector32~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector32~0 .extended_lut = "off";
defparam \Selector32~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Selector32~0 .shared_arith = "off";

dffeas \current_col[8] (
	.clk(ctl_clk),
	.d(pipe_8_0),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fetch1),
	.q(\current_col[8]~q ),
	.prn(vcc));
defparam \current_col[8] .is_wysiwyg = "true";
defparam \current_col[8] .power_up = "low";

arriaii_lcell_comb \Selector31~0 (
	.dataa(!pipe_21_0),
	.datab(!pipe_21_1),
	.datac(!pipe_21_3),
	.datad(!pipe_21_2),
	.datae(!\to_row_addr_r[5]~0_combout ),
	.dataf(!\to_row_addr_r[5]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector31~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector31~0 .extended_lut = "off";
defparam \Selector31~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Selector31~0 .shared_arith = "off";

dffeas \current_col[9] (
	.clk(ctl_clk),
	.d(pipe_9_0),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fetch1),
	.q(\current_col[9]~q ),
	.prn(vcc));
defparam \current_col[9] .is_wysiwyg = "true";
defparam \current_col[9] .power_up = "low";

arriaii_lcell_comb \Selector30~0 (
	.dataa(!pipe_22_0),
	.datab(!pipe_22_1),
	.datac(!pipe_22_3),
	.datad(!pipe_22_2),
	.datae(!\to_row_addr_r[5]~0_combout ),
	.dataf(!\to_row_addr_r[5]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector30~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector30~0 .extended_lut = "off";
defparam \Selector30~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Selector30~0 .shared_arith = "off";

arriaii_lcell_comb \Selector29~0 (
	.dataa(!pipe_23_0),
	.datab(!pipe_23_1),
	.datac(!pipe_23_3),
	.datad(!pipe_23_2),
	.datae(!\to_row_addr_r[5]~0_combout ),
	.dataf(!\to_row_addr_r[5]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector29~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector29~0 .extended_lut = "off";
defparam \Selector29~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Selector29~0 .shared_arith = "off";

arriaii_lcell_comb \Selector28~0 (
	.dataa(!pipe_24_0),
	.datab(!pipe_24_1),
	.datac(!pipe_24_3),
	.datad(!pipe_24_2),
	.datae(!\to_row_addr_r[5]~0_combout ),
	.dataf(!\to_row_addr_r[5]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector28~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector28~0 .extended_lut = "off";
defparam \Selector28~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Selector28~0 .shared_arith = "off";

arriaii_lcell_comb \Selector27~0 (
	.dataa(!pipe_25_0),
	.datab(!pipe_25_1),
	.datac(!pipe_25_3),
	.datad(!pipe_25_2),
	.datae(!\to_row_addr_r[5]~0_combout ),
	.dataf(!\to_row_addr_r[5]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector27~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector27~0 .extended_lut = "off";
defparam \Selector27~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Selector27~0 .shared_arith = "off";

arriaii_lcell_comb \Selector26~0 (
	.dataa(!pipe_26_0),
	.datab(!pipe_26_1),
	.datac(!pipe_26_3),
	.datad(!pipe_26_2),
	.datae(!\to_row_addr_r[5]~0_combout ),
	.dataf(!\to_row_addr_r[5]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector26~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector26~0 .extended_lut = "off";
defparam \Selector26~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Selector26~0 .shared_arith = "off";

arriaii_lcell_comb \Selector2~0 (
	.dataa(!\state.FETCH~q ),
	.datab(!do_refresh_r1),
	.datac(!auto_refresh_logic_per_chip0int_refresh_req),
	.datad(!\state.READWRITE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'hAE00AE00AE00AE00;
defparam \Selector2~0 .shared_arith = "off";

arriaii_lcell_comb \Selector15~0 (
	.dataa(!\state.REFRESH~q ),
	.datab(!\state.FETCH~q ),
	.datac(!\for_chip_refresh_req~q ),
	.datad(!\state.PCHALL~q ),
	.datae(!\Selector7~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector15~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector15~0 .extended_lut = "off";
defparam \Selector15~0 .lut_mask = 64'h0B0FFFFF0B0FFFFF;
defparam \Selector15~0 .shared_arith = "off";

dffeas for_chip_refresh_req(
	.clk(ctl_clk),
	.d(\Selector15~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\for_chip_refresh_req~q ),
	.prn(vcc));
defparam for_chip_refresh_req.is_wysiwyg = "true";
defparam for_chip_refresh_req.power_up = "low";

arriaii_lcell_comb \Selector2~1 (
	.dataa(!\for_chip[0]~q ),
	.datab(!\state.REFRESH~q ),
	.datac(!\for_chip_refresh_req~q ),
	.datad(!\state.PCHALL~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~1 .extended_lut = "off";
defparam \Selector2~1 .lut_mask = 64'h22F222F222F222F2;
defparam \Selector2~1 .shared_arith = "off";

arriaii_lcell_comb \Selector2~2 (
	.dataa(!ctl_init_success),
	.datab(!fetch1),
	.datac(!\state.INIT~q ),
	.datad(!\Selector2~0_combout ),
	.datae(!\Selector2~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~2 .extended_lut = "off";
defparam \Selector2~2 .lut_mask = 64'hDC50FFFFDC50FFFF;
defparam \Selector2~2 .shared_arith = "off";

dffeas \state.FETCH (
	.clk(ctl_clk),
	.d(\Selector2~2_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.FETCH~q ),
	.prn(vcc));
defparam \state.FETCH .is_wysiwyg = "true";
defparam \state.FETCH .power_up = "low";

arriaii_lcell_comb \Selector7~0 (
	.dataa(!fetch1),
	.datab(!\state.FETCH~q ),
	.datac(!do_refresh_r1),
	.datad(!auto_refresh_logic_per_chip0int_refresh_req),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector7~0 .extended_lut = "off";
defparam \Selector7~0 .lut_mask = 64'h0020002000200020;
defparam \Selector7~0 .shared_arith = "off";

arriaii_lcell_comb \Selector4~1 (
	.dataa(!\for_chip[0]~q ),
	.datab(!auto_refresh_logic_per_chip0int_refresh_req),
	.datac(!\Selector4~0_combout ),
	.datad(!\Selector7~0_combout ),
	.datae(!out_cs_all_banks_closed_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector4~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~1 .extended_lut = "off";
defparam \Selector4~1 .lut_mask = 64'h0537050505370505;
defparam \Selector4~1 .shared_arith = "off";

dffeas \state.PCHALL (
	.clk(ctl_clk),
	.d(\Selector4~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.PCHALL~q ),
	.prn(vcc));
defparam \state.PCHALL .is_wysiwyg = "true";
defparam \state.PCHALL .power_up = "low";

arriaii_lcell_comb \Selector4~0 (
	.dataa(!\for_chip_refresh_req~q ),
	.datab(!\state.PCHALL~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~0 .extended_lut = "off";
defparam \Selector4~0 .lut_mask = 64'h1111111111111111;
defparam \Selector4~0 .shared_arith = "off";

arriaii_lcell_comb \Selector7~1 (
	.dataa(!\for_chip[0]~q ),
	.datab(!\state.REFRESH~q ),
	.datac(!\Selector4~0_combout ),
	.datad(!\Selector7~0_combout ),
	.datae(!out_cs_all_banks_closed_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector7~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector7~1 .extended_lut = "off";
defparam \Selector7~1 .lut_mask = 64'h1B1B1BFF1B1B1BFF;
defparam \Selector7~1 .shared_arith = "off";

dffeas \state.REFRESH (
	.clk(ctl_clk),
	.d(\Selector7~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.REFRESH~q ),
	.prn(vcc));
defparam \state.REFRESH .is_wysiwyg = "true";
defparam \state.REFRESH .power_up = "low";

arriaii_lcell_comb \Selector0~0 (
	.dataa(!\state.DO2~q ),
	.datab(!\always38~15_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h4444444444444444;
defparam \Selector0~0 .shared_arith = "off";

arriaii_lcell_comb \Selector0~1 (
	.dataa(!fetch1),
	.datab(!\state.FETCH~q ),
	.datac(!\Selector0~0_combout ),
	.datad(!\state.READWRITE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~1 .extended_lut = "off";
defparam \Selector0~1 .lut_mask = 64'h1F5F1F5F1F5F1F5F;
defparam \Selector0~1 .shared_arith = "off";

dffeas \state.DO2 (
	.clk(ctl_clk),
	.d(\Selector0~1_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.DO2~q ),
	.prn(vcc));
defparam \state.DO2 .is_wysiwyg = "true";
defparam \state.DO2 .power_up = "low";

arriaii_lcell_comb \Selector11~1 (
	.dataa(!\state.FETCH~q ),
	.datab(!\state.DO2~q ),
	.datac(!\state.READWRITE~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector11~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector11~1 .extended_lut = "off";
defparam \Selector11~1 .lut_mask = 64'h8080808080808080;
defparam \Selector11~1 .shared_arith = "off";

arriaii_lcell_comb \Selector14~0 (
	.dataa(!do_precharge_all_r1),
	.datab(!out_cs_can_refresh_0),
	.datac(!\for_chip[0]~q ),
	.datad(!\state.REFRESH~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector14~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector14~0 .extended_lut = "off";
defparam \Selector14~0 .lut_mask = 64'h005D005D005D005D;
defparam \Selector14~0 .shared_arith = "off";

arriaii_lcell_comb \Selector14~1 (
	.dataa(!out_cs_can_precharge_all_0),
	.datab(!\for_chip_refresh_req~q ),
	.datac(!\state.PCHALL~q ),
	.datad(!\Selector14~0_combout ),
	.datae(!\state.INIT~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector14~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector14~1 .extended_lut = "off";
defparam \Selector14~1 .lut_mask = 64'h0000F1000000F100;
defparam \Selector14~1 .shared_arith = "off";

arriaii_lcell_comb \for_chip_saved[0]~0 (
	.dataa(!fetch1),
	.datab(!\state.FETCH~q ),
	.datac(!do_refresh_r1),
	.datad(!auto_refresh_logic_per_chip0int_refresh_req),
	.datae(!\for_chip_saved[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\for_chip_saved[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \for_chip_saved[0]~0 .extended_lut = "off";
defparam \for_chip_saved[0]~0 .lut_mask = 64'h0020FFFF0020FFFF;
defparam \for_chip_saved[0]~0 .shared_arith = "off";

dffeas \for_chip_saved[0] (
	.clk(ctl_clk),
	.d(\for_chip_saved[0]~0_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\for_chip_saved[0]~q ),
	.prn(vcc));
defparam \for_chip_saved[0] .is_wysiwyg = "true";
defparam \for_chip_saved[0] .power_up = "low";

arriaii_lcell_comb \Selector14~2 (
	.dataa(!\for_chip[0]~q ),
	.datab(!\state.REFRESH~q ),
	.datac(!\for_chip_refresh_req~q ),
	.datad(!\state.PCHALL~q ),
	.datae(!\for_chip_saved[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector14~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector14~2 .extended_lut = "off";
defparam \Selector14~2 .lut_mask = 64'h0000222A0000222A;
defparam \Selector14~2 .shared_arith = "off";

arriaii_lcell_comb \Selector14~3 (
	.dataa(!\for_chip[0]~q ),
	.datab(!\Selector11~1_combout ),
	.datac(!\Selector7~0_combout ),
	.datad(!\Selector14~1_combout ),
	.datae(!\Selector14~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector14~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector14~3 .extended_lut = "off";
defparam \Selector14~3 .lut_mask = 64'h5F4FFFFF5F4FFFFF;
defparam \Selector14~3 .shared_arith = "off";

dffeas \for_chip[0] (
	.clk(ctl_clk),
	.d(\Selector14~3_combout ),
	.asdata(vcc),
	.clrn(ctl_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\for_chip[0]~q ),
	.prn(vcc));
defparam \for_chip[0] .is_wysiwyg = "true";
defparam \for_chip[0] .power_up = "low";

arriaii_lcell_comb \Selector10~0 (
	.dataa(!do_precharge_all_r1),
	.datab(!out_cs_can_refresh_0),
	.datac(!\for_chip[0]~q ),
	.datad(!\state.REFRESH~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector10~0 .extended_lut = "off";
defparam \Selector10~0 .lut_mask = 64'h0002000200020002;
defparam \Selector10~0 .shared_arith = "off";

arriaii_lcell_comb \Selector10~1 (
	.dataa(!int_refresh_ack1),
	.datab(!\state.REFRESH~q ),
	.datac(!\Selector10~0_combout ),
	.datad(!\state.FETCH~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector10~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector10~1 .extended_lut = "off";
defparam \Selector10~1 .lut_mask = 64'h4F0F4F0F4F0F4F0F;
defparam \Selector10~1 .shared_arith = "off";

arriaii_lcell_comb \Selector11~0 (
	.dataa(!fetch1),
	.datab(!\state.FETCH~q ),
	.datac(!do_refresh_r1),
	.datad(!auto_refresh_logic_per_chip0int_refresh_req),
	.datae(!\state.DO2~q ),
	.dataf(!\always38~15_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector11~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector11~0 .extended_lut = "off";
defparam \Selector11~0 .lut_mask = 64'h220222022202FF02;
defparam \Selector11~0 .shared_arith = "off";

arriaii_lcell_comb \Selector11~2 (
	.dataa(!fetch1),
	.datab(!always38),
	.datac(!pipefull_0),
	.datad(!\Selector11~0_combout ),
	.datae(!\Selector0~0_combout ),
	.dataf(!\Selector11~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector11~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector11~2 .extended_lut = "off";
defparam \Selector11~2 .lut_mask = 64'h00CF55DF55DF55DF;
defparam \Selector11~2 .shared_arith = "off";

arriaii_lcell_comb \do_precharge_all~0 (
	.dataa(!\for_chip[0]~q ),
	.datab(!out_cs_can_precharge_all_0),
	.datac(!\for_chip_refresh_req~q ),
	.datad(!\state.PCHALL~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\do_precharge_all~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \do_precharge_all~0 .extended_lut = "off";
defparam \do_precharge_all~0 .lut_mask = 64'h0001000100010001;
defparam \do_precharge_all~0 .shared_arith = "off";

arriaii_lcell_comb \Selector22~0 (
	.dataa(!\state.READWRITE~q ),
	.datab(!\do_precharge_all~0_combout ),
	.datac(!\Selector20~1_combout ),
	.datad(!\Selector10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector22~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector22~0 .extended_lut = "off";
defparam \Selector22~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \Selector22~0 .shared_arith = "off";

arriaii_lcell_comb \Selector23~0 (
	.dataa(!\always39~0_combout ),
	.datab(!\always39~1_combout ),
	.datac(!\to_bank_addr_r[2]~0_combout ),
	.datad(!pipe_12_2),
	.datae(!pipe_12_3),
	.dataf(!pipe_12_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector23~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector23~0 .extended_lut = "off";
defparam \Selector23~0 .lut_mask = 64'h002280A25577D5F7;
defparam \Selector23~0 .shared_arith = "off";

arriaii_lcell_comb \Selector23~1 (
	.dataa(!current_bank_2),
	.datab(!\always39~2_combout ),
	.datac(!pipe_12_0),
	.datad(!\Selector23~0_combout ),
	.datae(!\to_bank_addr_r[2]~1_combout ),
	.dataf(!\to_bank_addr_r[2]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector23~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector23~1 .extended_lut = "off";
defparam \Selector23~1 .lut_mask = 64'h03CF000003CF5555;
defparam \Selector23~1 .shared_arith = "off";

arriaii_lcell_comb \Selector25~0 (
	.dataa(!\always39~0_combout ),
	.datab(!\always39~1_combout ),
	.datac(!\to_bank_addr_r[2]~0_combout ),
	.datad(!pipe_10_2),
	.datae(!pipe_10_3),
	.dataf(!pipe_10_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector25~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector25~0 .extended_lut = "off";
defparam \Selector25~0 .lut_mask = 64'h002280A25577D5F7;
defparam \Selector25~0 .shared_arith = "off";

arriaii_lcell_comb \Selector25~1 (
	.dataa(!current_bank_0),
	.datab(!\always39~2_combout ),
	.datac(!pipe_10_0),
	.datad(!\to_bank_addr_r[2]~1_combout ),
	.datae(!\to_bank_addr_r[2]~2_combout ),
	.dataf(!\Selector25~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector25~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector25~1 .extended_lut = "off";
defparam \Selector25~1 .lut_mask = 64'h03000355CF00CF55;
defparam \Selector25~1 .shared_arith = "off";

arriaii_lcell_comb \Selector24~0 (
	.dataa(!\always39~0_combout ),
	.datab(!\always39~1_combout ),
	.datac(!\to_bank_addr_r[2]~0_combout ),
	.datad(!pipe_11_2),
	.datae(!pipe_11_3),
	.dataf(!pipe_11_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector24~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector24~0 .extended_lut = "off";
defparam \Selector24~0 .lut_mask = 64'h002280A25577D5F7;
defparam \Selector24~0 .shared_arith = "off";

arriaii_lcell_comb \Selector24~1 (
	.dataa(!current_bank_1),
	.datab(!\always39~2_combout ),
	.datac(!pipe_11_0),
	.datad(!\to_bank_addr_r[2]~1_combout ),
	.datae(!\to_bank_addr_r[2]~2_combout ),
	.dataf(!\Selector24~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector24~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector24~1 .extended_lut = "off";
defparam \Selector24~1 .lut_mask = 64'h03000355CF00CF55;
defparam \Selector24~1 .shared_arith = "off";

arriaii_lcell_comb \new_gen_rdwr_data_valid~0 (
	.dataa(!\state.READWRITE~q ),
	.datab(!\always29~0_combout ),
	.datac(!\always39~3_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\new_gen_rdwr_data_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \new_gen_rdwr_data_valid~0 .extended_lut = "off";
defparam \new_gen_rdwr_data_valid~0 .lut_mask = 64'h3737373737373737;
defparam \new_gen_rdwr_data_valid~0 .shared_arith = "off";

endmodule

module ddr3_int_ddr3_int_phy (
	q_b_0,
	q_b_64,
	q_b_1,
	q_b_65,
	q_b_2,
	q_b_66,
	q_b_3,
	q_b_67,
	q_b_4,
	q_b_68,
	q_b_5,
	q_b_69,
	q_b_6,
	q_b_70,
	q_b_7,
	q_b_71,
	q_b_16,
	q_b_80,
	q_b_17,
	q_b_81,
	q_b_18,
	q_b_82,
	q_b_19,
	q_b_83,
	q_b_20,
	q_b_84,
	q_b_21,
	q_b_85,
	q_b_22,
	q_b_86,
	q_b_23,
	q_b_87,
	q_b_32,
	q_b_96,
	q_b_33,
	q_b_97,
	q_b_34,
	q_b_98,
	q_b_35,
	q_b_99,
	q_b_36,
	q_b_100,
	q_b_37,
	q_b_101,
	q_b_38,
	q_b_102,
	q_b_39,
	q_b_103,
	q_b_48,
	q_b_112,
	q_b_49,
	q_b_113,
	q_b_50,
	q_b_114,
	q_b_51,
	q_b_115,
	q_b_52,
	q_b_116,
	q_b_53,
	q_b_117,
	q_b_54,
	q_b_118,
	q_b_55,
	q_b_119,
	q_b_8,
	q_b_72,
	q_b_9,
	q_b_73,
	q_b_10,
	q_b_74,
	q_b_11,
	q_b_75,
	q_b_12,
	q_b_76,
	q_b_13,
	q_b_77,
	q_b_14,
	q_b_78,
	q_b_15,
	q_b_79,
	q_b_24,
	q_b_88,
	q_b_25,
	q_b_89,
	q_b_26,
	q_b_90,
	q_b_27,
	q_b_91,
	q_b_28,
	q_b_92,
	q_b_29,
	q_b_93,
	q_b_30,
	q_b_94,
	q_b_31,
	q_b_95,
	q_b_40,
	q_b_104,
	q_b_41,
	q_b_105,
	q_b_42,
	q_b_106,
	q_b_43,
	q_b_107,
	q_b_44,
	q_b_108,
	q_b_45,
	q_b_109,
	q_b_46,
	q_b_110,
	q_b_47,
	q_b_111,
	q_b_56,
	q_b_120,
	q_b_57,
	q_b_121,
	q_b_58,
	q_b_122,
	q_b_59,
	q_b_123,
	q_b_60,
	q_b_124,
	q_b_61,
	q_b_125,
	q_b_62,
	q_b_126,
	q_b_63,
	q_b_127,
	clk_0,
	clk_1,
	dataout_0,
	dataout_01,
	dataout_02,
	dataout_03,
	dataout_04,
	dataout_05,
	dataout_06,
	dataout_07,
	dataout_08,
	dataout_09,
	dataout_010,
	dataout_011,
	dataout_012,
	dataout_013,
	dataout_014,
	dataout_015,
	dataout_016,
	dataout_017,
	dataout_018,
	dataout_019,
	dataout_020,
	dataout_021,
	dataout_022,
	dataout_023,
	dqs_delay_ctrl_0,
	dqs_delay_ctrl_1,
	dqs_delay_ctrl_2,
	dqs_delay_ctrl_3,
	dqs_delay_ctrl_4,
	dqs_delay_ctrl_5,
	wire_output_dq_0_output_ddio_out_inst_dataout,
	wire_output_dq_0_output_ddio_out_inst_dataout1,
	wire_output_dq_0_output_ddio_out_inst_dataout2,
	wire_output_dq_0_output_ddio_out_inst_dataout3,
	do_read_r,
	mem_clk_buf_in_0,
	mem_clk_n_buf_in_0,
	wire_bidir_dq_0_output_ddio_out_inst_dataout,
	wire_bidir_dq_1_output_ddio_out_inst_dataout,
	wire_bidir_dq_2_output_ddio_out_inst_dataout,
	wire_bidir_dq_3_output_ddio_out_inst_dataout,
	wire_bidir_dq_4_output_ddio_out_inst_dataout,
	wire_bidir_dq_5_output_ddio_out_inst_dataout,
	wire_bidir_dq_6_output_ddio_out_inst_dataout,
	wire_bidir_dq_7_output_ddio_out_inst_dataout,
	wire_bidir_dq_0_output_ddio_out_inst_dataout1,
	wire_bidir_dq_1_output_ddio_out_inst_dataout1,
	wire_bidir_dq_2_output_ddio_out_inst_dataout1,
	wire_bidir_dq_3_output_ddio_out_inst_dataout1,
	wire_bidir_dq_4_output_ddio_out_inst_dataout1,
	wire_bidir_dq_5_output_ddio_out_inst_dataout1,
	wire_bidir_dq_6_output_ddio_out_inst_dataout1,
	wire_bidir_dq_7_output_ddio_out_inst_dataout1,
	wire_bidir_dq_0_output_ddio_out_inst_dataout2,
	wire_bidir_dq_1_output_ddio_out_inst_dataout2,
	wire_bidir_dq_2_output_ddio_out_inst_dataout2,
	wire_bidir_dq_3_output_ddio_out_inst_dataout2,
	wire_bidir_dq_4_output_ddio_out_inst_dataout2,
	wire_bidir_dq_5_output_ddio_out_inst_dataout2,
	wire_bidir_dq_6_output_ddio_out_inst_dataout2,
	wire_bidir_dq_7_output_ddio_out_inst_dataout2,
	wire_bidir_dq_0_output_ddio_out_inst_dataout3,
	wire_bidir_dq_1_output_ddio_out_inst_dataout3,
	wire_bidir_dq_2_output_ddio_out_inst_dataout3,
	wire_bidir_dq_3_output_ddio_out_inst_dataout3,
	wire_bidir_dq_4_output_ddio_out_inst_dataout3,
	wire_bidir_dq_5_output_ddio_out_inst_dataout3,
	wire_bidir_dq_6_output_ddio_out_inst_dataout3,
	wire_bidir_dq_7_output_ddio_out_inst_dataout3,
	dqs_pseudo_diff_out_0,
	dqsn_pseudo_diff_out_0,
	dqs_pseudo_diff_out_1,
	dqsn_pseudo_diff_out_1,
	dqs_pseudo_diff_out_2,
	dqsn_pseudo_diff_out_2,
	dqs_pseudo_diff_out_3,
	dqsn_pseudo_diff_out_3,
	dq_datain_0,
	dq_datain_1,
	dq_datain_2,
	dq_datain_3,
	dq_datain_4,
	dq_datain_5,
	dq_datain_6,
	dq_datain_7,
	dq_datain_8,
	dq_datain_9,
	dq_datain_10,
	dq_datain_11,
	dq_datain_12,
	dq_datain_13,
	dq_datain_14,
	dq_datain_15,
	dq_datain_16,
	dq_datain_17,
	dq_datain_18,
	dq_datain_19,
	dq_datain_20,
	dq_datain_21,
	dq_datain_22,
	dq_datain_23,
	dq_datain_24,
	dq_datain_25,
	dq_datain_26,
	dq_datain_27,
	dq_datain_28,
	dq_datain_29,
	dq_datain_30,
	dq_datain_31,
	dqs_buffered_0,
	dqs_buffered_1,
	dqs_buffered_2,
	dqs_buffered_3,
	q_b_961,
	q_b_321,
	q_b_641,
	q_b_01,
	q_b_971,
	q_b_331,
	q_b_651,
	q_b_128,
	q_b_981,
	q_b_341,
	q_b_661,
	q_b_210,
	q_b_991,
	q_b_351,
	q_b_671,
	q_b_310,
	q_b_1001,
	q_b_361,
	q_b_681,
	q_b_410,
	q_b_1011,
	q_b_371,
	q_b_691,
	q_b_510,
	q_b_1021,
	q_b_381,
	q_b_701,
	q_b_610,
	q_b_1031,
	q_b_391,
	q_b_711,
	q_b_710,
	q_b_1041,
	q_b_401,
	q_b_721,
	q_b_810,
	q_b_1051,
	q_b_411,
	q_b_731,
	q_b_910,
	q_b_1061,
	q_b_421,
	q_b_741,
	q_b_1010,
	q_b_1071,
	q_b_431,
	q_b_751,
	q_b_1110,
	q_b_1081,
	q_b_441,
	q_b_761,
	q_b_129,
	q_b_1091,
	q_b_451,
	q_b_771,
	q_b_131,
	q_b_1101,
	q_b_461,
	q_b_781,
	q_b_141,
	q_b_1111,
	q_b_471,
	q_b_791,
	q_b_151,
	q_b_1121,
	q_b_481,
	q_b_801,
	q_b_161,
	q_b_1131,
	q_b_491,
	q_b_811,
	q_b_171,
	q_b_1141,
	q_b_501,
	q_b_821,
	q_b_181,
	q_b_1151,
	q_b_511,
	q_b_831,
	q_b_191,
	q_b_1161,
	q_b_521,
	q_b_841,
	q_b_201,
	q_b_1171,
	q_b_531,
	q_b_851,
	q_b_211,
	q_b_1181,
	q_b_541,
	q_b_861,
	q_b_221,
	q_b_1191,
	q_b_551,
	q_b_871,
	q_b_231,
	q_b_1201,
	q_b_561,
	q_b_881,
	q_b_241,
	q_b_1211,
	q_b_571,
	q_b_891,
	q_b_251,
	q_b_1221,
	q_b_581,
	q_b_901,
	q_b_261,
	q_b_1231,
	q_b_591,
	q_b_911,
	q_b_271,
	q_b_1241,
	q_b_601,
	q_b_921,
	q_b_281,
	q_b_1251,
	q_b_611,
	q_b_931,
	q_b_291,
	q_b_1261,
	q_b_621,
	q_b_941,
	q_b_301,
	q_b_1271,
	q_b_631,
	q_b_951,
	q_b_311,
	fb_clk,
	ctl_rdata_valid_0,
	reset_request_n,
	ctl_init_fail,
	ctl_init_success,
	reset_phy_clk_1x_n,
	rdwr_data_valid_r,
	doing_read,
	bidir_dq_0_oe_ff_inst,
	bidir_dq_1_oe_ff_inst,
	bidir_dq_2_oe_ff_inst,
	bidir_dq_3_oe_ff_inst,
	bidir_dq_4_oe_ff_inst,
	bidir_dq_5_oe_ff_inst,
	bidir_dq_6_oe_ff_inst,
	bidir_dq_7_oe_ff_inst,
	bidir_dq_0_oe_ff_inst1,
	bidir_dq_1_oe_ff_inst1,
	bidir_dq_2_oe_ff_inst1,
	bidir_dq_3_oe_ff_inst1,
	bidir_dq_4_oe_ff_inst1,
	bidir_dq_5_oe_ff_inst1,
	bidir_dq_6_oe_ff_inst1,
	bidir_dq_7_oe_ff_inst1,
	bidir_dq_0_oe_ff_inst2,
	bidir_dq_1_oe_ff_inst2,
	bidir_dq_2_oe_ff_inst2,
	bidir_dq_3_oe_ff_inst2,
	bidir_dq_4_oe_ff_inst2,
	bidir_dq_5_oe_ff_inst2,
	bidir_dq_6_oe_ff_inst2,
	bidir_dq_7_oe_ff_inst2,
	bidir_dq_0_oe_ff_inst3,
	bidir_dq_1_oe_ff_inst3,
	bidir_dq_2_oe_ff_inst3,
	bidir_dq_3_oe_ff_inst3,
	bidir_dq_4_oe_ff_inst3,
	bidir_dq_5_oe_ff_inst3,
	bidir_dq_6_oe_ff_inst3,
	bidir_dq_7_oe_ff_inst3,
	dqs_0_oe_ff_inst,
	dqs_0_oe_ff_inst1,
	dqs_0_oe_ff_inst2,
	dqs_0_oe_ff_inst3,
	dqsn_0_oe_ff_inst,
	dqsn_0_oe_ff_inst1,
	dqsn_0_oe_ff_inst2,
	dqsn_0_oe_ff_inst3,
	wd_lat_2,
	wd_lat_1,
	wd_lat_0,
	wd_lat_3,
	wd_lat_4,
	afi_cs_n_1,
	int_cke_r_0,
	afi_addr_0,
	afi_addr_1,
	afi_addr_2,
	afi_addr_3,
	afi_addr_4,
	afi_addr_5,
	afi_addr_6,
	afi_addr_7,
	afi_addr_8,
	afi_addr_9,
	afi_addr_10,
	afi_addr_11,
	afi_addr_12,
	afi_addr_13,
	afi_ba_0,
	afi_ba_1,
	afi_ba_2,
	afi_ras_n_0,
	afi_cas_n_0,
	afi_we_n_0,
	afi_dm_4,
	afi_dm_12,
	afi_dm_0,
	afi_dm_8,
	afi_dm_5,
	afi_dm_13,
	afi_dm_1,
	afi_dm_9,
	afi_dm_6,
	afi_dm_14,
	afi_dm_2,
	afi_dm_10,
	afi_dm_7,
	afi_dm_15,
	afi_dm_3,
	afi_dm_11,
	int_wdata_valid,
	int_dqs_burst,
	int_dqs_burst_hr,
	GND_port,
	global_reset_n,
	pll_ref_clk,
	soft_reset_n)/* synthesis synthesis_greybox=0 */;
output 	q_b_0;
output 	q_b_64;
output 	q_b_1;
output 	q_b_65;
output 	q_b_2;
output 	q_b_66;
output 	q_b_3;
output 	q_b_67;
output 	q_b_4;
output 	q_b_68;
output 	q_b_5;
output 	q_b_69;
output 	q_b_6;
output 	q_b_70;
output 	q_b_7;
output 	q_b_71;
output 	q_b_16;
output 	q_b_80;
output 	q_b_17;
output 	q_b_81;
output 	q_b_18;
output 	q_b_82;
output 	q_b_19;
output 	q_b_83;
output 	q_b_20;
output 	q_b_84;
output 	q_b_21;
output 	q_b_85;
output 	q_b_22;
output 	q_b_86;
output 	q_b_23;
output 	q_b_87;
output 	q_b_32;
output 	q_b_96;
output 	q_b_33;
output 	q_b_97;
output 	q_b_34;
output 	q_b_98;
output 	q_b_35;
output 	q_b_99;
output 	q_b_36;
output 	q_b_100;
output 	q_b_37;
output 	q_b_101;
output 	q_b_38;
output 	q_b_102;
output 	q_b_39;
output 	q_b_103;
output 	q_b_48;
output 	q_b_112;
output 	q_b_49;
output 	q_b_113;
output 	q_b_50;
output 	q_b_114;
output 	q_b_51;
output 	q_b_115;
output 	q_b_52;
output 	q_b_116;
output 	q_b_53;
output 	q_b_117;
output 	q_b_54;
output 	q_b_118;
output 	q_b_55;
output 	q_b_119;
output 	q_b_8;
output 	q_b_72;
output 	q_b_9;
output 	q_b_73;
output 	q_b_10;
output 	q_b_74;
output 	q_b_11;
output 	q_b_75;
output 	q_b_12;
output 	q_b_76;
output 	q_b_13;
output 	q_b_77;
output 	q_b_14;
output 	q_b_78;
output 	q_b_15;
output 	q_b_79;
output 	q_b_24;
output 	q_b_88;
output 	q_b_25;
output 	q_b_89;
output 	q_b_26;
output 	q_b_90;
output 	q_b_27;
output 	q_b_91;
output 	q_b_28;
output 	q_b_92;
output 	q_b_29;
output 	q_b_93;
output 	q_b_30;
output 	q_b_94;
output 	q_b_31;
output 	q_b_95;
output 	q_b_40;
output 	q_b_104;
output 	q_b_41;
output 	q_b_105;
output 	q_b_42;
output 	q_b_106;
output 	q_b_43;
output 	q_b_107;
output 	q_b_44;
output 	q_b_108;
output 	q_b_45;
output 	q_b_109;
output 	q_b_46;
output 	q_b_110;
output 	q_b_47;
output 	q_b_111;
output 	q_b_56;
output 	q_b_120;
output 	q_b_57;
output 	q_b_121;
output 	q_b_58;
output 	q_b_122;
output 	q_b_59;
output 	q_b_123;
output 	q_b_60;
output 	q_b_124;
output 	q_b_61;
output 	q_b_125;
output 	q_b_62;
output 	q_b_126;
output 	q_b_63;
output 	q_b_127;
output 	clk_0;
output 	clk_1;
output 	dataout_0;
output 	dataout_01;
output 	dataout_02;
output 	dataout_03;
output 	dataout_04;
output 	dataout_05;
output 	dataout_06;
output 	dataout_07;
output 	dataout_08;
output 	dataout_09;
output 	dataout_010;
output 	dataout_011;
output 	dataout_012;
output 	dataout_013;
output 	dataout_014;
output 	dataout_015;
output 	dataout_016;
output 	dataout_017;
output 	dataout_018;
output 	dataout_019;
output 	dataout_020;
output 	dataout_021;
output 	dataout_022;
output 	dataout_023;
output 	dqs_delay_ctrl_0;
output 	dqs_delay_ctrl_1;
output 	dqs_delay_ctrl_2;
output 	dqs_delay_ctrl_3;
output 	dqs_delay_ctrl_4;
output 	dqs_delay_ctrl_5;
output 	wire_output_dq_0_output_ddio_out_inst_dataout;
output 	wire_output_dq_0_output_ddio_out_inst_dataout1;
output 	wire_output_dq_0_output_ddio_out_inst_dataout2;
output 	wire_output_dq_0_output_ddio_out_inst_dataout3;
input 	do_read_r;
output 	mem_clk_buf_in_0;
output 	mem_clk_n_buf_in_0;
output 	wire_bidir_dq_0_output_ddio_out_inst_dataout;
output 	wire_bidir_dq_1_output_ddio_out_inst_dataout;
output 	wire_bidir_dq_2_output_ddio_out_inst_dataout;
output 	wire_bidir_dq_3_output_ddio_out_inst_dataout;
output 	wire_bidir_dq_4_output_ddio_out_inst_dataout;
output 	wire_bidir_dq_5_output_ddio_out_inst_dataout;
output 	wire_bidir_dq_6_output_ddio_out_inst_dataout;
output 	wire_bidir_dq_7_output_ddio_out_inst_dataout;
output 	wire_bidir_dq_0_output_ddio_out_inst_dataout1;
output 	wire_bidir_dq_1_output_ddio_out_inst_dataout1;
output 	wire_bidir_dq_2_output_ddio_out_inst_dataout1;
output 	wire_bidir_dq_3_output_ddio_out_inst_dataout1;
output 	wire_bidir_dq_4_output_ddio_out_inst_dataout1;
output 	wire_bidir_dq_5_output_ddio_out_inst_dataout1;
output 	wire_bidir_dq_6_output_ddio_out_inst_dataout1;
output 	wire_bidir_dq_7_output_ddio_out_inst_dataout1;
output 	wire_bidir_dq_0_output_ddio_out_inst_dataout2;
output 	wire_bidir_dq_1_output_ddio_out_inst_dataout2;
output 	wire_bidir_dq_2_output_ddio_out_inst_dataout2;
output 	wire_bidir_dq_3_output_ddio_out_inst_dataout2;
output 	wire_bidir_dq_4_output_ddio_out_inst_dataout2;
output 	wire_bidir_dq_5_output_ddio_out_inst_dataout2;
output 	wire_bidir_dq_6_output_ddio_out_inst_dataout2;
output 	wire_bidir_dq_7_output_ddio_out_inst_dataout2;
output 	wire_bidir_dq_0_output_ddio_out_inst_dataout3;
output 	wire_bidir_dq_1_output_ddio_out_inst_dataout3;
output 	wire_bidir_dq_2_output_ddio_out_inst_dataout3;
output 	wire_bidir_dq_3_output_ddio_out_inst_dataout3;
output 	wire_bidir_dq_4_output_ddio_out_inst_dataout3;
output 	wire_bidir_dq_5_output_ddio_out_inst_dataout3;
output 	wire_bidir_dq_6_output_ddio_out_inst_dataout3;
output 	wire_bidir_dq_7_output_ddio_out_inst_dataout3;
output 	dqs_pseudo_diff_out_0;
output 	dqsn_pseudo_diff_out_0;
output 	dqs_pseudo_diff_out_1;
output 	dqsn_pseudo_diff_out_1;
output 	dqs_pseudo_diff_out_2;
output 	dqsn_pseudo_diff_out_2;
output 	dqs_pseudo_diff_out_3;
output 	dqsn_pseudo_diff_out_3;
input 	dq_datain_0;
input 	dq_datain_1;
input 	dq_datain_2;
input 	dq_datain_3;
input 	dq_datain_4;
input 	dq_datain_5;
input 	dq_datain_6;
input 	dq_datain_7;
input 	dq_datain_8;
input 	dq_datain_9;
input 	dq_datain_10;
input 	dq_datain_11;
input 	dq_datain_12;
input 	dq_datain_13;
input 	dq_datain_14;
input 	dq_datain_15;
input 	dq_datain_16;
input 	dq_datain_17;
input 	dq_datain_18;
input 	dq_datain_19;
input 	dq_datain_20;
input 	dq_datain_21;
input 	dq_datain_22;
input 	dq_datain_23;
input 	dq_datain_24;
input 	dq_datain_25;
input 	dq_datain_26;
input 	dq_datain_27;
input 	dq_datain_28;
input 	dq_datain_29;
input 	dq_datain_30;
input 	dq_datain_31;
input 	dqs_buffered_0;
input 	dqs_buffered_1;
input 	dqs_buffered_2;
input 	dqs_buffered_3;
input 	q_b_961;
input 	q_b_321;
input 	q_b_641;
input 	q_b_01;
input 	q_b_971;
input 	q_b_331;
input 	q_b_651;
input 	q_b_128;
input 	q_b_981;
input 	q_b_341;
input 	q_b_661;
input 	q_b_210;
input 	q_b_991;
input 	q_b_351;
input 	q_b_671;
input 	q_b_310;
input 	q_b_1001;
input 	q_b_361;
input 	q_b_681;
input 	q_b_410;
input 	q_b_1011;
input 	q_b_371;
input 	q_b_691;
input 	q_b_510;
input 	q_b_1021;
input 	q_b_381;
input 	q_b_701;
input 	q_b_610;
input 	q_b_1031;
input 	q_b_391;
input 	q_b_711;
input 	q_b_710;
input 	q_b_1041;
input 	q_b_401;
input 	q_b_721;
input 	q_b_810;
input 	q_b_1051;
input 	q_b_411;
input 	q_b_731;
input 	q_b_910;
input 	q_b_1061;
input 	q_b_421;
input 	q_b_741;
input 	q_b_1010;
input 	q_b_1071;
input 	q_b_431;
input 	q_b_751;
input 	q_b_1110;
input 	q_b_1081;
input 	q_b_441;
input 	q_b_761;
input 	q_b_129;
input 	q_b_1091;
input 	q_b_451;
input 	q_b_771;
input 	q_b_131;
input 	q_b_1101;
input 	q_b_461;
input 	q_b_781;
input 	q_b_141;
input 	q_b_1111;
input 	q_b_471;
input 	q_b_791;
input 	q_b_151;
input 	q_b_1121;
input 	q_b_481;
input 	q_b_801;
input 	q_b_161;
input 	q_b_1131;
input 	q_b_491;
input 	q_b_811;
input 	q_b_171;
input 	q_b_1141;
input 	q_b_501;
input 	q_b_821;
input 	q_b_181;
input 	q_b_1151;
input 	q_b_511;
input 	q_b_831;
input 	q_b_191;
input 	q_b_1161;
input 	q_b_521;
input 	q_b_841;
input 	q_b_201;
input 	q_b_1171;
input 	q_b_531;
input 	q_b_851;
input 	q_b_211;
input 	q_b_1181;
input 	q_b_541;
input 	q_b_861;
input 	q_b_221;
input 	q_b_1191;
input 	q_b_551;
input 	q_b_871;
input 	q_b_231;
input 	q_b_1201;
input 	q_b_561;
input 	q_b_881;
input 	q_b_241;
input 	q_b_1211;
input 	q_b_571;
input 	q_b_891;
input 	q_b_251;
input 	q_b_1221;
input 	q_b_581;
input 	q_b_901;
input 	q_b_261;
input 	q_b_1231;
input 	q_b_591;
input 	q_b_911;
input 	q_b_271;
input 	q_b_1241;
input 	q_b_601;
input 	q_b_921;
input 	q_b_281;
input 	q_b_1251;
input 	q_b_611;
input 	q_b_931;
input 	q_b_291;
input 	q_b_1261;
input 	q_b_621;
input 	q_b_941;
input 	q_b_301;
input 	q_b_1271;
input 	q_b_631;
input 	q_b_951;
input 	q_b_311;
input 	fb_clk;
output 	ctl_rdata_valid_0;
output 	reset_request_n;
output 	ctl_init_fail;
output 	ctl_init_success;
output 	reset_phy_clk_1x_n;
input 	rdwr_data_valid_r;
input 	doing_read;
output 	bidir_dq_0_oe_ff_inst;
output 	bidir_dq_1_oe_ff_inst;
output 	bidir_dq_2_oe_ff_inst;
output 	bidir_dq_3_oe_ff_inst;
output 	bidir_dq_4_oe_ff_inst;
output 	bidir_dq_5_oe_ff_inst;
output 	bidir_dq_6_oe_ff_inst;
output 	bidir_dq_7_oe_ff_inst;
output 	bidir_dq_0_oe_ff_inst1;
output 	bidir_dq_1_oe_ff_inst1;
output 	bidir_dq_2_oe_ff_inst1;
output 	bidir_dq_3_oe_ff_inst1;
output 	bidir_dq_4_oe_ff_inst1;
output 	bidir_dq_5_oe_ff_inst1;
output 	bidir_dq_6_oe_ff_inst1;
output 	bidir_dq_7_oe_ff_inst1;
output 	bidir_dq_0_oe_ff_inst2;
output 	bidir_dq_1_oe_ff_inst2;
output 	bidir_dq_2_oe_ff_inst2;
output 	bidir_dq_3_oe_ff_inst2;
output 	bidir_dq_4_oe_ff_inst2;
output 	bidir_dq_5_oe_ff_inst2;
output 	bidir_dq_6_oe_ff_inst2;
output 	bidir_dq_7_oe_ff_inst2;
output 	bidir_dq_0_oe_ff_inst3;
output 	bidir_dq_1_oe_ff_inst3;
output 	bidir_dq_2_oe_ff_inst3;
output 	bidir_dq_3_oe_ff_inst3;
output 	bidir_dq_4_oe_ff_inst3;
output 	bidir_dq_5_oe_ff_inst3;
output 	bidir_dq_6_oe_ff_inst3;
output 	bidir_dq_7_oe_ff_inst3;
output 	dqs_0_oe_ff_inst;
output 	dqs_0_oe_ff_inst1;
output 	dqs_0_oe_ff_inst2;
output 	dqs_0_oe_ff_inst3;
output 	dqsn_0_oe_ff_inst;
output 	dqsn_0_oe_ff_inst1;
output 	dqsn_0_oe_ff_inst2;
output 	dqsn_0_oe_ff_inst3;
output 	wd_lat_2;
output 	wd_lat_1;
output 	wd_lat_0;
output 	wd_lat_3;
output 	wd_lat_4;
input 	afi_cs_n_1;
input 	int_cke_r_0;
input 	afi_addr_0;
input 	afi_addr_1;
input 	afi_addr_2;
input 	afi_addr_3;
input 	afi_addr_4;
input 	afi_addr_5;
input 	afi_addr_6;
input 	afi_addr_7;
input 	afi_addr_8;
input 	afi_addr_9;
input 	afi_addr_10;
input 	afi_addr_11;
input 	afi_addr_12;
input 	afi_addr_13;
input 	afi_ba_0;
input 	afi_ba_1;
input 	afi_ba_2;
input 	afi_ras_n_0;
input 	afi_cas_n_0;
input 	afi_we_n_0;
input 	afi_dm_4;
input 	afi_dm_12;
input 	afi_dm_0;
input 	afi_dm_8;
input 	afi_dm_5;
input 	afi_dm_13;
input 	afi_dm_1;
input 	afi_dm_9;
input 	afi_dm_6;
input 	afi_dm_14;
input 	afi_dm_2;
input 	afi_dm_10;
input 	afi_dm_7;
input 	afi_dm_15;
input 	afi_dm_3;
input 	afi_dm_11;
input 	int_wdata_valid;
input 	int_dqs_burst;
input 	int_dqs_burst_hr;
input 	GND_port;
input 	global_reset_n;
input 	pll_ref_clk;
input 	soft_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_ddr3_int_phy_alt_mem_phy ddr3_int_phy_alt_mem_phy_inst(
	.q_b_0(q_b_0),
	.q_b_64(q_b_64),
	.q_b_1(q_b_1),
	.q_b_65(q_b_65),
	.q_b_2(q_b_2),
	.q_b_66(q_b_66),
	.q_b_3(q_b_3),
	.q_b_67(q_b_67),
	.q_b_4(q_b_4),
	.q_b_68(q_b_68),
	.q_b_5(q_b_5),
	.q_b_69(q_b_69),
	.q_b_6(q_b_6),
	.q_b_70(q_b_70),
	.q_b_7(q_b_7),
	.q_b_71(q_b_71),
	.q_b_16(q_b_16),
	.q_b_80(q_b_80),
	.q_b_17(q_b_17),
	.q_b_81(q_b_81),
	.q_b_18(q_b_18),
	.q_b_82(q_b_82),
	.q_b_19(q_b_19),
	.q_b_83(q_b_83),
	.q_b_20(q_b_20),
	.q_b_84(q_b_84),
	.q_b_21(q_b_21),
	.q_b_85(q_b_85),
	.q_b_22(q_b_22),
	.q_b_86(q_b_86),
	.q_b_23(q_b_23),
	.q_b_87(q_b_87),
	.q_b_32(q_b_32),
	.q_b_96(q_b_96),
	.q_b_33(q_b_33),
	.q_b_97(q_b_97),
	.q_b_34(q_b_34),
	.q_b_98(q_b_98),
	.q_b_35(q_b_35),
	.q_b_99(q_b_99),
	.q_b_36(q_b_36),
	.q_b_100(q_b_100),
	.q_b_37(q_b_37),
	.q_b_101(q_b_101),
	.q_b_38(q_b_38),
	.q_b_102(q_b_102),
	.q_b_39(q_b_39),
	.q_b_103(q_b_103),
	.q_b_48(q_b_48),
	.q_b_112(q_b_112),
	.q_b_49(q_b_49),
	.q_b_113(q_b_113),
	.q_b_50(q_b_50),
	.q_b_114(q_b_114),
	.q_b_51(q_b_51),
	.q_b_115(q_b_115),
	.q_b_52(q_b_52),
	.q_b_116(q_b_116),
	.q_b_53(q_b_53),
	.q_b_117(q_b_117),
	.q_b_54(q_b_54),
	.q_b_118(q_b_118),
	.q_b_55(q_b_55),
	.q_b_119(q_b_119),
	.q_b_8(q_b_8),
	.q_b_72(q_b_72),
	.q_b_9(q_b_9),
	.q_b_73(q_b_73),
	.q_b_10(q_b_10),
	.q_b_74(q_b_74),
	.q_b_11(q_b_11),
	.q_b_75(q_b_75),
	.q_b_12(q_b_12),
	.q_b_76(q_b_76),
	.q_b_13(q_b_13),
	.q_b_77(q_b_77),
	.q_b_14(q_b_14),
	.q_b_78(q_b_78),
	.q_b_15(q_b_15),
	.q_b_79(q_b_79),
	.q_b_24(q_b_24),
	.q_b_88(q_b_88),
	.q_b_25(q_b_25),
	.q_b_89(q_b_89),
	.q_b_26(q_b_26),
	.q_b_90(q_b_90),
	.q_b_27(q_b_27),
	.q_b_91(q_b_91),
	.q_b_28(q_b_28),
	.q_b_92(q_b_92),
	.q_b_29(q_b_29),
	.q_b_93(q_b_93),
	.q_b_30(q_b_30),
	.q_b_94(q_b_94),
	.q_b_31(q_b_31),
	.q_b_95(q_b_95),
	.q_b_40(q_b_40),
	.q_b_104(q_b_104),
	.q_b_41(q_b_41),
	.q_b_105(q_b_105),
	.q_b_42(q_b_42),
	.q_b_106(q_b_106),
	.q_b_43(q_b_43),
	.q_b_107(q_b_107),
	.q_b_44(q_b_44),
	.q_b_108(q_b_108),
	.q_b_45(q_b_45),
	.q_b_109(q_b_109),
	.q_b_46(q_b_46),
	.q_b_110(q_b_110),
	.q_b_47(q_b_47),
	.q_b_111(q_b_111),
	.q_b_56(q_b_56),
	.q_b_120(q_b_120),
	.q_b_57(q_b_57),
	.q_b_121(q_b_121),
	.q_b_58(q_b_58),
	.q_b_122(q_b_122),
	.q_b_59(q_b_59),
	.q_b_123(q_b_123),
	.q_b_60(q_b_60),
	.q_b_124(q_b_124),
	.q_b_61(q_b_61),
	.q_b_125(q_b_125),
	.q_b_62(q_b_62),
	.q_b_126(q_b_126),
	.q_b_63(q_b_63),
	.q_b_127(q_b_127),
	.clk_0(clk_0),
	.clk_1(clk_1),
	.dataout_0(dataout_0),
	.dataout_01(dataout_01),
	.dataout_02(dataout_02),
	.dataout_03(dataout_03),
	.dataout_04(dataout_04),
	.dataout_05(dataout_05),
	.dataout_06(dataout_06),
	.dataout_07(dataout_07),
	.dataout_08(dataout_08),
	.dataout_09(dataout_09),
	.dataout_010(dataout_010),
	.dataout_011(dataout_011),
	.dataout_012(dataout_012),
	.dataout_013(dataout_013),
	.dataout_014(dataout_014),
	.dataout_015(dataout_015),
	.dataout_016(dataout_016),
	.dataout_017(dataout_017),
	.dataout_018(dataout_018),
	.dataout_019(dataout_019),
	.dataout_020(dataout_020),
	.dataout_021(dataout_021),
	.dataout_022(dataout_022),
	.dataout_023(dataout_023),
	.dqs_delay_ctrl_0(dqs_delay_ctrl_0),
	.dqs_delay_ctrl_1(dqs_delay_ctrl_1),
	.dqs_delay_ctrl_2(dqs_delay_ctrl_2),
	.dqs_delay_ctrl_3(dqs_delay_ctrl_3),
	.dqs_delay_ctrl_4(dqs_delay_ctrl_4),
	.dqs_delay_ctrl_5(dqs_delay_ctrl_5),
	.wire_output_dq_0_output_ddio_out_inst_dataout(wire_output_dq_0_output_ddio_out_inst_dataout),
	.wire_output_dq_0_output_ddio_out_inst_dataout1(wire_output_dq_0_output_ddio_out_inst_dataout1),
	.wire_output_dq_0_output_ddio_out_inst_dataout2(wire_output_dq_0_output_ddio_out_inst_dataout2),
	.wire_output_dq_0_output_ddio_out_inst_dataout3(wire_output_dq_0_output_ddio_out_inst_dataout3),
	.do_read_r(do_read_r),
	.mem_clk_buf_in_0(mem_clk_buf_in_0),
	.mem_clk_n_buf_in_0(mem_clk_n_buf_in_0),
	.wire_bidir_dq_0_output_ddio_out_inst_dataout(wire_bidir_dq_0_output_ddio_out_inst_dataout),
	.wire_bidir_dq_1_output_ddio_out_inst_dataout(wire_bidir_dq_1_output_ddio_out_inst_dataout),
	.wire_bidir_dq_2_output_ddio_out_inst_dataout(wire_bidir_dq_2_output_ddio_out_inst_dataout),
	.wire_bidir_dq_3_output_ddio_out_inst_dataout(wire_bidir_dq_3_output_ddio_out_inst_dataout),
	.wire_bidir_dq_4_output_ddio_out_inst_dataout(wire_bidir_dq_4_output_ddio_out_inst_dataout),
	.wire_bidir_dq_5_output_ddio_out_inst_dataout(wire_bidir_dq_5_output_ddio_out_inst_dataout),
	.wire_bidir_dq_6_output_ddio_out_inst_dataout(wire_bidir_dq_6_output_ddio_out_inst_dataout),
	.wire_bidir_dq_7_output_ddio_out_inst_dataout(wire_bidir_dq_7_output_ddio_out_inst_dataout),
	.wire_bidir_dq_0_output_ddio_out_inst_dataout1(wire_bidir_dq_0_output_ddio_out_inst_dataout1),
	.wire_bidir_dq_1_output_ddio_out_inst_dataout1(wire_bidir_dq_1_output_ddio_out_inst_dataout1),
	.wire_bidir_dq_2_output_ddio_out_inst_dataout1(wire_bidir_dq_2_output_ddio_out_inst_dataout1),
	.wire_bidir_dq_3_output_ddio_out_inst_dataout1(wire_bidir_dq_3_output_ddio_out_inst_dataout1),
	.wire_bidir_dq_4_output_ddio_out_inst_dataout1(wire_bidir_dq_4_output_ddio_out_inst_dataout1),
	.wire_bidir_dq_5_output_ddio_out_inst_dataout1(wire_bidir_dq_5_output_ddio_out_inst_dataout1),
	.wire_bidir_dq_6_output_ddio_out_inst_dataout1(wire_bidir_dq_6_output_ddio_out_inst_dataout1),
	.wire_bidir_dq_7_output_ddio_out_inst_dataout1(wire_bidir_dq_7_output_ddio_out_inst_dataout1),
	.wire_bidir_dq_0_output_ddio_out_inst_dataout2(wire_bidir_dq_0_output_ddio_out_inst_dataout2),
	.wire_bidir_dq_1_output_ddio_out_inst_dataout2(wire_bidir_dq_1_output_ddio_out_inst_dataout2),
	.wire_bidir_dq_2_output_ddio_out_inst_dataout2(wire_bidir_dq_2_output_ddio_out_inst_dataout2),
	.wire_bidir_dq_3_output_ddio_out_inst_dataout2(wire_bidir_dq_3_output_ddio_out_inst_dataout2),
	.wire_bidir_dq_4_output_ddio_out_inst_dataout2(wire_bidir_dq_4_output_ddio_out_inst_dataout2),
	.wire_bidir_dq_5_output_ddio_out_inst_dataout2(wire_bidir_dq_5_output_ddio_out_inst_dataout2),
	.wire_bidir_dq_6_output_ddio_out_inst_dataout2(wire_bidir_dq_6_output_ddio_out_inst_dataout2),
	.wire_bidir_dq_7_output_ddio_out_inst_dataout2(wire_bidir_dq_7_output_ddio_out_inst_dataout2),
	.wire_bidir_dq_0_output_ddio_out_inst_dataout3(wire_bidir_dq_0_output_ddio_out_inst_dataout3),
	.wire_bidir_dq_1_output_ddio_out_inst_dataout3(wire_bidir_dq_1_output_ddio_out_inst_dataout3),
	.wire_bidir_dq_2_output_ddio_out_inst_dataout3(wire_bidir_dq_2_output_ddio_out_inst_dataout3),
	.wire_bidir_dq_3_output_ddio_out_inst_dataout3(wire_bidir_dq_3_output_ddio_out_inst_dataout3),
	.wire_bidir_dq_4_output_ddio_out_inst_dataout3(wire_bidir_dq_4_output_ddio_out_inst_dataout3),
	.wire_bidir_dq_5_output_ddio_out_inst_dataout3(wire_bidir_dq_5_output_ddio_out_inst_dataout3),
	.wire_bidir_dq_6_output_ddio_out_inst_dataout3(wire_bidir_dq_6_output_ddio_out_inst_dataout3),
	.wire_bidir_dq_7_output_ddio_out_inst_dataout3(wire_bidir_dq_7_output_ddio_out_inst_dataout3),
	.dqs_pseudo_diff_out_0(dqs_pseudo_diff_out_0),
	.dqsn_pseudo_diff_out_0(dqsn_pseudo_diff_out_0),
	.dqs_pseudo_diff_out_1(dqs_pseudo_diff_out_1),
	.dqsn_pseudo_diff_out_1(dqsn_pseudo_diff_out_1),
	.dqs_pseudo_diff_out_2(dqs_pseudo_diff_out_2),
	.dqsn_pseudo_diff_out_2(dqsn_pseudo_diff_out_2),
	.dqs_pseudo_diff_out_3(dqs_pseudo_diff_out_3),
	.dqsn_pseudo_diff_out_3(dqsn_pseudo_diff_out_3),
	.dq_datain_0(dq_datain_0),
	.dq_datain_1(dq_datain_1),
	.dq_datain_2(dq_datain_2),
	.dq_datain_3(dq_datain_3),
	.dq_datain_4(dq_datain_4),
	.dq_datain_5(dq_datain_5),
	.dq_datain_6(dq_datain_6),
	.dq_datain_7(dq_datain_7),
	.dq_datain_8(dq_datain_8),
	.dq_datain_9(dq_datain_9),
	.dq_datain_10(dq_datain_10),
	.dq_datain_11(dq_datain_11),
	.dq_datain_12(dq_datain_12),
	.dq_datain_13(dq_datain_13),
	.dq_datain_14(dq_datain_14),
	.dq_datain_15(dq_datain_15),
	.dq_datain_16(dq_datain_16),
	.dq_datain_17(dq_datain_17),
	.dq_datain_18(dq_datain_18),
	.dq_datain_19(dq_datain_19),
	.dq_datain_20(dq_datain_20),
	.dq_datain_21(dq_datain_21),
	.dq_datain_22(dq_datain_22),
	.dq_datain_23(dq_datain_23),
	.dq_datain_24(dq_datain_24),
	.dq_datain_25(dq_datain_25),
	.dq_datain_26(dq_datain_26),
	.dq_datain_27(dq_datain_27),
	.dq_datain_28(dq_datain_28),
	.dq_datain_29(dq_datain_29),
	.dq_datain_30(dq_datain_30),
	.dq_datain_31(dq_datain_31),
	.dqs_buffered_0(dqs_buffered_0),
	.dqs_buffered_1(dqs_buffered_1),
	.dqs_buffered_2(dqs_buffered_2),
	.dqs_buffered_3(dqs_buffered_3),
	.q_b_961(q_b_961),
	.q_b_321(q_b_321),
	.q_b_641(q_b_641),
	.q_b_01(q_b_01),
	.q_b_971(q_b_971),
	.q_b_331(q_b_331),
	.q_b_651(q_b_651),
	.q_b_128(q_b_128),
	.q_b_981(q_b_981),
	.q_b_341(q_b_341),
	.q_b_661(q_b_661),
	.q_b_210(q_b_210),
	.q_b_991(q_b_991),
	.q_b_351(q_b_351),
	.q_b_671(q_b_671),
	.q_b_310(q_b_310),
	.q_b_1001(q_b_1001),
	.q_b_361(q_b_361),
	.q_b_681(q_b_681),
	.q_b_410(q_b_410),
	.q_b_1011(q_b_1011),
	.q_b_371(q_b_371),
	.q_b_691(q_b_691),
	.q_b_510(q_b_510),
	.q_b_1021(q_b_1021),
	.q_b_381(q_b_381),
	.q_b_701(q_b_701),
	.q_b_610(q_b_610),
	.q_b_1031(q_b_1031),
	.q_b_391(q_b_391),
	.q_b_711(q_b_711),
	.q_b_710(q_b_710),
	.q_b_1041(q_b_1041),
	.q_b_401(q_b_401),
	.q_b_721(q_b_721),
	.q_b_810(q_b_810),
	.q_b_1051(q_b_1051),
	.q_b_411(q_b_411),
	.q_b_731(q_b_731),
	.q_b_910(q_b_910),
	.q_b_1061(q_b_1061),
	.q_b_421(q_b_421),
	.q_b_741(q_b_741),
	.q_b_1010(q_b_1010),
	.q_b_1071(q_b_1071),
	.q_b_431(q_b_431),
	.q_b_751(q_b_751),
	.q_b_1110(q_b_1110),
	.q_b_1081(q_b_1081),
	.q_b_441(q_b_441),
	.q_b_761(q_b_761),
	.q_b_129(q_b_129),
	.q_b_1091(q_b_1091),
	.q_b_451(q_b_451),
	.q_b_771(q_b_771),
	.q_b_131(q_b_131),
	.q_b_1101(q_b_1101),
	.q_b_461(q_b_461),
	.q_b_781(q_b_781),
	.q_b_141(q_b_141),
	.q_b_1111(q_b_1111),
	.q_b_471(q_b_471),
	.q_b_791(q_b_791),
	.q_b_151(q_b_151),
	.q_b_1121(q_b_1121),
	.q_b_481(q_b_481),
	.q_b_801(q_b_801),
	.q_b_161(q_b_161),
	.q_b_1131(q_b_1131),
	.q_b_491(q_b_491),
	.q_b_811(q_b_811),
	.q_b_171(q_b_171),
	.q_b_1141(q_b_1141),
	.q_b_501(q_b_501),
	.q_b_821(q_b_821),
	.q_b_181(q_b_181),
	.q_b_1151(q_b_1151),
	.q_b_511(q_b_511),
	.q_b_831(q_b_831),
	.q_b_191(q_b_191),
	.q_b_1161(q_b_1161),
	.q_b_521(q_b_521),
	.q_b_841(q_b_841),
	.q_b_201(q_b_201),
	.q_b_1171(q_b_1171),
	.q_b_531(q_b_531),
	.q_b_851(q_b_851),
	.q_b_211(q_b_211),
	.q_b_1181(q_b_1181),
	.q_b_541(q_b_541),
	.q_b_861(q_b_861),
	.q_b_221(q_b_221),
	.q_b_1191(q_b_1191),
	.q_b_551(q_b_551),
	.q_b_871(q_b_871),
	.q_b_231(q_b_231),
	.q_b_1201(q_b_1201),
	.q_b_561(q_b_561),
	.q_b_881(q_b_881),
	.q_b_241(q_b_241),
	.q_b_1211(q_b_1211),
	.q_b_571(q_b_571),
	.q_b_891(q_b_891),
	.q_b_251(q_b_251),
	.q_b_1221(q_b_1221),
	.q_b_581(q_b_581),
	.q_b_901(q_b_901),
	.q_b_261(q_b_261),
	.q_b_1231(q_b_1231),
	.q_b_591(q_b_591),
	.q_b_911(q_b_911),
	.q_b_271(q_b_271),
	.q_b_1241(q_b_1241),
	.q_b_601(q_b_601),
	.q_b_921(q_b_921),
	.q_b_281(q_b_281),
	.q_b_1251(q_b_1251),
	.q_b_611(q_b_611),
	.q_b_931(q_b_931),
	.q_b_291(q_b_291),
	.q_b_1261(q_b_1261),
	.q_b_621(q_b_621),
	.q_b_941(q_b_941),
	.q_b_301(q_b_301),
	.q_b_1271(q_b_1271),
	.q_b_631(q_b_631),
	.q_b_951(q_b_951),
	.q_b_311(q_b_311),
	.fb_clk(fb_clk),
	.ctl_rdata_valid_0(ctl_rdata_valid_0),
	.reset_request_n(reset_request_n),
	.ctl_init_fail(ctl_init_fail),
	.ctl_init_success(ctl_init_success),
	.reset_phy_clk_1x_n(reset_phy_clk_1x_n),
	.rdwr_data_valid_r(rdwr_data_valid_r),
	.doing_read(doing_read),
	.bidir_dq_0_oe_ff_inst(bidir_dq_0_oe_ff_inst),
	.bidir_dq_1_oe_ff_inst(bidir_dq_1_oe_ff_inst),
	.bidir_dq_2_oe_ff_inst(bidir_dq_2_oe_ff_inst),
	.bidir_dq_3_oe_ff_inst(bidir_dq_3_oe_ff_inst),
	.bidir_dq_4_oe_ff_inst(bidir_dq_4_oe_ff_inst),
	.bidir_dq_5_oe_ff_inst(bidir_dq_5_oe_ff_inst),
	.bidir_dq_6_oe_ff_inst(bidir_dq_6_oe_ff_inst),
	.bidir_dq_7_oe_ff_inst(bidir_dq_7_oe_ff_inst),
	.bidir_dq_0_oe_ff_inst1(bidir_dq_0_oe_ff_inst1),
	.bidir_dq_1_oe_ff_inst1(bidir_dq_1_oe_ff_inst1),
	.bidir_dq_2_oe_ff_inst1(bidir_dq_2_oe_ff_inst1),
	.bidir_dq_3_oe_ff_inst1(bidir_dq_3_oe_ff_inst1),
	.bidir_dq_4_oe_ff_inst1(bidir_dq_4_oe_ff_inst1),
	.bidir_dq_5_oe_ff_inst1(bidir_dq_5_oe_ff_inst1),
	.bidir_dq_6_oe_ff_inst1(bidir_dq_6_oe_ff_inst1),
	.bidir_dq_7_oe_ff_inst1(bidir_dq_7_oe_ff_inst1),
	.bidir_dq_0_oe_ff_inst2(bidir_dq_0_oe_ff_inst2),
	.bidir_dq_1_oe_ff_inst2(bidir_dq_1_oe_ff_inst2),
	.bidir_dq_2_oe_ff_inst2(bidir_dq_2_oe_ff_inst2),
	.bidir_dq_3_oe_ff_inst2(bidir_dq_3_oe_ff_inst2),
	.bidir_dq_4_oe_ff_inst2(bidir_dq_4_oe_ff_inst2),
	.bidir_dq_5_oe_ff_inst2(bidir_dq_5_oe_ff_inst2),
	.bidir_dq_6_oe_ff_inst2(bidir_dq_6_oe_ff_inst2),
	.bidir_dq_7_oe_ff_inst2(bidir_dq_7_oe_ff_inst2),
	.bidir_dq_0_oe_ff_inst3(bidir_dq_0_oe_ff_inst3),
	.bidir_dq_1_oe_ff_inst3(bidir_dq_1_oe_ff_inst3),
	.bidir_dq_2_oe_ff_inst3(bidir_dq_2_oe_ff_inst3),
	.bidir_dq_3_oe_ff_inst3(bidir_dq_3_oe_ff_inst3),
	.bidir_dq_4_oe_ff_inst3(bidir_dq_4_oe_ff_inst3),
	.bidir_dq_5_oe_ff_inst3(bidir_dq_5_oe_ff_inst3),
	.bidir_dq_6_oe_ff_inst3(bidir_dq_6_oe_ff_inst3),
	.bidir_dq_7_oe_ff_inst3(bidir_dq_7_oe_ff_inst3),
	.dqs_0_oe_ff_inst(dqs_0_oe_ff_inst),
	.dqs_0_oe_ff_inst1(dqs_0_oe_ff_inst1),
	.dqs_0_oe_ff_inst2(dqs_0_oe_ff_inst2),
	.dqs_0_oe_ff_inst3(dqs_0_oe_ff_inst3),
	.dqsn_0_oe_ff_inst(dqsn_0_oe_ff_inst),
	.dqsn_0_oe_ff_inst1(dqsn_0_oe_ff_inst1),
	.dqsn_0_oe_ff_inst2(dqsn_0_oe_ff_inst2),
	.dqsn_0_oe_ff_inst3(dqsn_0_oe_ff_inst3),
	.wd_lat_2(wd_lat_2),
	.wd_lat_1(wd_lat_1),
	.wd_lat_0(wd_lat_0),
	.wd_lat_3(wd_lat_3),
	.wd_lat_4(wd_lat_4),
	.afi_cs_n_1(afi_cs_n_1),
	.int_cke_r_0(int_cke_r_0),
	.afi_addr_0(afi_addr_0),
	.afi_addr_1(afi_addr_1),
	.afi_addr_2(afi_addr_2),
	.afi_addr_3(afi_addr_3),
	.afi_addr_4(afi_addr_4),
	.afi_addr_5(afi_addr_5),
	.afi_addr_6(afi_addr_6),
	.afi_addr_7(afi_addr_7),
	.afi_addr_8(afi_addr_8),
	.afi_addr_9(afi_addr_9),
	.afi_addr_10(afi_addr_10),
	.afi_addr_11(afi_addr_11),
	.afi_addr_12(afi_addr_12),
	.afi_addr_13(afi_addr_13),
	.afi_ba_0(afi_ba_0),
	.afi_ba_1(afi_ba_1),
	.afi_ba_2(afi_ba_2),
	.afi_ras_n_0(afi_ras_n_0),
	.afi_cas_n_0(afi_cas_n_0),
	.afi_we_n_0(afi_we_n_0),
	.afi_dm_4(afi_dm_4),
	.afi_dm_12(afi_dm_12),
	.afi_dm_0(afi_dm_0),
	.afi_dm_8(afi_dm_8),
	.afi_dm_5(afi_dm_5),
	.afi_dm_13(afi_dm_13),
	.afi_dm_1(afi_dm_1),
	.afi_dm_9(afi_dm_9),
	.afi_dm_6(afi_dm_6),
	.afi_dm_14(afi_dm_14),
	.afi_dm_2(afi_dm_2),
	.afi_dm_10(afi_dm_10),
	.afi_dm_7(afi_dm_7),
	.afi_dm_15(afi_dm_15),
	.afi_dm_3(afi_dm_3),
	.afi_dm_11(afi_dm_11),
	.int_wdata_valid(int_wdata_valid),
	.int_dqs_burst(int_dqs_burst),
	.int_dqs_burst_hr(int_dqs_burst_hr),
	.GND_port(GND_port),
	.global_reset_n(global_reset_n),
	.pll_ref_clk(pll_ref_clk),
	.soft_reset_n(soft_reset_n));

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy (
	q_b_0,
	q_b_64,
	q_b_1,
	q_b_65,
	q_b_2,
	q_b_66,
	q_b_3,
	q_b_67,
	q_b_4,
	q_b_68,
	q_b_5,
	q_b_69,
	q_b_6,
	q_b_70,
	q_b_7,
	q_b_71,
	q_b_16,
	q_b_80,
	q_b_17,
	q_b_81,
	q_b_18,
	q_b_82,
	q_b_19,
	q_b_83,
	q_b_20,
	q_b_84,
	q_b_21,
	q_b_85,
	q_b_22,
	q_b_86,
	q_b_23,
	q_b_87,
	q_b_32,
	q_b_96,
	q_b_33,
	q_b_97,
	q_b_34,
	q_b_98,
	q_b_35,
	q_b_99,
	q_b_36,
	q_b_100,
	q_b_37,
	q_b_101,
	q_b_38,
	q_b_102,
	q_b_39,
	q_b_103,
	q_b_48,
	q_b_112,
	q_b_49,
	q_b_113,
	q_b_50,
	q_b_114,
	q_b_51,
	q_b_115,
	q_b_52,
	q_b_116,
	q_b_53,
	q_b_117,
	q_b_54,
	q_b_118,
	q_b_55,
	q_b_119,
	q_b_8,
	q_b_72,
	q_b_9,
	q_b_73,
	q_b_10,
	q_b_74,
	q_b_11,
	q_b_75,
	q_b_12,
	q_b_76,
	q_b_13,
	q_b_77,
	q_b_14,
	q_b_78,
	q_b_15,
	q_b_79,
	q_b_24,
	q_b_88,
	q_b_25,
	q_b_89,
	q_b_26,
	q_b_90,
	q_b_27,
	q_b_91,
	q_b_28,
	q_b_92,
	q_b_29,
	q_b_93,
	q_b_30,
	q_b_94,
	q_b_31,
	q_b_95,
	q_b_40,
	q_b_104,
	q_b_41,
	q_b_105,
	q_b_42,
	q_b_106,
	q_b_43,
	q_b_107,
	q_b_44,
	q_b_108,
	q_b_45,
	q_b_109,
	q_b_46,
	q_b_110,
	q_b_47,
	q_b_111,
	q_b_56,
	q_b_120,
	q_b_57,
	q_b_121,
	q_b_58,
	q_b_122,
	q_b_59,
	q_b_123,
	q_b_60,
	q_b_124,
	q_b_61,
	q_b_125,
	q_b_62,
	q_b_126,
	q_b_63,
	q_b_127,
	clk_0,
	clk_1,
	dataout_0,
	dataout_01,
	dataout_02,
	dataout_03,
	dataout_04,
	dataout_05,
	dataout_06,
	dataout_07,
	dataout_08,
	dataout_09,
	dataout_010,
	dataout_011,
	dataout_012,
	dataout_013,
	dataout_014,
	dataout_015,
	dataout_016,
	dataout_017,
	dataout_018,
	dataout_019,
	dataout_020,
	dataout_021,
	dataout_022,
	dataout_023,
	dqs_delay_ctrl_0,
	dqs_delay_ctrl_1,
	dqs_delay_ctrl_2,
	dqs_delay_ctrl_3,
	dqs_delay_ctrl_4,
	dqs_delay_ctrl_5,
	wire_output_dq_0_output_ddio_out_inst_dataout,
	wire_output_dq_0_output_ddio_out_inst_dataout1,
	wire_output_dq_0_output_ddio_out_inst_dataout2,
	wire_output_dq_0_output_ddio_out_inst_dataout3,
	do_read_r,
	mem_clk_buf_in_0,
	mem_clk_n_buf_in_0,
	wire_bidir_dq_0_output_ddio_out_inst_dataout,
	wire_bidir_dq_1_output_ddio_out_inst_dataout,
	wire_bidir_dq_2_output_ddio_out_inst_dataout,
	wire_bidir_dq_3_output_ddio_out_inst_dataout,
	wire_bidir_dq_4_output_ddio_out_inst_dataout,
	wire_bidir_dq_5_output_ddio_out_inst_dataout,
	wire_bidir_dq_6_output_ddio_out_inst_dataout,
	wire_bidir_dq_7_output_ddio_out_inst_dataout,
	wire_bidir_dq_0_output_ddio_out_inst_dataout1,
	wire_bidir_dq_1_output_ddio_out_inst_dataout1,
	wire_bidir_dq_2_output_ddio_out_inst_dataout1,
	wire_bidir_dq_3_output_ddio_out_inst_dataout1,
	wire_bidir_dq_4_output_ddio_out_inst_dataout1,
	wire_bidir_dq_5_output_ddio_out_inst_dataout1,
	wire_bidir_dq_6_output_ddio_out_inst_dataout1,
	wire_bidir_dq_7_output_ddio_out_inst_dataout1,
	wire_bidir_dq_0_output_ddio_out_inst_dataout2,
	wire_bidir_dq_1_output_ddio_out_inst_dataout2,
	wire_bidir_dq_2_output_ddio_out_inst_dataout2,
	wire_bidir_dq_3_output_ddio_out_inst_dataout2,
	wire_bidir_dq_4_output_ddio_out_inst_dataout2,
	wire_bidir_dq_5_output_ddio_out_inst_dataout2,
	wire_bidir_dq_6_output_ddio_out_inst_dataout2,
	wire_bidir_dq_7_output_ddio_out_inst_dataout2,
	wire_bidir_dq_0_output_ddio_out_inst_dataout3,
	wire_bidir_dq_1_output_ddio_out_inst_dataout3,
	wire_bidir_dq_2_output_ddio_out_inst_dataout3,
	wire_bidir_dq_3_output_ddio_out_inst_dataout3,
	wire_bidir_dq_4_output_ddio_out_inst_dataout3,
	wire_bidir_dq_5_output_ddio_out_inst_dataout3,
	wire_bidir_dq_6_output_ddio_out_inst_dataout3,
	wire_bidir_dq_7_output_ddio_out_inst_dataout3,
	dqs_pseudo_diff_out_0,
	dqsn_pseudo_diff_out_0,
	dqs_pseudo_diff_out_1,
	dqsn_pseudo_diff_out_1,
	dqs_pseudo_diff_out_2,
	dqsn_pseudo_diff_out_2,
	dqs_pseudo_diff_out_3,
	dqsn_pseudo_diff_out_3,
	dq_datain_0,
	dq_datain_1,
	dq_datain_2,
	dq_datain_3,
	dq_datain_4,
	dq_datain_5,
	dq_datain_6,
	dq_datain_7,
	dq_datain_8,
	dq_datain_9,
	dq_datain_10,
	dq_datain_11,
	dq_datain_12,
	dq_datain_13,
	dq_datain_14,
	dq_datain_15,
	dq_datain_16,
	dq_datain_17,
	dq_datain_18,
	dq_datain_19,
	dq_datain_20,
	dq_datain_21,
	dq_datain_22,
	dq_datain_23,
	dq_datain_24,
	dq_datain_25,
	dq_datain_26,
	dq_datain_27,
	dq_datain_28,
	dq_datain_29,
	dq_datain_30,
	dq_datain_31,
	dqs_buffered_0,
	dqs_buffered_1,
	dqs_buffered_2,
	dqs_buffered_3,
	q_b_961,
	q_b_321,
	q_b_641,
	q_b_01,
	q_b_971,
	q_b_331,
	q_b_651,
	q_b_128,
	q_b_981,
	q_b_341,
	q_b_661,
	q_b_210,
	q_b_991,
	q_b_351,
	q_b_671,
	q_b_310,
	q_b_1001,
	q_b_361,
	q_b_681,
	q_b_410,
	q_b_1011,
	q_b_371,
	q_b_691,
	q_b_510,
	q_b_1021,
	q_b_381,
	q_b_701,
	q_b_610,
	q_b_1031,
	q_b_391,
	q_b_711,
	q_b_710,
	q_b_1041,
	q_b_401,
	q_b_721,
	q_b_810,
	q_b_1051,
	q_b_411,
	q_b_731,
	q_b_910,
	q_b_1061,
	q_b_421,
	q_b_741,
	q_b_1010,
	q_b_1071,
	q_b_431,
	q_b_751,
	q_b_1110,
	q_b_1081,
	q_b_441,
	q_b_761,
	q_b_129,
	q_b_1091,
	q_b_451,
	q_b_771,
	q_b_131,
	q_b_1101,
	q_b_461,
	q_b_781,
	q_b_141,
	q_b_1111,
	q_b_471,
	q_b_791,
	q_b_151,
	q_b_1121,
	q_b_481,
	q_b_801,
	q_b_161,
	q_b_1131,
	q_b_491,
	q_b_811,
	q_b_171,
	q_b_1141,
	q_b_501,
	q_b_821,
	q_b_181,
	q_b_1151,
	q_b_511,
	q_b_831,
	q_b_191,
	q_b_1161,
	q_b_521,
	q_b_841,
	q_b_201,
	q_b_1171,
	q_b_531,
	q_b_851,
	q_b_211,
	q_b_1181,
	q_b_541,
	q_b_861,
	q_b_221,
	q_b_1191,
	q_b_551,
	q_b_871,
	q_b_231,
	q_b_1201,
	q_b_561,
	q_b_881,
	q_b_241,
	q_b_1211,
	q_b_571,
	q_b_891,
	q_b_251,
	q_b_1221,
	q_b_581,
	q_b_901,
	q_b_261,
	q_b_1231,
	q_b_591,
	q_b_911,
	q_b_271,
	q_b_1241,
	q_b_601,
	q_b_921,
	q_b_281,
	q_b_1251,
	q_b_611,
	q_b_931,
	q_b_291,
	q_b_1261,
	q_b_621,
	q_b_941,
	q_b_301,
	q_b_1271,
	q_b_631,
	q_b_951,
	q_b_311,
	fb_clk,
	ctl_rdata_valid_0,
	reset_request_n,
	ctl_init_fail,
	ctl_init_success,
	reset_phy_clk_1x_n,
	rdwr_data_valid_r,
	doing_read,
	bidir_dq_0_oe_ff_inst,
	bidir_dq_1_oe_ff_inst,
	bidir_dq_2_oe_ff_inst,
	bidir_dq_3_oe_ff_inst,
	bidir_dq_4_oe_ff_inst,
	bidir_dq_5_oe_ff_inst,
	bidir_dq_6_oe_ff_inst,
	bidir_dq_7_oe_ff_inst,
	bidir_dq_0_oe_ff_inst1,
	bidir_dq_1_oe_ff_inst1,
	bidir_dq_2_oe_ff_inst1,
	bidir_dq_3_oe_ff_inst1,
	bidir_dq_4_oe_ff_inst1,
	bidir_dq_5_oe_ff_inst1,
	bidir_dq_6_oe_ff_inst1,
	bidir_dq_7_oe_ff_inst1,
	bidir_dq_0_oe_ff_inst2,
	bidir_dq_1_oe_ff_inst2,
	bidir_dq_2_oe_ff_inst2,
	bidir_dq_3_oe_ff_inst2,
	bidir_dq_4_oe_ff_inst2,
	bidir_dq_5_oe_ff_inst2,
	bidir_dq_6_oe_ff_inst2,
	bidir_dq_7_oe_ff_inst2,
	bidir_dq_0_oe_ff_inst3,
	bidir_dq_1_oe_ff_inst3,
	bidir_dq_2_oe_ff_inst3,
	bidir_dq_3_oe_ff_inst3,
	bidir_dq_4_oe_ff_inst3,
	bidir_dq_5_oe_ff_inst3,
	bidir_dq_6_oe_ff_inst3,
	bidir_dq_7_oe_ff_inst3,
	dqs_0_oe_ff_inst,
	dqs_0_oe_ff_inst1,
	dqs_0_oe_ff_inst2,
	dqs_0_oe_ff_inst3,
	dqsn_0_oe_ff_inst,
	dqsn_0_oe_ff_inst1,
	dqsn_0_oe_ff_inst2,
	dqsn_0_oe_ff_inst3,
	wd_lat_2,
	wd_lat_1,
	wd_lat_0,
	wd_lat_3,
	wd_lat_4,
	afi_cs_n_1,
	int_cke_r_0,
	afi_addr_0,
	afi_addr_1,
	afi_addr_2,
	afi_addr_3,
	afi_addr_4,
	afi_addr_5,
	afi_addr_6,
	afi_addr_7,
	afi_addr_8,
	afi_addr_9,
	afi_addr_10,
	afi_addr_11,
	afi_addr_12,
	afi_addr_13,
	afi_ba_0,
	afi_ba_1,
	afi_ba_2,
	afi_ras_n_0,
	afi_cas_n_0,
	afi_we_n_0,
	afi_dm_4,
	afi_dm_12,
	afi_dm_0,
	afi_dm_8,
	afi_dm_5,
	afi_dm_13,
	afi_dm_1,
	afi_dm_9,
	afi_dm_6,
	afi_dm_14,
	afi_dm_2,
	afi_dm_10,
	afi_dm_7,
	afi_dm_15,
	afi_dm_3,
	afi_dm_11,
	int_wdata_valid,
	int_dqs_burst,
	int_dqs_burst_hr,
	GND_port,
	global_reset_n,
	pll_ref_clk,
	soft_reset_n)/* synthesis synthesis_greybox=0 */;
output 	q_b_0;
output 	q_b_64;
output 	q_b_1;
output 	q_b_65;
output 	q_b_2;
output 	q_b_66;
output 	q_b_3;
output 	q_b_67;
output 	q_b_4;
output 	q_b_68;
output 	q_b_5;
output 	q_b_69;
output 	q_b_6;
output 	q_b_70;
output 	q_b_7;
output 	q_b_71;
output 	q_b_16;
output 	q_b_80;
output 	q_b_17;
output 	q_b_81;
output 	q_b_18;
output 	q_b_82;
output 	q_b_19;
output 	q_b_83;
output 	q_b_20;
output 	q_b_84;
output 	q_b_21;
output 	q_b_85;
output 	q_b_22;
output 	q_b_86;
output 	q_b_23;
output 	q_b_87;
output 	q_b_32;
output 	q_b_96;
output 	q_b_33;
output 	q_b_97;
output 	q_b_34;
output 	q_b_98;
output 	q_b_35;
output 	q_b_99;
output 	q_b_36;
output 	q_b_100;
output 	q_b_37;
output 	q_b_101;
output 	q_b_38;
output 	q_b_102;
output 	q_b_39;
output 	q_b_103;
output 	q_b_48;
output 	q_b_112;
output 	q_b_49;
output 	q_b_113;
output 	q_b_50;
output 	q_b_114;
output 	q_b_51;
output 	q_b_115;
output 	q_b_52;
output 	q_b_116;
output 	q_b_53;
output 	q_b_117;
output 	q_b_54;
output 	q_b_118;
output 	q_b_55;
output 	q_b_119;
output 	q_b_8;
output 	q_b_72;
output 	q_b_9;
output 	q_b_73;
output 	q_b_10;
output 	q_b_74;
output 	q_b_11;
output 	q_b_75;
output 	q_b_12;
output 	q_b_76;
output 	q_b_13;
output 	q_b_77;
output 	q_b_14;
output 	q_b_78;
output 	q_b_15;
output 	q_b_79;
output 	q_b_24;
output 	q_b_88;
output 	q_b_25;
output 	q_b_89;
output 	q_b_26;
output 	q_b_90;
output 	q_b_27;
output 	q_b_91;
output 	q_b_28;
output 	q_b_92;
output 	q_b_29;
output 	q_b_93;
output 	q_b_30;
output 	q_b_94;
output 	q_b_31;
output 	q_b_95;
output 	q_b_40;
output 	q_b_104;
output 	q_b_41;
output 	q_b_105;
output 	q_b_42;
output 	q_b_106;
output 	q_b_43;
output 	q_b_107;
output 	q_b_44;
output 	q_b_108;
output 	q_b_45;
output 	q_b_109;
output 	q_b_46;
output 	q_b_110;
output 	q_b_47;
output 	q_b_111;
output 	q_b_56;
output 	q_b_120;
output 	q_b_57;
output 	q_b_121;
output 	q_b_58;
output 	q_b_122;
output 	q_b_59;
output 	q_b_123;
output 	q_b_60;
output 	q_b_124;
output 	q_b_61;
output 	q_b_125;
output 	q_b_62;
output 	q_b_126;
output 	q_b_63;
output 	q_b_127;
output 	clk_0;
output 	clk_1;
output 	dataout_0;
output 	dataout_01;
output 	dataout_02;
output 	dataout_03;
output 	dataout_04;
output 	dataout_05;
output 	dataout_06;
output 	dataout_07;
output 	dataout_08;
output 	dataout_09;
output 	dataout_010;
output 	dataout_011;
output 	dataout_012;
output 	dataout_013;
output 	dataout_014;
output 	dataout_015;
output 	dataout_016;
output 	dataout_017;
output 	dataout_018;
output 	dataout_019;
output 	dataout_020;
output 	dataout_021;
output 	dataout_022;
output 	dataout_023;
output 	dqs_delay_ctrl_0;
output 	dqs_delay_ctrl_1;
output 	dqs_delay_ctrl_2;
output 	dqs_delay_ctrl_3;
output 	dqs_delay_ctrl_4;
output 	dqs_delay_ctrl_5;
output 	wire_output_dq_0_output_ddio_out_inst_dataout;
output 	wire_output_dq_0_output_ddio_out_inst_dataout1;
output 	wire_output_dq_0_output_ddio_out_inst_dataout2;
output 	wire_output_dq_0_output_ddio_out_inst_dataout3;
input 	do_read_r;
output 	mem_clk_buf_in_0;
output 	mem_clk_n_buf_in_0;
output 	wire_bidir_dq_0_output_ddio_out_inst_dataout;
output 	wire_bidir_dq_1_output_ddio_out_inst_dataout;
output 	wire_bidir_dq_2_output_ddio_out_inst_dataout;
output 	wire_bidir_dq_3_output_ddio_out_inst_dataout;
output 	wire_bidir_dq_4_output_ddio_out_inst_dataout;
output 	wire_bidir_dq_5_output_ddio_out_inst_dataout;
output 	wire_bidir_dq_6_output_ddio_out_inst_dataout;
output 	wire_bidir_dq_7_output_ddio_out_inst_dataout;
output 	wire_bidir_dq_0_output_ddio_out_inst_dataout1;
output 	wire_bidir_dq_1_output_ddio_out_inst_dataout1;
output 	wire_bidir_dq_2_output_ddio_out_inst_dataout1;
output 	wire_bidir_dq_3_output_ddio_out_inst_dataout1;
output 	wire_bidir_dq_4_output_ddio_out_inst_dataout1;
output 	wire_bidir_dq_5_output_ddio_out_inst_dataout1;
output 	wire_bidir_dq_6_output_ddio_out_inst_dataout1;
output 	wire_bidir_dq_7_output_ddio_out_inst_dataout1;
output 	wire_bidir_dq_0_output_ddio_out_inst_dataout2;
output 	wire_bidir_dq_1_output_ddio_out_inst_dataout2;
output 	wire_bidir_dq_2_output_ddio_out_inst_dataout2;
output 	wire_bidir_dq_3_output_ddio_out_inst_dataout2;
output 	wire_bidir_dq_4_output_ddio_out_inst_dataout2;
output 	wire_bidir_dq_5_output_ddio_out_inst_dataout2;
output 	wire_bidir_dq_6_output_ddio_out_inst_dataout2;
output 	wire_bidir_dq_7_output_ddio_out_inst_dataout2;
output 	wire_bidir_dq_0_output_ddio_out_inst_dataout3;
output 	wire_bidir_dq_1_output_ddio_out_inst_dataout3;
output 	wire_bidir_dq_2_output_ddio_out_inst_dataout3;
output 	wire_bidir_dq_3_output_ddio_out_inst_dataout3;
output 	wire_bidir_dq_4_output_ddio_out_inst_dataout3;
output 	wire_bidir_dq_5_output_ddio_out_inst_dataout3;
output 	wire_bidir_dq_6_output_ddio_out_inst_dataout3;
output 	wire_bidir_dq_7_output_ddio_out_inst_dataout3;
output 	dqs_pseudo_diff_out_0;
output 	dqsn_pseudo_diff_out_0;
output 	dqs_pseudo_diff_out_1;
output 	dqsn_pseudo_diff_out_1;
output 	dqs_pseudo_diff_out_2;
output 	dqsn_pseudo_diff_out_2;
output 	dqs_pseudo_diff_out_3;
output 	dqsn_pseudo_diff_out_3;
input 	dq_datain_0;
input 	dq_datain_1;
input 	dq_datain_2;
input 	dq_datain_3;
input 	dq_datain_4;
input 	dq_datain_5;
input 	dq_datain_6;
input 	dq_datain_7;
input 	dq_datain_8;
input 	dq_datain_9;
input 	dq_datain_10;
input 	dq_datain_11;
input 	dq_datain_12;
input 	dq_datain_13;
input 	dq_datain_14;
input 	dq_datain_15;
input 	dq_datain_16;
input 	dq_datain_17;
input 	dq_datain_18;
input 	dq_datain_19;
input 	dq_datain_20;
input 	dq_datain_21;
input 	dq_datain_22;
input 	dq_datain_23;
input 	dq_datain_24;
input 	dq_datain_25;
input 	dq_datain_26;
input 	dq_datain_27;
input 	dq_datain_28;
input 	dq_datain_29;
input 	dq_datain_30;
input 	dq_datain_31;
input 	dqs_buffered_0;
input 	dqs_buffered_1;
input 	dqs_buffered_2;
input 	dqs_buffered_3;
input 	q_b_961;
input 	q_b_321;
input 	q_b_641;
input 	q_b_01;
input 	q_b_971;
input 	q_b_331;
input 	q_b_651;
input 	q_b_128;
input 	q_b_981;
input 	q_b_341;
input 	q_b_661;
input 	q_b_210;
input 	q_b_991;
input 	q_b_351;
input 	q_b_671;
input 	q_b_310;
input 	q_b_1001;
input 	q_b_361;
input 	q_b_681;
input 	q_b_410;
input 	q_b_1011;
input 	q_b_371;
input 	q_b_691;
input 	q_b_510;
input 	q_b_1021;
input 	q_b_381;
input 	q_b_701;
input 	q_b_610;
input 	q_b_1031;
input 	q_b_391;
input 	q_b_711;
input 	q_b_710;
input 	q_b_1041;
input 	q_b_401;
input 	q_b_721;
input 	q_b_810;
input 	q_b_1051;
input 	q_b_411;
input 	q_b_731;
input 	q_b_910;
input 	q_b_1061;
input 	q_b_421;
input 	q_b_741;
input 	q_b_1010;
input 	q_b_1071;
input 	q_b_431;
input 	q_b_751;
input 	q_b_1110;
input 	q_b_1081;
input 	q_b_441;
input 	q_b_761;
input 	q_b_129;
input 	q_b_1091;
input 	q_b_451;
input 	q_b_771;
input 	q_b_131;
input 	q_b_1101;
input 	q_b_461;
input 	q_b_781;
input 	q_b_141;
input 	q_b_1111;
input 	q_b_471;
input 	q_b_791;
input 	q_b_151;
input 	q_b_1121;
input 	q_b_481;
input 	q_b_801;
input 	q_b_161;
input 	q_b_1131;
input 	q_b_491;
input 	q_b_811;
input 	q_b_171;
input 	q_b_1141;
input 	q_b_501;
input 	q_b_821;
input 	q_b_181;
input 	q_b_1151;
input 	q_b_511;
input 	q_b_831;
input 	q_b_191;
input 	q_b_1161;
input 	q_b_521;
input 	q_b_841;
input 	q_b_201;
input 	q_b_1171;
input 	q_b_531;
input 	q_b_851;
input 	q_b_211;
input 	q_b_1181;
input 	q_b_541;
input 	q_b_861;
input 	q_b_221;
input 	q_b_1191;
input 	q_b_551;
input 	q_b_871;
input 	q_b_231;
input 	q_b_1201;
input 	q_b_561;
input 	q_b_881;
input 	q_b_241;
input 	q_b_1211;
input 	q_b_571;
input 	q_b_891;
input 	q_b_251;
input 	q_b_1221;
input 	q_b_581;
input 	q_b_901;
input 	q_b_261;
input 	q_b_1231;
input 	q_b_591;
input 	q_b_911;
input 	q_b_271;
input 	q_b_1241;
input 	q_b_601;
input 	q_b_921;
input 	q_b_281;
input 	q_b_1251;
input 	q_b_611;
input 	q_b_931;
input 	q_b_291;
input 	q_b_1261;
input 	q_b_621;
input 	q_b_941;
input 	q_b_301;
input 	q_b_1271;
input 	q_b_631;
input 	q_b_951;
input 	q_b_311;
input 	fb_clk;
output 	ctl_rdata_valid_0;
output 	reset_request_n;
output 	ctl_init_fail;
output 	ctl_init_success;
output 	reset_phy_clk_1x_n;
input 	rdwr_data_valid_r;
input 	doing_read;
output 	bidir_dq_0_oe_ff_inst;
output 	bidir_dq_1_oe_ff_inst;
output 	bidir_dq_2_oe_ff_inst;
output 	bidir_dq_3_oe_ff_inst;
output 	bidir_dq_4_oe_ff_inst;
output 	bidir_dq_5_oe_ff_inst;
output 	bidir_dq_6_oe_ff_inst;
output 	bidir_dq_7_oe_ff_inst;
output 	bidir_dq_0_oe_ff_inst1;
output 	bidir_dq_1_oe_ff_inst1;
output 	bidir_dq_2_oe_ff_inst1;
output 	bidir_dq_3_oe_ff_inst1;
output 	bidir_dq_4_oe_ff_inst1;
output 	bidir_dq_5_oe_ff_inst1;
output 	bidir_dq_6_oe_ff_inst1;
output 	bidir_dq_7_oe_ff_inst1;
output 	bidir_dq_0_oe_ff_inst2;
output 	bidir_dq_1_oe_ff_inst2;
output 	bidir_dq_2_oe_ff_inst2;
output 	bidir_dq_3_oe_ff_inst2;
output 	bidir_dq_4_oe_ff_inst2;
output 	bidir_dq_5_oe_ff_inst2;
output 	bidir_dq_6_oe_ff_inst2;
output 	bidir_dq_7_oe_ff_inst2;
output 	bidir_dq_0_oe_ff_inst3;
output 	bidir_dq_1_oe_ff_inst3;
output 	bidir_dq_2_oe_ff_inst3;
output 	bidir_dq_3_oe_ff_inst3;
output 	bidir_dq_4_oe_ff_inst3;
output 	bidir_dq_5_oe_ff_inst3;
output 	bidir_dq_6_oe_ff_inst3;
output 	bidir_dq_7_oe_ff_inst3;
output 	dqs_0_oe_ff_inst;
output 	dqs_0_oe_ff_inst1;
output 	dqs_0_oe_ff_inst2;
output 	dqs_0_oe_ff_inst3;
output 	dqsn_0_oe_ff_inst;
output 	dqsn_0_oe_ff_inst1;
output 	dqsn_0_oe_ff_inst2;
output 	dqsn_0_oe_ff_inst3;
output 	wd_lat_2;
output 	wd_lat_1;
output 	wd_lat_0;
output 	wd_lat_3;
output 	wd_lat_4;
input 	afi_cs_n_1;
input 	int_cke_r_0;
input 	afi_addr_0;
input 	afi_addr_1;
input 	afi_addr_2;
input 	afi_addr_3;
input 	afi_addr_4;
input 	afi_addr_5;
input 	afi_addr_6;
input 	afi_addr_7;
input 	afi_addr_8;
input 	afi_addr_9;
input 	afi_addr_10;
input 	afi_addr_11;
input 	afi_addr_12;
input 	afi_addr_13;
input 	afi_ba_0;
input 	afi_ba_1;
input 	afi_ba_2;
input 	afi_ras_n_0;
input 	afi_cas_n_0;
input 	afi_we_n_0;
input 	afi_dm_4;
input 	afi_dm_12;
input 	afi_dm_0;
input 	afi_dm_8;
input 	afi_dm_5;
input 	afi_dm_13;
input 	afi_dm_1;
input 	afi_dm_9;
input 	afi_dm_6;
input 	afi_dm_14;
input 	afi_dm_2;
input 	afi_dm_10;
input 	afi_dm_7;
input 	afi_dm_15;
input 	afi_dm_3;
input 	afi_dm_11;
input 	int_wdata_valid;
input 	int_dqs_burst;
input 	int_dqs_burst_hr;
input 	GND_port;
input 	global_reset_n;
input 	pll_ref_clk;
input 	soft_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \clk|half_rate.pll|altpll_component|auto_generated|clk[3] ;
wire \clk|half_rate.pll|altpll_component|auto_generated|clk[4] ;
wire \clk|half_rate.pll|altpll_component|auto_generated|clk[5] ;
wire \half_rate_wdp_gen.wdp|wdp_dm_l_2x[0]~q ;
wire \half_rate_wdp_gen.wdp|wdp_dm_h_2x[0]~q ;
wire \half_rate_wdp_gen.wdp|wdp_dm_l_2x[1]~q ;
wire \half_rate_wdp_gen.wdp|wdp_dm_h_2x[1]~q ;
wire \half_rate_wdp_gen.wdp|wdp_dm_l_2x[2]~q ;
wire \half_rate_wdp_gen.wdp|wdp_dm_h_2x[2]~q ;
wire \half_rate_wdp_gen.wdp|wdp_dm_l_2x[3]~q ;
wire \half_rate_wdp_gen.wdp|wdp_dm_h_2x[3]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_l_2x[0]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_h_2x[0]~q ;
wire \half_rate_wdp_gen.wdp|dq_oe_2x[0]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_l_2x[1]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_h_2x[1]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_l_2x[2]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_h_2x[2]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_l_2x[3]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_h_2x[3]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_l_2x[4]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_h_2x[4]~q ;
wire \half_rate_wdp_gen.wdp|dq_oe_2x[1]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_l_2x[5]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_h_2x[5]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_l_2x[6]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_h_2x[6]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_l_2x[7]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_h_2x[7]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_l_2x[8]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_h_2x[8]~q ;
wire \half_rate_wdp_gen.wdp|dq_oe_2x[2]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_l_2x[9]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_h_2x[9]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_l_2x[10]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_h_2x[10]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_l_2x[11]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_h_2x[11]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_l_2x[12]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_h_2x[12]~q ;
wire \half_rate_wdp_gen.wdp|dq_oe_2x[3]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_l_2x[13]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_h_2x[13]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_l_2x[14]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_h_2x[14]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_l_2x[15]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_h_2x[15]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_l_2x[16]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_h_2x[16]~q ;
wire \half_rate_wdp_gen.wdp|dq_oe_2x[4]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_l_2x[17]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_h_2x[17]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_l_2x[18]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_h_2x[18]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_l_2x[19]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_h_2x[19]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_l_2x[20]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_h_2x[20]~q ;
wire \half_rate_wdp_gen.wdp|dq_oe_2x[5]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_l_2x[21]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_h_2x[21]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_l_2x[22]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_h_2x[22]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_l_2x[23]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_h_2x[23]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_l_2x[24]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_h_2x[24]~q ;
wire \half_rate_wdp_gen.wdp|dq_oe_2x[6]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_l_2x[25]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_h_2x[25]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_l_2x[26]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_h_2x[26]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_l_2x[27]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_h_2x[27]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_l_2x[28]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_h_2x[28]~q ;
wire \half_rate_wdp_gen.wdp|dq_oe_2x[7]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_l_2x[29]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_h_2x[29]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_l_2x[30]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_h_2x[30]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_l_2x[31]~q ;
wire \half_rate_wdp_gen.wdp|wdp_wdata_h_2x[31]~q ;
wire \seq_wrapper|seq_inst|seq_ac_cke[1]~q ;
wire \seq_wrapper|seq_inst|seq_ac_addr[0]~q ;
wire \seq_wrapper|seq_inst|seq_ac_addr[14]~q ;
wire \seq_wrapper|seq_inst|seq_ac_addr[1]~q ;
wire \seq_wrapper|seq_inst|seq_ac_addr[15]~q ;
wire \seq_wrapper|seq_inst|seq_ac_addr[16]~q ;
wire \seq_wrapper|seq_inst|seq_ac_addr[17]~q ;
wire \seq_wrapper|seq_inst|seq_ac_addr[18]~q ;
wire \seq_wrapper|seq_inst|seq_ac_addr[5]~q ;
wire \seq_wrapper|seq_inst|seq_ac_addr[19]~q ;
wire \seq_wrapper|seq_inst|seq_ac_addr[8]~q ;
wire \seq_wrapper|seq_inst|seq_ac_addr[22]~q ;
wire \seq_wrapper|seq_inst|seq_ac_addr[10]~q ;
wire \seq_wrapper|seq_inst|seq_ac_addr[24]~q ;
wire \seq_wrapper|seq_inst|seq_ac_addr[12]~q ;
wire \seq_wrapper|seq_inst|seq_ac_addr[26]~q ;
wire \seq_wrapper|seq_inst|seq_ac_ba[0]~q ;
wire \seq_wrapper|seq_inst|seq_ac_ba[3]~q ;
wire \seq_wrapper|seq_inst|seq_ac_ba[1]~q ;
wire \seq_wrapper|seq_inst|seq_ac_ba[4]~q ;
wire \seq_wrapper|seq_inst|seq_ac_rst_n[0]~q ;
wire \clk|mimic_data_2x ;
wire \dpio|dio_rdata_h_2x[0]~q ;
wire \poa|rd_addr_2x[0]~q ;
wire \rdv_pipe|rd_addr[0]~q ;
wire \dpio|dio_rdata_h_2x[1]~q ;
wire \dpio|dio_rdata_h_2x[2]~q ;
wire \dpio|dio_rdata_h_2x[3]~q ;
wire \dpio|dio_rdata_h_2x[4]~q ;
wire \dpio|dio_rdata_h_2x[5]~q ;
wire \dpio|dio_rdata_h_2x[6]~q ;
wire \dpio|dio_rdata_h_2x[7]~q ;
wire \dpio|dio_rdata_h_2x[8]~q ;
wire \dpio|dio_rdata_h_2x[9]~q ;
wire \dpio|dio_rdata_h_2x[10]~q ;
wire \dpio|dio_rdata_h_2x[11]~q ;
wire \dpio|dio_rdata_h_2x[12]~q ;
wire \dpio|dio_rdata_h_2x[13]~q ;
wire \dpio|dio_rdata_h_2x[14]~q ;
wire \dpio|dio_rdata_h_2x[15]~q ;
wire \dpio|dio_rdata_h_2x[16]~q ;
wire \dpio|dio_rdata_h_2x[17]~q ;
wire \dpio|dio_rdata_h_2x[18]~q ;
wire \dpio|dio_rdata_h_2x[19]~q ;
wire \dpio|dio_rdata_h_2x[20]~q ;
wire \dpio|dio_rdata_h_2x[21]~q ;
wire \dpio|dio_rdata_h_2x[22]~q ;
wire \dpio|dio_rdata_h_2x[23]~q ;
wire \dpio|dio_rdata_h_2x[24]~q ;
wire \dpio|dio_rdata_h_2x[25]~q ;
wire \dpio|dio_rdata_h_2x[26]~q ;
wire \dpio|dio_rdata_h_2x[27]~q ;
wire \dpio|dio_rdata_h_2x[28]~q ;
wire \dpio|dio_rdata_h_2x[29]~q ;
wire \dpio|dio_rdata_h_2x[30]~q ;
wire \dpio|dio_rdata_h_2x[31]~q ;
wire \dpio|dio_rdata_l_2x[0]~q ;
wire \dpio|dio_rdata_l_2x[1]~q ;
wire \dpio|dio_rdata_l_2x[2]~q ;
wire \dpio|dio_rdata_l_2x[3]~q ;
wire \dpio|dio_rdata_l_2x[4]~q ;
wire \dpio|dio_rdata_l_2x[5]~q ;
wire \dpio|dio_rdata_l_2x[6]~q ;
wire \dpio|dio_rdata_l_2x[7]~q ;
wire \dpio|dio_rdata_l_2x[8]~q ;
wire \dpio|dio_rdata_l_2x[9]~q ;
wire \dpio|dio_rdata_l_2x[10]~q ;
wire \dpio|dio_rdata_l_2x[11]~q ;
wire \dpio|dio_rdata_l_2x[12]~q ;
wire \dpio|dio_rdata_l_2x[13]~q ;
wire \dpio|dio_rdata_l_2x[14]~q ;
wire \dpio|dio_rdata_l_2x[15]~q ;
wire \dpio|dio_rdata_l_2x[16]~q ;
wire \dpio|dio_rdata_l_2x[17]~q ;
wire \dpio|dio_rdata_l_2x[18]~q ;
wire \dpio|dio_rdata_l_2x[19]~q ;
wire \dpio|dio_rdata_l_2x[20]~q ;
wire \dpio|dio_rdata_l_2x[21]~q ;
wire \dpio|dio_rdata_l_2x[22]~q ;
wire \dpio|dio_rdata_l_2x[23]~q ;
wire \dpio|dio_rdata_l_2x[24]~q ;
wire \dpio|dio_rdata_l_2x[25]~q ;
wire \dpio|dio_rdata_l_2x[26]~q ;
wire \dpio|dio_rdata_l_2x[27]~q ;
wire \dpio|dio_rdata_l_2x[28]~q ;
wire \dpio|dio_rdata_l_2x[29]~q ;
wire \dpio|dio_rdata_l_2x[30]~q ;
wire \dpio|dio_rdata_l_2x[31]~q ;
wire \clk|reset_rdp_phy_clk_pipe|ams_pipe[1]~q ;
wire \clk|ac_clk_pipe_2x|ams_pipe[1]~q ;
wire \seq_wrapper|seq_inst|ctrl|ctl_init_fail~q ;
wire \seq_wrapper|seq_inst|ctrl|ctl_init_success~q ;
wire \clk|resync_clk_2x_pipe|ams_pipe[1]~q ;
wire \seq_wrapper|seq_inst|seq_rdv_doing_rd[7]~q ;
wire \rdv_pipe|merged_doing_rd~0_combout ;
wire \seq_wrapper|seq_inst|seq_rdp_reset_req_n~q ;
wire \seq_wrapper|seq_inst|seq_ac_add_1t_ac_lat_internal~q ;
wire \seq_wrapper|seq_inst|seq_rdata_valid_lat_dec~q ;
wire \seq_wrapper|seq_inst|seq_rdv_doing_rd[4]~q ;
wire \seq_wrapper|seq_inst|seq_pll_inc_dec_n~q ;
wire \seq_wrapper|seq_inst|seq_pll_start_reconfig~q ;
wire \clk|write_clk_pipe|ams_pipe[3]~q ;
wire \half_rate_wdp_gen.wdp|dqs_burst_2x_r3[0]~q ;
wire \half_rate_wdp_gen.wdp|dqs_burst_2x_r3[1]~q ;
wire \half_rate_wdp_gen.wdp|dqs_burst_2x_r3[2]~q ;
wire \half_rate_wdp_gen.wdp|dqs_burst_2x_r3[3]~q ;
wire \seq_wrapper|seq_inst|seq_pll_select[2]~q ;
wire \seq_wrapper|seq_inst|seq_pll_select[1]~q ;
wire \seq_wrapper|seq_inst|seq_mem_clk_disable~q ;
wire \clk|mem_clk_pipe|ams_pipe[3]~q ;
wire \rdv_pipe|seq_rdata_valid[0]~q ;
wire \rdv_pipe|seq_rdata_valid[1]~q ;
wire \seq_wrapper|seq_inst|seq_ac_cs_n[0]~q ;
wire \seq_wrapper|seq_inst|admin|seq_ac_sel~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdp_ovride~q ;
wire \seq_wrapper|seq_inst|seq_wdp_ovride~0_combout ;
wire \poa|postamble_en_pos_2x[0]~q ;
wire \poa|postamble_en_pos_2x[1]~q ;
wire \poa|postamble_en_pos_2x[2]~q ;
wire \poa|postamble_en_pos_2x[3]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[120]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[56]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[88]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[24]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[121]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[57]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[89]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[25]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[122]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[58]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[90]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[26]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[123]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[59]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[91]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[27]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[124]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[60]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[92]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[28]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[125]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[61]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[93]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[29]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[126]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[62]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[94]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[30]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[127]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[63]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[95]~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdata[31]~q ;
wire \seq_wrapper|seq_inst|seq_poa_protection_override_1x~q ;
wire \seq_wrapper|seq_inst|seq_poa_lat_dec_1x[0]~q ;
wire \merged_doing_rd[4]~combout ;
wire \mmc|mimic_done_out~q ;
wire \clk|measure_clk_pipe|ams_pipe[1]~q ;
wire \clk|phs_shft_busy_siii~q ;
wire \seq_wrapper|seq_inst|dgrb|seq_mmc_start~q ;
wire \mmc|mimic_value_captured~q ;
wire \seq_wrapper|seq_inst|dgwb|dgwb_wdp_ovride~_wirecell_combout ;
wire \seq_wrapper|seq_inst|seq_ac_cas_n[0]~_wirecell_combout ;
wire \seq_wrapper|seq_inst|seq_ac_cas_n[1]~_wirecell_combout ;
wire \seq_wrapper|seq_inst|seq_ac_cs_n[1]~_wirecell_combout ;
wire \seq_wrapper|seq_inst|seq_ac_ras_n[0]~_wirecell_combout ;
wire \seq_wrapper|seq_inst|seq_ac_ras_n[1]~_wirecell_combout ;
wire \seq_wrapper|seq_inst|seq_ac_we_n[0]~_wirecell_combout ;
wire \seq_wrapper|seq_inst|seq_ac_we_n[1]~_wirecell_combout ;


ddr3_int_ddr3_int_phy_alt_mem_phy_rdata_valid rdv_pipe(
	.clk_0(clk_0),
	.do_read_r(do_read_r),
	.ctl_rdata_valid_0(ctl_rdata_valid_0),
	.ctl_init_success(ctl_init_success),
	.rd_addr_0(\rdv_pipe|rd_addr[0]~q ),
	.reset_phy_clk_1x_n(\clk|reset_rdp_phy_clk_pipe|ams_pipe[1]~q ),
	.rdwr_data_valid_r(rdwr_data_valid_r),
	.seq_rdv_doing_rd_7(\seq_wrapper|seq_inst|seq_rdv_doing_rd[7]~q ),
	.doing_read(doing_read),
	.merged_doing_rd(\rdv_pipe|merged_doing_rd~0_combout ),
	.seq_rdata_valid_lat_dec(\seq_wrapper|seq_inst|seq_rdata_valid_lat_dec~q ),
	.seq_rdv_doing_rd_4(\seq_wrapper|seq_inst|seq_rdv_doing_rd[4]~q ),
	.seq_rdata_valid_0(\rdv_pipe|seq_rdata_valid[0]~q ),
	.seq_rdata_valid_1(\rdv_pipe|seq_rdata_valid[1]~q ));

ddr3_int_ddr3_int_phy_alt_mem_phy_clk_reset clk(
	.clk_0(clk_0),
	.clk_1(clk_1),
	.clk_3(\clk|half_rate.pll|altpll_component|auto_generated|clk[3] ),
	.clk_4(\clk|half_rate.pll|altpll_component|auto_generated|clk[4] ),
	.clk_5(\clk|half_rate.pll|altpll_component|auto_generated|clk[5] ),
	.dqs_delay_ctrl({dqs_delay_ctrl_5,dqs_delay_ctrl_4,dqs_delay_ctrl_3,dqs_delay_ctrl_2,dqs_delay_ctrl_1,dqs_delay_ctrl_0}),
	.mem_clk_buf_in_0(mem_clk_buf_in_0),
	.mem_clk_n_buf_in_0(mem_clk_n_buf_in_0),
	.mimic_data_2x(\clk|mimic_data_2x ),
	.fb_clk(fb_clk),
	.reset_request_n(reset_request_n),
	.reset_phy_clk_1x_n1(reset_phy_clk_1x_n),
	.ams_pipe_1(\clk|reset_rdp_phy_clk_pipe|ams_pipe[1]~q ),
	.ams_pipe_11(\clk|ac_clk_pipe_2x|ams_pipe[1]~q ),
	.ams_pipe_12(\clk|resync_clk_2x_pipe|ams_pipe[1]~q ),
	.seq_rdp_reset_req_n(\seq_wrapper|seq_inst|seq_rdp_reset_req_n~q ),
	.seq_pll_inc_dec_n(\seq_wrapper|seq_inst|seq_pll_inc_dec_n~q ),
	.seq_pll_start_reconfig(\seq_wrapper|seq_inst|seq_pll_start_reconfig~q ),
	.ams_pipe_3(\clk|write_clk_pipe|ams_pipe[3]~q ),
	.seq_pll_select({\seq_wrapper|seq_inst|seq_pll_select[2]~q ,\seq_wrapper|seq_inst|seq_pll_select[1]~q ,\seq_wrapper|seq_inst|seq_pll_select[2]~q }),
	.seq_mem_clk_disable(\seq_wrapper|seq_inst|seq_mem_clk_disable~q ),
	.ams_pipe_31(\clk|mem_clk_pipe|ams_pipe[3]~q ),
	.ams_pipe_13(\clk|measure_clk_pipe|ams_pipe[1]~q ),
	.phs_shft_busy_siii1(\clk|phs_shft_busy_siii~q ),
	.global_reset_n(global_reset_n),
	.pll_ref_clk(pll_ref_clk),
	.soft_reset_n(soft_reset_n));

ddr3_int_ddr3_int_phy_alt_mem_phy_mimic mmc(
	.measure_clk(\clk|half_rate.pll|altpll_component|auto_generated|clk[5] ),
	.mimic_data_in(\clk|mimic_data_2x ),
	.mimic_done_out1(\mmc|mimic_done_out~q ),
	.reset_measure_clk_n(\clk|measure_clk_pipe|ams_pipe[1]~q ),
	.seq_mmc_start(\seq_wrapper|seq_inst|dgrb|seq_mmc_start~q ),
	.mimic_value_captured1(\mmc|mimic_value_captured~q ));

ddr3_int_ddr3_int_phy_alt_mem_phy_postamble poa(
	.clk_0(clk_0),
	.clk_4(\clk|half_rate.pll|altpll_component|auto_generated|clk[4] ),
	.rd_addr_2x_0(\poa|rd_addr_2x[0]~q ),
	.reset_phy_clk_1x_n(\clk|reset_rdp_phy_clk_pipe|ams_pipe[1]~q ),
	.reset_poa_clk_2x_n(\clk|resync_clk_2x_pipe|ams_pipe[1]~q ),
	.seq_rdv_doing_rd_7(\seq_wrapper|seq_inst|seq_rdv_doing_rd[7]~q ),
	.merged_doing_rd(\rdv_pipe|merged_doing_rd~0_combout ),
	.seq_rdv_doing_rd_4(\seq_wrapper|seq_inst|seq_rdv_doing_rd[4]~q ),
	.postamble_en_pos_2x_0(\poa|postamble_en_pos_2x[0]~q ),
	.postamble_en_pos_2x_1(\poa|postamble_en_pos_2x[1]~q ),
	.postamble_en_pos_2x_2(\poa|postamble_en_pos_2x[2]~q ),
	.postamble_en_pos_2x_3(\poa|postamble_en_pos_2x[3]~q ),
	.seq_poa_protection_override_1x(\seq_wrapper|seq_inst|seq_poa_protection_override_1x~q ),
	.seq_poa_lat_dec_1x(\seq_wrapper|seq_inst|seq_poa_lat_dec_1x[0]~q ),
	.ctl_doing_rd_beat2_1x(\merged_doing_rd[4]~combout ));

ddr3_int_ddr3_int_phy_alt_mem_phy_seq_wrapper seq_wrapper(
	.q_b_0(q_b_0),
	.q_b_64(q_b_64),
	.q_b_1(q_b_1),
	.q_b_65(q_b_65),
	.q_b_2(q_b_2),
	.q_b_66(q_b_66),
	.q_b_3(q_b_3),
	.q_b_67(q_b_67),
	.q_b_4(q_b_4),
	.q_b_68(q_b_68),
	.q_b_5(q_b_5),
	.q_b_69(q_b_69),
	.q_b_6(q_b_6),
	.q_b_70(q_b_70),
	.q_b_7(q_b_7),
	.q_b_71(q_b_71),
	.q_b_16(q_b_16),
	.q_b_80(q_b_80),
	.q_b_17(q_b_17),
	.q_b_81(q_b_81),
	.q_b_18(q_b_18),
	.q_b_82(q_b_82),
	.q_b_19(q_b_19),
	.q_b_83(q_b_83),
	.q_b_20(q_b_20),
	.q_b_84(q_b_84),
	.q_b_21(q_b_21),
	.q_b_85(q_b_85),
	.q_b_22(q_b_22),
	.q_b_86(q_b_86),
	.q_b_23(q_b_23),
	.q_b_87(q_b_87),
	.q_b_32(q_b_32),
	.q_b_96(q_b_96),
	.q_b_33(q_b_33),
	.q_b_97(q_b_97),
	.q_b_34(q_b_34),
	.q_b_98(q_b_98),
	.q_b_35(q_b_35),
	.q_b_99(q_b_99),
	.q_b_36(q_b_36),
	.q_b_100(q_b_100),
	.q_b_37(q_b_37),
	.q_b_101(q_b_101),
	.q_b_38(q_b_38),
	.q_b_102(q_b_102),
	.q_b_39(q_b_39),
	.q_b_103(q_b_103),
	.q_b_48(q_b_48),
	.q_b_112(q_b_112),
	.q_b_49(q_b_49),
	.q_b_113(q_b_113),
	.q_b_50(q_b_50),
	.q_b_114(q_b_114),
	.q_b_51(q_b_51),
	.q_b_115(q_b_115),
	.q_b_52(q_b_52),
	.q_b_116(q_b_116),
	.q_b_53(q_b_53),
	.q_b_117(q_b_117),
	.q_b_54(q_b_54),
	.q_b_118(q_b_118),
	.q_b_55(q_b_55),
	.q_b_119(q_b_119),
	.q_b_8(q_b_8),
	.q_b_72(q_b_72),
	.q_b_9(q_b_9),
	.q_b_73(q_b_73),
	.q_b_10(q_b_10),
	.q_b_74(q_b_74),
	.q_b_11(q_b_11),
	.q_b_75(q_b_75),
	.q_b_12(q_b_12),
	.q_b_76(q_b_76),
	.q_b_13(q_b_13),
	.q_b_77(q_b_77),
	.q_b_14(q_b_14),
	.q_b_78(q_b_78),
	.q_b_15(q_b_15),
	.q_b_79(q_b_79),
	.q_b_24(q_b_24),
	.q_b_88(q_b_88),
	.q_b_25(q_b_25),
	.q_b_89(q_b_89),
	.q_b_26(q_b_26),
	.q_b_90(q_b_90),
	.q_b_27(q_b_27),
	.q_b_91(q_b_91),
	.q_b_28(q_b_28),
	.q_b_92(q_b_92),
	.q_b_29(q_b_29),
	.q_b_93(q_b_93),
	.q_b_30(q_b_30),
	.q_b_94(q_b_94),
	.q_b_31(q_b_31),
	.q_b_95(q_b_95),
	.q_b_40(q_b_40),
	.q_b_104(q_b_104),
	.q_b_41(q_b_41),
	.q_b_105(q_b_105),
	.q_b_42(q_b_42),
	.q_b_106(q_b_106),
	.q_b_43(q_b_43),
	.q_b_107(q_b_107),
	.q_b_44(q_b_44),
	.q_b_108(q_b_108),
	.q_b_45(q_b_45),
	.q_b_109(q_b_109),
	.q_b_46(q_b_46),
	.q_b_110(q_b_110),
	.q_b_47(q_b_47),
	.q_b_111(q_b_111),
	.q_b_56(q_b_56),
	.q_b_120(q_b_120),
	.q_b_57(q_b_57),
	.q_b_121(q_b_121),
	.q_b_58(q_b_58),
	.q_b_122(q_b_122),
	.q_b_59(q_b_59),
	.q_b_123(q_b_123),
	.q_b_60(q_b_60),
	.q_b_124(q_b_124),
	.q_b_61(q_b_61),
	.q_b_125(q_b_125),
	.q_b_62(q_b_62),
	.q_b_126(q_b_126),
	.q_b_63(q_b_63),
	.q_b_127(q_b_127),
	.clk_0(clk_0),
	.seq_ac_cke_1(\seq_wrapper|seq_inst|seq_ac_cke[1]~q ),
	.seq_ac_addr_0(\seq_wrapper|seq_inst|seq_ac_addr[0]~q ),
	.seq_ac_addr_14(\seq_wrapper|seq_inst|seq_ac_addr[14]~q ),
	.seq_ac_addr_1(\seq_wrapper|seq_inst|seq_ac_addr[1]~q ),
	.seq_ac_addr_15(\seq_wrapper|seq_inst|seq_ac_addr[15]~q ),
	.seq_ac_addr_16(\seq_wrapper|seq_inst|seq_ac_addr[16]~q ),
	.seq_ac_addr_17(\seq_wrapper|seq_inst|seq_ac_addr[17]~q ),
	.seq_ac_addr_18(\seq_wrapper|seq_inst|seq_ac_addr[18]~q ),
	.seq_ac_addr_5(\seq_wrapper|seq_inst|seq_ac_addr[5]~q ),
	.seq_ac_addr_19(\seq_wrapper|seq_inst|seq_ac_addr[19]~q ),
	.seq_ac_addr_8(\seq_wrapper|seq_inst|seq_ac_addr[8]~q ),
	.seq_ac_addr_22(\seq_wrapper|seq_inst|seq_ac_addr[22]~q ),
	.seq_ac_addr_10(\seq_wrapper|seq_inst|seq_ac_addr[10]~q ),
	.seq_ac_addr_24(\seq_wrapper|seq_inst|seq_ac_addr[24]~q ),
	.seq_ac_addr_12(\seq_wrapper|seq_inst|seq_ac_addr[12]~q ),
	.seq_ac_addr_26(\seq_wrapper|seq_inst|seq_ac_addr[26]~q ),
	.seq_ac_ba_0(\seq_wrapper|seq_inst|seq_ac_ba[0]~q ),
	.seq_ac_ba_3(\seq_wrapper|seq_inst|seq_ac_ba[3]~q ),
	.seq_ac_ba_1(\seq_wrapper|seq_inst|seq_ac_ba[1]~q ),
	.seq_ac_ba_4(\seq_wrapper|seq_inst|seq_ac_ba[4]~q ),
	.seq_ac_rst_n_0(\seq_wrapper|seq_inst|seq_ac_rst_n[0]~q ),
	.ctl_init_fail(ctl_init_fail),
	.ctl_init_success(ctl_init_success),
	.reset_phy_clk_1x_n(reset_phy_clk_1x_n),
	.ctl_init_fail1(\seq_wrapper|seq_inst|ctrl|ctl_init_fail~q ),
	.ctl_init_success1(\seq_wrapper|seq_inst|ctrl|ctl_init_success~q ),
	.seq_rdv_doing_rd_7(\seq_wrapper|seq_inst|seq_rdv_doing_rd[7]~q ),
	.seq_rdp_reset_req_n(\seq_wrapper|seq_inst|seq_rdp_reset_req_n~q ),
	.seq_ac_add_1t_ac_lat_internal(\seq_wrapper|seq_inst|seq_ac_add_1t_ac_lat_internal~q ),
	.wd_lat_2(wd_lat_2),
	.wd_lat_1(wd_lat_1),
	.wd_lat_0(wd_lat_0),
	.wd_lat_3(wd_lat_3),
	.wd_lat_4(wd_lat_4),
	.seq_rdata_valid_lat_dec(\seq_wrapper|seq_inst|seq_rdata_valid_lat_dec~q ),
	.seq_rdv_doing_rd_4(\seq_wrapper|seq_inst|seq_rdv_doing_rd[4]~q ),
	.seq_pll_inc_dec_n(\seq_wrapper|seq_inst|seq_pll_inc_dec_n~q ),
	.seq_pll_start_reconfig(\seq_wrapper|seq_inst|seq_pll_start_reconfig~q ),
	.seq_pll_select_2(\seq_wrapper|seq_inst|seq_pll_select[2]~q ),
	.seq_pll_select_1(\seq_wrapper|seq_inst|seq_pll_select[1]~q ),
	.seq_mem_clk_disable(\seq_wrapper|seq_inst|seq_mem_clk_disable~q ),
	.seq_rdata_valid_0(\rdv_pipe|seq_rdata_valid[0]~q ),
	.seq_rdata_valid_1(\rdv_pipe|seq_rdata_valid[1]~q ),
	.seq_ac_cs_n_0(\seq_wrapper|seq_inst|seq_ac_cs_n[0]~q ),
	.seq_ac_sel(\seq_wrapper|seq_inst|admin|seq_ac_sel~q ),
	.dgwb_wdp_ovride(\seq_wrapper|seq_inst|dgwb|dgwb_wdp_ovride~q ),
	.seq_wdp_ovride(\seq_wrapper|seq_inst|seq_wdp_ovride~0_combout ),
	.dgwb_wdata_120(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[120]~q ),
	.dgwb_wdata_56(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[56]~q ),
	.dgwb_wdata_88(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[88]~q ),
	.dgwb_wdata_24(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[24]~q ),
	.dgwb_wdata_121(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[121]~q ),
	.dgwb_wdata_57(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[57]~q ),
	.dgwb_wdata_89(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[89]~q ),
	.dgwb_wdata_25(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[25]~q ),
	.dgwb_wdata_122(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[122]~q ),
	.dgwb_wdata_58(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[58]~q ),
	.dgwb_wdata_90(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[90]~q ),
	.dgwb_wdata_26(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[26]~q ),
	.dgwb_wdata_123(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[123]~q ),
	.dgwb_wdata_59(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[59]~q ),
	.dgwb_wdata_91(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[91]~q ),
	.dgwb_wdata_27(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[27]~q ),
	.dgwb_wdata_124(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[124]~q ),
	.dgwb_wdata_60(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[60]~q ),
	.dgwb_wdata_92(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[92]~q ),
	.dgwb_wdata_28(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[28]~q ),
	.dgwb_wdata_125(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[125]~q ),
	.dgwb_wdata_61(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[61]~q ),
	.dgwb_wdata_93(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[93]~q ),
	.dgwb_wdata_29(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[29]~q ),
	.dgwb_wdata_126(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[126]~q ),
	.dgwb_wdata_62(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[62]~q ),
	.dgwb_wdata_94(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[94]~q ),
	.dgwb_wdata_30(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[30]~q ),
	.dgwb_wdata_127(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[127]~q ),
	.dgwb_wdata_63(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[63]~q ),
	.dgwb_wdata_95(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[95]~q ),
	.dgwb_wdata_31(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[31]~q ),
	.seq_poa_protection_override_1x(\seq_wrapper|seq_inst|seq_poa_protection_override_1x~q ),
	.seq_poa_lat_dec_1x_0(\seq_wrapper|seq_inst|seq_poa_lat_dec_1x[0]~q ),
	.mimic_done_out(\mmc|mimic_done_out~q ),
	.phs_shft_busy_siii(\clk|phs_shft_busy_siii~q ),
	.seq_mmc_start(\seq_wrapper|seq_inst|dgrb|seq_mmc_start~q ),
	.mimic_value_captured(\mmc|mimic_value_captured~q ),
	.GND_port(GND_port),
	.dgwb_wdp_ovride1(\seq_wrapper|seq_inst|dgwb|dgwb_wdp_ovride~_wirecell_combout ),
	.seq_ac_cas_n_0(\seq_wrapper|seq_inst|seq_ac_cas_n[0]~_wirecell_combout ),
	.seq_ac_cas_n_1(\seq_wrapper|seq_inst|seq_ac_cas_n[1]~_wirecell_combout ),
	.seq_ac_cs_n_1(\seq_wrapper|seq_inst|seq_ac_cs_n[1]~_wirecell_combout ),
	.seq_ac_ras_n_0(\seq_wrapper|seq_inst|seq_ac_ras_n[0]~_wirecell_combout ),
	.seq_ac_ras_n_1(\seq_wrapper|seq_inst|seq_ac_ras_n[1]~_wirecell_combout ),
	.seq_ac_we_n_0(\seq_wrapper|seq_inst|seq_ac_we_n[0]~_wirecell_combout ),
	.seq_ac_we_n_1(\seq_wrapper|seq_inst|seq_ac_we_n[1]~_wirecell_combout ));

ddr3_int_ddr3_int_phy_alt_mem_phy_write_dp \half_rate_wdp_gen.wdp (
	.phy_clk_1x(clk_0),
	.mem_clk_2x(clk_1),
	.write_clk_2x(\clk|half_rate.pll|altpll_component|auto_generated|clk[3] ),
	.wdp_dm_l_2x_0(\half_rate_wdp_gen.wdp|wdp_dm_l_2x[0]~q ),
	.wdp_dm_h_2x_0(\half_rate_wdp_gen.wdp|wdp_dm_h_2x[0]~q ),
	.wdp_dm_l_2x_1(\half_rate_wdp_gen.wdp|wdp_dm_l_2x[1]~q ),
	.wdp_dm_h_2x_1(\half_rate_wdp_gen.wdp|wdp_dm_h_2x[1]~q ),
	.wdp_dm_l_2x_2(\half_rate_wdp_gen.wdp|wdp_dm_l_2x[2]~q ),
	.wdp_dm_h_2x_2(\half_rate_wdp_gen.wdp|wdp_dm_h_2x[2]~q ),
	.wdp_dm_l_2x_3(\half_rate_wdp_gen.wdp|wdp_dm_l_2x[3]~q ),
	.wdp_dm_h_2x_3(\half_rate_wdp_gen.wdp|wdp_dm_h_2x[3]~q ),
	.wdp_wdata_l_2x_0(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[0]~q ),
	.wdp_wdata_h_2x_0(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[0]~q ),
	.dq_oe_2x_0(\half_rate_wdp_gen.wdp|dq_oe_2x[0]~q ),
	.wdp_wdata_l_2x_1(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[1]~q ),
	.wdp_wdata_h_2x_1(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[1]~q ),
	.wdp_wdata_l_2x_2(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[2]~q ),
	.wdp_wdata_h_2x_2(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[2]~q ),
	.wdp_wdata_l_2x_3(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[3]~q ),
	.wdp_wdata_h_2x_3(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[3]~q ),
	.wdp_wdata_l_2x_4(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[4]~q ),
	.wdp_wdata_h_2x_4(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[4]~q ),
	.dq_oe_2x_1(\half_rate_wdp_gen.wdp|dq_oe_2x[1]~q ),
	.wdp_wdata_l_2x_5(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[5]~q ),
	.wdp_wdata_h_2x_5(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[5]~q ),
	.wdp_wdata_l_2x_6(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[6]~q ),
	.wdp_wdata_h_2x_6(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[6]~q ),
	.wdp_wdata_l_2x_7(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[7]~q ),
	.wdp_wdata_h_2x_7(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[7]~q ),
	.wdp_wdata_l_2x_8(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[8]~q ),
	.wdp_wdata_h_2x_8(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[8]~q ),
	.dq_oe_2x_2(\half_rate_wdp_gen.wdp|dq_oe_2x[2]~q ),
	.wdp_wdata_l_2x_9(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[9]~q ),
	.wdp_wdata_h_2x_9(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[9]~q ),
	.wdp_wdata_l_2x_10(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[10]~q ),
	.wdp_wdata_h_2x_10(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[10]~q ),
	.wdp_wdata_l_2x_11(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[11]~q ),
	.wdp_wdata_h_2x_11(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[11]~q ),
	.wdp_wdata_l_2x_12(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[12]~q ),
	.wdp_wdata_h_2x_12(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[12]~q ),
	.dq_oe_2x_3(\half_rate_wdp_gen.wdp|dq_oe_2x[3]~q ),
	.wdp_wdata_l_2x_13(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[13]~q ),
	.wdp_wdata_h_2x_13(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[13]~q ),
	.wdp_wdata_l_2x_14(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[14]~q ),
	.wdp_wdata_h_2x_14(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[14]~q ),
	.wdp_wdata_l_2x_15(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[15]~q ),
	.wdp_wdata_h_2x_15(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[15]~q ),
	.wdp_wdata_l_2x_16(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[16]~q ),
	.wdp_wdata_h_2x_16(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[16]~q ),
	.dq_oe_2x_4(\half_rate_wdp_gen.wdp|dq_oe_2x[4]~q ),
	.wdp_wdata_l_2x_17(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[17]~q ),
	.wdp_wdata_h_2x_17(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[17]~q ),
	.wdp_wdata_l_2x_18(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[18]~q ),
	.wdp_wdata_h_2x_18(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[18]~q ),
	.wdp_wdata_l_2x_19(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[19]~q ),
	.wdp_wdata_h_2x_19(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[19]~q ),
	.wdp_wdata_l_2x_20(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[20]~q ),
	.wdp_wdata_h_2x_20(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[20]~q ),
	.dq_oe_2x_5(\half_rate_wdp_gen.wdp|dq_oe_2x[5]~q ),
	.wdp_wdata_l_2x_21(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[21]~q ),
	.wdp_wdata_h_2x_21(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[21]~q ),
	.wdp_wdata_l_2x_22(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[22]~q ),
	.wdp_wdata_h_2x_22(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[22]~q ),
	.wdp_wdata_l_2x_23(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[23]~q ),
	.wdp_wdata_h_2x_23(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[23]~q ),
	.wdp_wdata_l_2x_24(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[24]~q ),
	.wdp_wdata_h_2x_24(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[24]~q ),
	.dq_oe_2x_6(\half_rate_wdp_gen.wdp|dq_oe_2x[6]~q ),
	.wdp_wdata_l_2x_25(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[25]~q ),
	.wdp_wdata_h_2x_25(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[25]~q ),
	.wdp_wdata_l_2x_26(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[26]~q ),
	.wdp_wdata_h_2x_26(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[26]~q ),
	.wdp_wdata_l_2x_27(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[27]~q ),
	.wdp_wdata_h_2x_27(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[27]~q ),
	.wdp_wdata_l_2x_28(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[28]~q ),
	.wdp_wdata_h_2x_28(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[28]~q ),
	.dq_oe_2x_7(\half_rate_wdp_gen.wdp|dq_oe_2x[7]~q ),
	.wdp_wdata_l_2x_29(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[29]~q ),
	.wdp_wdata_h_2x_29(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[29]~q ),
	.wdp_wdata_l_2x_30(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[30]~q ),
	.wdp_wdata_h_2x_30(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[30]~q ),
	.wdp_wdata_l_2x_31(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[31]~q ),
	.wdp_wdata_h_2x_31(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[31]~q ),
	.q_b_96(q_b_961),
	.q_b_32(q_b_321),
	.q_b_64(q_b_641),
	.q_b_0(q_b_01),
	.q_b_97(q_b_971),
	.q_b_33(q_b_331),
	.q_b_65(q_b_651),
	.q_b_1(q_b_128),
	.q_b_98(q_b_981),
	.q_b_34(q_b_341),
	.q_b_66(q_b_661),
	.q_b_2(q_b_210),
	.q_b_99(q_b_991),
	.q_b_35(q_b_351),
	.q_b_67(q_b_671),
	.q_b_3(q_b_310),
	.q_b_100(q_b_1001),
	.q_b_36(q_b_361),
	.q_b_68(q_b_681),
	.q_b_4(q_b_410),
	.q_b_101(q_b_1011),
	.q_b_37(q_b_371),
	.q_b_69(q_b_691),
	.q_b_5(q_b_510),
	.q_b_102(q_b_1021),
	.q_b_38(q_b_381),
	.q_b_70(q_b_701),
	.q_b_6(q_b_610),
	.q_b_103(q_b_1031),
	.q_b_39(q_b_391),
	.q_b_71(q_b_711),
	.q_b_7(q_b_710),
	.q_b_104(q_b_1041),
	.q_b_40(q_b_401),
	.q_b_72(q_b_721),
	.q_b_8(q_b_810),
	.q_b_105(q_b_1051),
	.q_b_41(q_b_411),
	.q_b_73(q_b_731),
	.q_b_9(q_b_910),
	.q_b_106(q_b_1061),
	.q_b_42(q_b_421),
	.q_b_74(q_b_741),
	.q_b_10(q_b_1010),
	.q_b_107(q_b_1071),
	.q_b_43(q_b_431),
	.q_b_75(q_b_751),
	.q_b_11(q_b_1110),
	.q_b_108(q_b_1081),
	.q_b_44(q_b_441),
	.q_b_76(q_b_761),
	.q_b_12(q_b_129),
	.q_b_109(q_b_1091),
	.q_b_45(q_b_451),
	.q_b_77(q_b_771),
	.q_b_13(q_b_131),
	.q_b_110(q_b_1101),
	.q_b_46(q_b_461),
	.q_b_78(q_b_781),
	.q_b_14(q_b_141),
	.q_b_111(q_b_1111),
	.q_b_47(q_b_471),
	.q_b_79(q_b_791),
	.q_b_15(q_b_151),
	.q_b_112(q_b_1121),
	.q_b_48(q_b_481),
	.q_b_80(q_b_801),
	.q_b_16(q_b_161),
	.q_b_113(q_b_1131),
	.q_b_49(q_b_491),
	.q_b_81(q_b_811),
	.q_b_17(q_b_171),
	.q_b_114(q_b_1141),
	.q_b_50(q_b_501),
	.q_b_82(q_b_821),
	.q_b_18(q_b_181),
	.q_b_115(q_b_1151),
	.q_b_51(q_b_511),
	.q_b_83(q_b_831),
	.q_b_19(q_b_191),
	.q_b_116(q_b_1161),
	.q_b_52(q_b_521),
	.q_b_84(q_b_841),
	.q_b_20(q_b_201),
	.q_b_117(q_b_1171),
	.q_b_53(q_b_531),
	.q_b_85(q_b_851),
	.q_b_21(q_b_211),
	.q_b_118(q_b_1181),
	.q_b_54(q_b_541),
	.q_b_86(q_b_861),
	.q_b_22(q_b_221),
	.q_b_119(q_b_1191),
	.q_b_55(q_b_551),
	.q_b_87(q_b_871),
	.q_b_23(q_b_231),
	.q_b_120(q_b_1201),
	.q_b_56(q_b_561),
	.q_b_88(q_b_881),
	.q_b_24(q_b_241),
	.q_b_121(q_b_1211),
	.q_b_57(q_b_571),
	.q_b_89(q_b_891),
	.q_b_25(q_b_251),
	.q_b_122(q_b_1221),
	.q_b_58(q_b_581),
	.q_b_90(q_b_901),
	.q_b_26(q_b_261),
	.q_b_123(q_b_1231),
	.q_b_59(q_b_591),
	.q_b_91(q_b_911),
	.q_b_27(q_b_271),
	.q_b_124(q_b_1241),
	.q_b_60(q_b_601),
	.q_b_92(q_b_921),
	.q_b_28(q_b_281),
	.q_b_125(q_b_1251),
	.q_b_61(q_b_611),
	.q_b_93(q_b_931),
	.q_b_29(q_b_291),
	.q_b_126(q_b_1261),
	.q_b_62(q_b_621),
	.q_b_94(q_b_941),
	.q_b_30(q_b_301),
	.q_b_127(q_b_1271),
	.q_b_63(q_b_631),
	.q_b_95(q_b_951),
	.q_b_31(q_b_311),
	.reset_phy_clk_1x_n(reset_phy_clk_1x_n),
	.ctl_init_fail(\seq_wrapper|seq_inst|ctrl|ctl_init_fail~q ),
	.ctl_init_success(\seq_wrapper|seq_inst|ctrl|ctl_init_success~q ),
	.reset_write_clk_2x_n(\clk|write_clk_pipe|ams_pipe[3]~q ),
	.dqs_burst_2x_r3_0(\half_rate_wdp_gen.wdp|dqs_burst_2x_r3[0]~q ),
	.dqs_burst_2x_r3_1(\half_rate_wdp_gen.wdp|dqs_burst_2x_r3[1]~q ),
	.dqs_burst_2x_r3_2(\half_rate_wdp_gen.wdp|dqs_burst_2x_r3[2]~q ),
	.dqs_burst_2x_r3_3(\half_rate_wdp_gen.wdp|dqs_burst_2x_r3[3]~q ),
	.reset_mem_clk_2x_n(\clk|mem_clk_pipe|ams_pipe[3]~q ),
	.afi_dm_4(afi_dm_4),
	.dgwb_wdp_ovride(\seq_wrapper|seq_inst|dgwb|dgwb_wdp_ovride~q ),
	.seq_wdp_ovride(\seq_wrapper|seq_inst|seq_wdp_ovride~0_combout ),
	.afi_dm_12(afi_dm_12),
	.afi_dm_0(afi_dm_0),
	.afi_dm_8(afi_dm_8),
	.afi_dm_5(afi_dm_5),
	.afi_dm_13(afi_dm_13),
	.afi_dm_1(afi_dm_1),
	.afi_dm_9(afi_dm_9),
	.afi_dm_6(afi_dm_6),
	.afi_dm_14(afi_dm_14),
	.afi_dm_2(afi_dm_2),
	.afi_dm_10(afi_dm_10),
	.afi_dm_7(afi_dm_7),
	.afi_dm_15(afi_dm_15),
	.afi_dm_3(afi_dm_3),
	.afi_dm_11(afi_dm_11),
	.int_wdata_valid(int_wdata_valid),
	.dgwb_wdata_120(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[120]~q ),
	.dgwb_wdata_56(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[56]~q ),
	.dgwb_wdata_88(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[88]~q ),
	.dgwb_wdata_24(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[24]~q ),
	.dgwb_wdata_121(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[121]~q ),
	.dgwb_wdata_57(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[57]~q ),
	.dgwb_wdata_89(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[89]~q ),
	.dgwb_wdata_25(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[25]~q ),
	.dgwb_wdata_122(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[122]~q ),
	.dgwb_wdata_58(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[58]~q ),
	.dgwb_wdata_90(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[90]~q ),
	.dgwb_wdata_26(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[26]~q ),
	.dgwb_wdata_123(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[123]~q ),
	.dgwb_wdata_59(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[59]~q ),
	.dgwb_wdata_91(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[91]~q ),
	.dgwb_wdata_27(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[27]~q ),
	.dgwb_wdata_124(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[124]~q ),
	.dgwb_wdata_60(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[60]~q ),
	.dgwb_wdata_92(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[92]~q ),
	.dgwb_wdata_28(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[28]~q ),
	.dgwb_wdata_125(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[125]~q ),
	.dgwb_wdata_61(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[61]~q ),
	.dgwb_wdata_93(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[93]~q ),
	.dgwb_wdata_29(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[29]~q ),
	.dgwb_wdata_126(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[126]~q ),
	.dgwb_wdata_62(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[62]~q ),
	.dgwb_wdata_94(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[94]~q ),
	.dgwb_wdata_30(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[30]~q ),
	.dgwb_wdata_127(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[127]~q ),
	.dgwb_wdata_63(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[63]~q ),
	.dgwb_wdata_95(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[95]~q ),
	.dgwb_wdata_31(\seq_wrapper|seq_inst|dgwb|dgwb_wdata[31]~q ),
	.int_dqs_burst(int_dqs_burst),
	.int_dqs_burst_hr(int_dqs_burst_hr),
	.dgwb_wdp_ovride1(\seq_wrapper|seq_inst|dgwb|dgwb_wdp_ovride~_wirecell_combout ));

ddr3_int_ddr3_int_phy_alt_mem_phy_addr_cmd \half_rate_adc_gen.adc (
	.clk_0(clk_0),
	.clk_3(\clk|half_rate.pll|altpll_component|auto_generated|clk[3] ),
	.dataout_0(dataout_0),
	.dataout_01(dataout_01),
	.dataout_02(dataout_02),
	.dataout_03(dataout_03),
	.dataout_04(dataout_04),
	.dataout_05(dataout_05),
	.dataout_06(dataout_06),
	.dataout_07(dataout_07),
	.dataout_08(dataout_08),
	.dataout_09(dataout_09),
	.dataout_010(dataout_010),
	.dataout_011(dataout_011),
	.dataout_012(dataout_012),
	.dataout_013(dataout_013),
	.dataout_014(dataout_014),
	.dataout_015(dataout_015),
	.dataout_016(dataout_016),
	.dataout_017(dataout_017),
	.dataout_018(dataout_018),
	.dataout_019(dataout_019),
	.dataout_020(dataout_020),
	.dataout_021(dataout_021),
	.dataout_022(dataout_022),
	.dataout_023(dataout_023),
	.seq_ac_cke_1(\seq_wrapper|seq_inst|seq_ac_cke[1]~q ),
	.seq_ac_addr_0(\seq_wrapper|seq_inst|seq_ac_addr[0]~q ),
	.seq_ac_addr_14(\seq_wrapper|seq_inst|seq_ac_addr[14]~q ),
	.seq_ac_addr_1(\seq_wrapper|seq_inst|seq_ac_addr[1]~q ),
	.seq_ac_addr_15(\seq_wrapper|seq_inst|seq_ac_addr[15]~q ),
	.seq_ac_addr_16(\seq_wrapper|seq_inst|seq_ac_addr[16]~q ),
	.seq_ac_addr_17(\seq_wrapper|seq_inst|seq_ac_addr[17]~q ),
	.seq_ac_addr_18(\seq_wrapper|seq_inst|seq_ac_addr[18]~q ),
	.seq_ac_addr_5(\seq_wrapper|seq_inst|seq_ac_addr[5]~q ),
	.seq_ac_addr_19(\seq_wrapper|seq_inst|seq_ac_addr[19]~q ),
	.seq_ac_addr_8(\seq_wrapper|seq_inst|seq_ac_addr[8]~q ),
	.seq_ac_addr_22(\seq_wrapper|seq_inst|seq_ac_addr[22]~q ),
	.seq_ac_addr_10(\seq_wrapper|seq_inst|seq_ac_addr[10]~q ),
	.seq_ac_addr_24(\seq_wrapper|seq_inst|seq_ac_addr[24]~q ),
	.seq_ac_addr_12(\seq_wrapper|seq_inst|seq_ac_addr[12]~q ),
	.seq_ac_addr_26(\seq_wrapper|seq_inst|seq_ac_addr[26]~q ),
	.seq_ac_ba_0(\seq_wrapper|seq_inst|seq_ac_ba[0]~q ),
	.seq_ac_ba_3(\seq_wrapper|seq_inst|seq_ac_ba[3]~q ),
	.seq_ac_ba_1(\seq_wrapper|seq_inst|seq_ac_ba[1]~q ),
	.seq_ac_ba_4(\seq_wrapper|seq_inst|seq_ac_ba[4]~q ),
	.seq_ac_rst_n_0(\seq_wrapper|seq_inst|seq_ac_rst_n[0]~q ),
	.ams_pipe_1(\clk|ac_clk_pipe_2x|ams_pipe[1]~q ),
	.seq_ac_add_1t_ac_lat_internal(\seq_wrapper|seq_inst|seq_ac_add_1t_ac_lat_internal~q ),
	.seq_ac_cs_n_0(\seq_wrapper|seq_inst|seq_ac_cs_n[0]~q ),
	.seq_ac_sel(\seq_wrapper|seq_inst|admin|seq_ac_sel~q ),
	.afi_cs_n_1(afi_cs_n_1),
	.int_cke_r_0(int_cke_r_0),
	.afi_addr_0(afi_addr_0),
	.afi_addr_1(afi_addr_1),
	.afi_addr_2(afi_addr_2),
	.afi_addr_3(afi_addr_3),
	.afi_addr_4(afi_addr_4),
	.afi_addr_5(afi_addr_5),
	.afi_addr_6(afi_addr_6),
	.afi_addr_7(afi_addr_7),
	.afi_addr_8(afi_addr_8),
	.afi_addr_9(afi_addr_9),
	.afi_addr_10(afi_addr_10),
	.afi_addr_11(afi_addr_11),
	.afi_addr_12(afi_addr_12),
	.afi_addr_13(afi_addr_13),
	.afi_ba_0(afi_ba_0),
	.afi_ba_1(afi_ba_1),
	.afi_ba_2(afi_ba_2),
	.afi_ras_n_0(afi_ras_n_0),
	.afi_cas_n_0(afi_cas_n_0),
	.afi_we_n_0(afi_we_n_0),
	.GND_port(GND_port),
	.seq_ac_cas_n_0(\seq_wrapper|seq_inst|seq_ac_cas_n[0]~_wirecell_combout ),
	.seq_ac_cas_n_1(\seq_wrapper|seq_inst|seq_ac_cas_n[1]~_wirecell_combout ),
	.seq_ac_cs_n_1(\seq_wrapper|seq_inst|seq_ac_cs_n[1]~_wirecell_combout ),
	.seq_ac_ras_n_0(\seq_wrapper|seq_inst|seq_ac_ras_n[0]~_wirecell_combout ),
	.seq_ac_ras_n_1(\seq_wrapper|seq_inst|seq_ac_ras_n[1]~_wirecell_combout ),
	.seq_ac_we_n_0(\seq_wrapper|seq_inst|seq_ac_we_n[0]~_wirecell_combout ),
	.seq_ac_we_n_1(\seq_wrapper|seq_inst|seq_ac_we_n[1]~_wirecell_combout ));

ddr3_int_ddr3_int_phy_alt_mem_phy_dp_io dpio(
	.clk_1(clk_1),
	.clk_3(\clk|half_rate.pll|altpll_component|auto_generated|clk[3] ),
	.resync_clk_2x(\clk|half_rate.pll|altpll_component|auto_generated|clk[4] ),
	.dqs_delay_ctrl_0(dqs_delay_ctrl_0),
	.dqs_delay_ctrl_1(dqs_delay_ctrl_1),
	.dqs_delay_ctrl_2(dqs_delay_ctrl_2),
	.dqs_delay_ctrl_3(dqs_delay_ctrl_3),
	.dqs_delay_ctrl_4(dqs_delay_ctrl_4),
	.dqs_delay_ctrl_5(dqs_delay_ctrl_5),
	.wire_output_dq_0_output_ddio_out_inst_dataout(wire_output_dq_0_output_ddio_out_inst_dataout),
	.wire_output_dq_0_output_ddio_out_inst_dataout1(wire_output_dq_0_output_ddio_out_inst_dataout1),
	.wire_output_dq_0_output_ddio_out_inst_dataout2(wire_output_dq_0_output_ddio_out_inst_dataout2),
	.wire_output_dq_0_output_ddio_out_inst_dataout3(wire_output_dq_0_output_ddio_out_inst_dataout3),
	.wdp_dm_l_2x_0(\half_rate_wdp_gen.wdp|wdp_dm_l_2x[0]~q ),
	.wdp_dm_h_2x_0(\half_rate_wdp_gen.wdp|wdp_dm_h_2x[0]~q ),
	.wdp_dm_l_2x_1(\half_rate_wdp_gen.wdp|wdp_dm_l_2x[1]~q ),
	.wdp_dm_h_2x_1(\half_rate_wdp_gen.wdp|wdp_dm_h_2x[1]~q ),
	.wdp_dm_l_2x_2(\half_rate_wdp_gen.wdp|wdp_dm_l_2x[2]~q ),
	.wdp_dm_h_2x_2(\half_rate_wdp_gen.wdp|wdp_dm_h_2x[2]~q ),
	.wdp_dm_l_2x_3(\half_rate_wdp_gen.wdp|wdp_dm_l_2x[3]~q ),
	.wdp_dm_h_2x_3(\half_rate_wdp_gen.wdp|wdp_dm_h_2x[3]~q ),
	.wire_bidir_dq_0_output_ddio_out_inst_dataout(wire_bidir_dq_0_output_ddio_out_inst_dataout),
	.wire_bidir_dq_1_output_ddio_out_inst_dataout(wire_bidir_dq_1_output_ddio_out_inst_dataout),
	.wire_bidir_dq_2_output_ddio_out_inst_dataout(wire_bidir_dq_2_output_ddio_out_inst_dataout),
	.wire_bidir_dq_3_output_ddio_out_inst_dataout(wire_bidir_dq_3_output_ddio_out_inst_dataout),
	.wire_bidir_dq_4_output_ddio_out_inst_dataout(wire_bidir_dq_4_output_ddio_out_inst_dataout),
	.wire_bidir_dq_5_output_ddio_out_inst_dataout(wire_bidir_dq_5_output_ddio_out_inst_dataout),
	.wire_bidir_dq_6_output_ddio_out_inst_dataout(wire_bidir_dq_6_output_ddio_out_inst_dataout),
	.wire_bidir_dq_7_output_ddio_out_inst_dataout(wire_bidir_dq_7_output_ddio_out_inst_dataout),
	.wire_bidir_dq_0_output_ddio_out_inst_dataout1(wire_bidir_dq_0_output_ddio_out_inst_dataout1),
	.wire_bidir_dq_1_output_ddio_out_inst_dataout1(wire_bidir_dq_1_output_ddio_out_inst_dataout1),
	.wire_bidir_dq_2_output_ddio_out_inst_dataout1(wire_bidir_dq_2_output_ddio_out_inst_dataout1),
	.wire_bidir_dq_3_output_ddio_out_inst_dataout1(wire_bidir_dq_3_output_ddio_out_inst_dataout1),
	.wire_bidir_dq_4_output_ddio_out_inst_dataout1(wire_bidir_dq_4_output_ddio_out_inst_dataout1),
	.wire_bidir_dq_5_output_ddio_out_inst_dataout1(wire_bidir_dq_5_output_ddio_out_inst_dataout1),
	.wire_bidir_dq_6_output_ddio_out_inst_dataout1(wire_bidir_dq_6_output_ddio_out_inst_dataout1),
	.wire_bidir_dq_7_output_ddio_out_inst_dataout1(wire_bidir_dq_7_output_ddio_out_inst_dataout1),
	.wire_bidir_dq_0_output_ddio_out_inst_dataout2(wire_bidir_dq_0_output_ddio_out_inst_dataout2),
	.wire_bidir_dq_1_output_ddio_out_inst_dataout2(wire_bidir_dq_1_output_ddio_out_inst_dataout2),
	.wire_bidir_dq_2_output_ddio_out_inst_dataout2(wire_bidir_dq_2_output_ddio_out_inst_dataout2),
	.wire_bidir_dq_3_output_ddio_out_inst_dataout2(wire_bidir_dq_3_output_ddio_out_inst_dataout2),
	.wire_bidir_dq_4_output_ddio_out_inst_dataout2(wire_bidir_dq_4_output_ddio_out_inst_dataout2),
	.wire_bidir_dq_5_output_ddio_out_inst_dataout2(wire_bidir_dq_5_output_ddio_out_inst_dataout2),
	.wire_bidir_dq_6_output_ddio_out_inst_dataout2(wire_bidir_dq_6_output_ddio_out_inst_dataout2),
	.wire_bidir_dq_7_output_ddio_out_inst_dataout2(wire_bidir_dq_7_output_ddio_out_inst_dataout2),
	.wire_bidir_dq_0_output_ddio_out_inst_dataout3(wire_bidir_dq_0_output_ddio_out_inst_dataout3),
	.wire_bidir_dq_1_output_ddio_out_inst_dataout3(wire_bidir_dq_1_output_ddio_out_inst_dataout3),
	.wire_bidir_dq_2_output_ddio_out_inst_dataout3(wire_bidir_dq_2_output_ddio_out_inst_dataout3),
	.wire_bidir_dq_3_output_ddio_out_inst_dataout3(wire_bidir_dq_3_output_ddio_out_inst_dataout3),
	.wire_bidir_dq_4_output_ddio_out_inst_dataout3(wire_bidir_dq_4_output_ddio_out_inst_dataout3),
	.wire_bidir_dq_5_output_ddio_out_inst_dataout3(wire_bidir_dq_5_output_ddio_out_inst_dataout3),
	.wire_bidir_dq_6_output_ddio_out_inst_dataout3(wire_bidir_dq_6_output_ddio_out_inst_dataout3),
	.wire_bidir_dq_7_output_ddio_out_inst_dataout3(wire_bidir_dq_7_output_ddio_out_inst_dataout3),
	.dqs_pseudo_diff_out_0(dqs_pseudo_diff_out_0),
	.dqsn_pseudo_diff_out_0(dqsn_pseudo_diff_out_0),
	.dqs_pseudo_diff_out_1(dqs_pseudo_diff_out_1),
	.dqsn_pseudo_diff_out_1(dqsn_pseudo_diff_out_1),
	.dqs_pseudo_diff_out_2(dqs_pseudo_diff_out_2),
	.dqsn_pseudo_diff_out_2(dqsn_pseudo_diff_out_2),
	.dqs_pseudo_diff_out_3(dqs_pseudo_diff_out_3),
	.dqsn_pseudo_diff_out_3(dqsn_pseudo_diff_out_3),
	.wdp_wdata_l_2x_0(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[0]~q ),
	.wdp_wdata_h_2x_0(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[0]~q ),
	.dq_oe_2x_0(\half_rate_wdp_gen.wdp|dq_oe_2x[0]~q ),
	.wdp_wdata_l_2x_1(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[1]~q ),
	.wdp_wdata_h_2x_1(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[1]~q ),
	.wdp_wdata_l_2x_2(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[2]~q ),
	.wdp_wdata_h_2x_2(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[2]~q ),
	.wdp_wdata_l_2x_3(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[3]~q ),
	.wdp_wdata_h_2x_3(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[3]~q ),
	.wdp_wdata_l_2x_4(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[4]~q ),
	.wdp_wdata_h_2x_4(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[4]~q ),
	.dq_oe_2x_1(\half_rate_wdp_gen.wdp|dq_oe_2x[1]~q ),
	.wdp_wdata_l_2x_5(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[5]~q ),
	.wdp_wdata_h_2x_5(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[5]~q ),
	.wdp_wdata_l_2x_6(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[6]~q ),
	.wdp_wdata_h_2x_6(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[6]~q ),
	.wdp_wdata_l_2x_7(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[7]~q ),
	.wdp_wdata_h_2x_7(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[7]~q ),
	.wdp_wdata_l_2x_8(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[8]~q ),
	.wdp_wdata_h_2x_8(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[8]~q ),
	.dq_oe_2x_2(\half_rate_wdp_gen.wdp|dq_oe_2x[2]~q ),
	.wdp_wdata_l_2x_9(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[9]~q ),
	.wdp_wdata_h_2x_9(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[9]~q ),
	.wdp_wdata_l_2x_10(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[10]~q ),
	.wdp_wdata_h_2x_10(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[10]~q ),
	.wdp_wdata_l_2x_11(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[11]~q ),
	.wdp_wdata_h_2x_11(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[11]~q ),
	.wdp_wdata_l_2x_12(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[12]~q ),
	.wdp_wdata_h_2x_12(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[12]~q ),
	.dq_oe_2x_3(\half_rate_wdp_gen.wdp|dq_oe_2x[3]~q ),
	.wdp_wdata_l_2x_13(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[13]~q ),
	.wdp_wdata_h_2x_13(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[13]~q ),
	.wdp_wdata_l_2x_14(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[14]~q ),
	.wdp_wdata_h_2x_14(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[14]~q ),
	.wdp_wdata_l_2x_15(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[15]~q ),
	.wdp_wdata_h_2x_15(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[15]~q ),
	.wdp_wdata_l_2x_16(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[16]~q ),
	.wdp_wdata_h_2x_16(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[16]~q ),
	.dq_oe_2x_4(\half_rate_wdp_gen.wdp|dq_oe_2x[4]~q ),
	.wdp_wdata_l_2x_17(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[17]~q ),
	.wdp_wdata_h_2x_17(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[17]~q ),
	.wdp_wdata_l_2x_18(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[18]~q ),
	.wdp_wdata_h_2x_18(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[18]~q ),
	.wdp_wdata_l_2x_19(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[19]~q ),
	.wdp_wdata_h_2x_19(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[19]~q ),
	.wdp_wdata_l_2x_20(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[20]~q ),
	.wdp_wdata_h_2x_20(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[20]~q ),
	.dq_oe_2x_5(\half_rate_wdp_gen.wdp|dq_oe_2x[5]~q ),
	.wdp_wdata_l_2x_21(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[21]~q ),
	.wdp_wdata_h_2x_21(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[21]~q ),
	.wdp_wdata_l_2x_22(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[22]~q ),
	.wdp_wdata_h_2x_22(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[22]~q ),
	.wdp_wdata_l_2x_23(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[23]~q ),
	.wdp_wdata_h_2x_23(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[23]~q ),
	.wdp_wdata_l_2x_24(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[24]~q ),
	.wdp_wdata_h_2x_24(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[24]~q ),
	.dq_oe_2x_6(\half_rate_wdp_gen.wdp|dq_oe_2x[6]~q ),
	.wdp_wdata_l_2x_25(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[25]~q ),
	.wdp_wdata_h_2x_25(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[25]~q ),
	.wdp_wdata_l_2x_26(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[26]~q ),
	.wdp_wdata_h_2x_26(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[26]~q ),
	.wdp_wdata_l_2x_27(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[27]~q ),
	.wdp_wdata_h_2x_27(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[27]~q ),
	.wdp_wdata_l_2x_28(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[28]~q ),
	.wdp_wdata_h_2x_28(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[28]~q ),
	.dq_oe_2x_7(\half_rate_wdp_gen.wdp|dq_oe_2x[7]~q ),
	.wdp_wdata_l_2x_29(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[29]~q ),
	.wdp_wdata_h_2x_29(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[29]~q ),
	.wdp_wdata_l_2x_30(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[30]~q ),
	.wdp_wdata_h_2x_30(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[30]~q ),
	.wdp_wdata_l_2x_31(\half_rate_wdp_gen.wdp|wdp_wdata_l_2x[31]~q ),
	.wdp_wdata_h_2x_31(\half_rate_wdp_gen.wdp|wdp_wdata_h_2x[31]~q ),
	.dq_datain_0(dq_datain_0),
	.dq_datain_1(dq_datain_1),
	.dq_datain_2(dq_datain_2),
	.dq_datain_3(dq_datain_3),
	.dq_datain_4(dq_datain_4),
	.dq_datain_5(dq_datain_5),
	.dq_datain_6(dq_datain_6),
	.dq_datain_7(dq_datain_7),
	.dq_datain_8(dq_datain_8),
	.dq_datain_9(dq_datain_9),
	.dq_datain_10(dq_datain_10),
	.dq_datain_11(dq_datain_11),
	.dq_datain_12(dq_datain_12),
	.dq_datain_13(dq_datain_13),
	.dq_datain_14(dq_datain_14),
	.dq_datain_15(dq_datain_15),
	.dq_datain_16(dq_datain_16),
	.dq_datain_17(dq_datain_17),
	.dq_datain_18(dq_datain_18),
	.dq_datain_19(dq_datain_19),
	.dq_datain_20(dq_datain_20),
	.dq_datain_21(dq_datain_21),
	.dq_datain_22(dq_datain_22),
	.dq_datain_23(dq_datain_23),
	.dq_datain_24(dq_datain_24),
	.dq_datain_25(dq_datain_25),
	.dq_datain_26(dq_datain_26),
	.dq_datain_27(dq_datain_27),
	.dq_datain_28(dq_datain_28),
	.dq_datain_29(dq_datain_29),
	.dq_datain_30(dq_datain_30),
	.dq_datain_31(dq_datain_31),
	.dqs_buffered_0(dqs_buffered_0),
	.dqs_buffered_1(dqs_buffered_1),
	.dqs_buffered_2(dqs_buffered_2),
	.dqs_buffered_3(dqs_buffered_3),
	.dio_rdata_h_2x_0(\dpio|dio_rdata_h_2x[0]~q ),
	.dio_rdata_h_2x_1(\dpio|dio_rdata_h_2x[1]~q ),
	.dio_rdata_h_2x_2(\dpio|dio_rdata_h_2x[2]~q ),
	.dio_rdata_h_2x_3(\dpio|dio_rdata_h_2x[3]~q ),
	.dio_rdata_h_2x_4(\dpio|dio_rdata_h_2x[4]~q ),
	.dio_rdata_h_2x_5(\dpio|dio_rdata_h_2x[5]~q ),
	.dio_rdata_h_2x_6(\dpio|dio_rdata_h_2x[6]~q ),
	.dio_rdata_h_2x_7(\dpio|dio_rdata_h_2x[7]~q ),
	.dio_rdata_h_2x_8(\dpio|dio_rdata_h_2x[8]~q ),
	.dio_rdata_h_2x_9(\dpio|dio_rdata_h_2x[9]~q ),
	.dio_rdata_h_2x_10(\dpio|dio_rdata_h_2x[10]~q ),
	.dio_rdata_h_2x_11(\dpio|dio_rdata_h_2x[11]~q ),
	.dio_rdata_h_2x_12(\dpio|dio_rdata_h_2x[12]~q ),
	.dio_rdata_h_2x_13(\dpio|dio_rdata_h_2x[13]~q ),
	.dio_rdata_h_2x_14(\dpio|dio_rdata_h_2x[14]~q ),
	.dio_rdata_h_2x_15(\dpio|dio_rdata_h_2x[15]~q ),
	.dio_rdata_h_2x_16(\dpio|dio_rdata_h_2x[16]~q ),
	.dio_rdata_h_2x_17(\dpio|dio_rdata_h_2x[17]~q ),
	.dio_rdata_h_2x_18(\dpio|dio_rdata_h_2x[18]~q ),
	.dio_rdata_h_2x_19(\dpio|dio_rdata_h_2x[19]~q ),
	.dio_rdata_h_2x_20(\dpio|dio_rdata_h_2x[20]~q ),
	.dio_rdata_h_2x_21(\dpio|dio_rdata_h_2x[21]~q ),
	.dio_rdata_h_2x_22(\dpio|dio_rdata_h_2x[22]~q ),
	.dio_rdata_h_2x_23(\dpio|dio_rdata_h_2x[23]~q ),
	.dio_rdata_h_2x_24(\dpio|dio_rdata_h_2x[24]~q ),
	.dio_rdata_h_2x_25(\dpio|dio_rdata_h_2x[25]~q ),
	.dio_rdata_h_2x_26(\dpio|dio_rdata_h_2x[26]~q ),
	.dio_rdata_h_2x_27(\dpio|dio_rdata_h_2x[27]~q ),
	.dio_rdata_h_2x_28(\dpio|dio_rdata_h_2x[28]~q ),
	.dio_rdata_h_2x_29(\dpio|dio_rdata_h_2x[29]~q ),
	.dio_rdata_h_2x_30(\dpio|dio_rdata_h_2x[30]~q ),
	.dio_rdata_h_2x_31(\dpio|dio_rdata_h_2x[31]~q ),
	.dio_rdata_l_2x_0(\dpio|dio_rdata_l_2x[0]~q ),
	.dio_rdata_l_2x_1(\dpio|dio_rdata_l_2x[1]~q ),
	.dio_rdata_l_2x_2(\dpio|dio_rdata_l_2x[2]~q ),
	.dio_rdata_l_2x_3(\dpio|dio_rdata_l_2x[3]~q ),
	.dio_rdata_l_2x_4(\dpio|dio_rdata_l_2x[4]~q ),
	.dio_rdata_l_2x_5(\dpio|dio_rdata_l_2x[5]~q ),
	.dio_rdata_l_2x_6(\dpio|dio_rdata_l_2x[6]~q ),
	.dio_rdata_l_2x_7(\dpio|dio_rdata_l_2x[7]~q ),
	.dio_rdata_l_2x_8(\dpio|dio_rdata_l_2x[8]~q ),
	.dio_rdata_l_2x_9(\dpio|dio_rdata_l_2x[9]~q ),
	.dio_rdata_l_2x_10(\dpio|dio_rdata_l_2x[10]~q ),
	.dio_rdata_l_2x_11(\dpio|dio_rdata_l_2x[11]~q ),
	.dio_rdata_l_2x_12(\dpio|dio_rdata_l_2x[12]~q ),
	.dio_rdata_l_2x_13(\dpio|dio_rdata_l_2x[13]~q ),
	.dio_rdata_l_2x_14(\dpio|dio_rdata_l_2x[14]~q ),
	.dio_rdata_l_2x_15(\dpio|dio_rdata_l_2x[15]~q ),
	.dio_rdata_l_2x_16(\dpio|dio_rdata_l_2x[16]~q ),
	.dio_rdata_l_2x_17(\dpio|dio_rdata_l_2x[17]~q ),
	.dio_rdata_l_2x_18(\dpio|dio_rdata_l_2x[18]~q ),
	.dio_rdata_l_2x_19(\dpio|dio_rdata_l_2x[19]~q ),
	.dio_rdata_l_2x_20(\dpio|dio_rdata_l_2x[20]~q ),
	.dio_rdata_l_2x_21(\dpio|dio_rdata_l_2x[21]~q ),
	.dio_rdata_l_2x_22(\dpio|dio_rdata_l_2x[22]~q ),
	.dio_rdata_l_2x_23(\dpio|dio_rdata_l_2x[23]~q ),
	.dio_rdata_l_2x_24(\dpio|dio_rdata_l_2x[24]~q ),
	.dio_rdata_l_2x_25(\dpio|dio_rdata_l_2x[25]~q ),
	.dio_rdata_l_2x_26(\dpio|dio_rdata_l_2x[26]~q ),
	.dio_rdata_l_2x_27(\dpio|dio_rdata_l_2x[27]~q ),
	.dio_rdata_l_2x_28(\dpio|dio_rdata_l_2x[28]~q ),
	.dio_rdata_l_2x_29(\dpio|dio_rdata_l_2x[29]~q ),
	.dio_rdata_l_2x_30(\dpio|dio_rdata_l_2x[30]~q ),
	.dio_rdata_l_2x_31(\dpio|dio_rdata_l_2x[31]~q ),
	.bidir_dq_0_oe_ff_inst(bidir_dq_0_oe_ff_inst),
	.bidir_dq_1_oe_ff_inst(bidir_dq_1_oe_ff_inst),
	.bidir_dq_2_oe_ff_inst(bidir_dq_2_oe_ff_inst),
	.bidir_dq_3_oe_ff_inst(bidir_dq_3_oe_ff_inst),
	.bidir_dq_4_oe_ff_inst(bidir_dq_4_oe_ff_inst),
	.bidir_dq_5_oe_ff_inst(bidir_dq_5_oe_ff_inst),
	.bidir_dq_6_oe_ff_inst(bidir_dq_6_oe_ff_inst),
	.bidir_dq_7_oe_ff_inst(bidir_dq_7_oe_ff_inst),
	.bidir_dq_0_oe_ff_inst1(bidir_dq_0_oe_ff_inst1),
	.bidir_dq_1_oe_ff_inst1(bidir_dq_1_oe_ff_inst1),
	.bidir_dq_2_oe_ff_inst1(bidir_dq_2_oe_ff_inst1),
	.bidir_dq_3_oe_ff_inst1(bidir_dq_3_oe_ff_inst1),
	.bidir_dq_4_oe_ff_inst1(bidir_dq_4_oe_ff_inst1),
	.bidir_dq_5_oe_ff_inst1(bidir_dq_5_oe_ff_inst1),
	.bidir_dq_6_oe_ff_inst1(bidir_dq_6_oe_ff_inst1),
	.bidir_dq_7_oe_ff_inst1(bidir_dq_7_oe_ff_inst1),
	.bidir_dq_0_oe_ff_inst2(bidir_dq_0_oe_ff_inst2),
	.bidir_dq_1_oe_ff_inst2(bidir_dq_1_oe_ff_inst2),
	.bidir_dq_2_oe_ff_inst2(bidir_dq_2_oe_ff_inst2),
	.bidir_dq_3_oe_ff_inst2(bidir_dq_3_oe_ff_inst2),
	.bidir_dq_4_oe_ff_inst2(bidir_dq_4_oe_ff_inst2),
	.bidir_dq_5_oe_ff_inst2(bidir_dq_5_oe_ff_inst2),
	.bidir_dq_6_oe_ff_inst2(bidir_dq_6_oe_ff_inst2),
	.bidir_dq_7_oe_ff_inst2(bidir_dq_7_oe_ff_inst2),
	.bidir_dq_0_oe_ff_inst3(bidir_dq_0_oe_ff_inst3),
	.bidir_dq_1_oe_ff_inst3(bidir_dq_1_oe_ff_inst3),
	.bidir_dq_2_oe_ff_inst3(bidir_dq_2_oe_ff_inst3),
	.bidir_dq_3_oe_ff_inst3(bidir_dq_3_oe_ff_inst3),
	.bidir_dq_4_oe_ff_inst3(bidir_dq_4_oe_ff_inst3),
	.bidir_dq_5_oe_ff_inst3(bidir_dq_5_oe_ff_inst3),
	.bidir_dq_6_oe_ff_inst3(bidir_dq_6_oe_ff_inst3),
	.bidir_dq_7_oe_ff_inst3(bidir_dq_7_oe_ff_inst3),
	.dqs_0_oe_ff_inst(dqs_0_oe_ff_inst),
	.dqs_0_oe_ff_inst1(dqs_0_oe_ff_inst1),
	.dqs_0_oe_ff_inst2(dqs_0_oe_ff_inst2),
	.dqs_0_oe_ff_inst3(dqs_0_oe_ff_inst3),
	.dqsn_0_oe_ff_inst(dqsn_0_oe_ff_inst),
	.dqsn_0_oe_ff_inst1(dqsn_0_oe_ff_inst1),
	.dqsn_0_oe_ff_inst2(dqsn_0_oe_ff_inst2),
	.dqsn_0_oe_ff_inst3(dqsn_0_oe_ff_inst3),
	.ams_pipe_3(\clk|write_clk_pipe|ams_pipe[3]~q ),
	.dqs_burst_2x_r3_0(\half_rate_wdp_gen.wdp|dqs_burst_2x_r3[0]~q ),
	.dqs_burst_2x_r3_1(\half_rate_wdp_gen.wdp|dqs_burst_2x_r3[1]~q ),
	.dqs_burst_2x_r3_2(\half_rate_wdp_gen.wdp|dqs_burst_2x_r3[2]~q ),
	.dqs_burst_2x_r3_3(\half_rate_wdp_gen.wdp|dqs_burst_2x_r3[3]~q ),
	.postamble_en_pos_2x_0(\poa|postamble_en_pos_2x[0]~q ),
	.postamble_en_pos_2x_1(\poa|postamble_en_pos_2x[1]~q ),
	.postamble_en_pos_2x_2(\poa|postamble_en_pos_2x[2]~q ),
	.postamble_en_pos_2x_3(\poa|postamble_en_pos_2x[3]~q ));

ddr3_int_ddr3_int_phy_alt_mem_phy_read_dp rdp(
	.q_b_0(q_b_0),
	.q_b_64(q_b_64),
	.q_b_1(q_b_1),
	.q_b_65(q_b_65),
	.q_b_2(q_b_2),
	.q_b_66(q_b_66),
	.q_b_3(q_b_3),
	.q_b_67(q_b_67),
	.q_b_4(q_b_4),
	.q_b_68(q_b_68),
	.q_b_5(q_b_5),
	.q_b_69(q_b_69),
	.q_b_6(q_b_6),
	.q_b_70(q_b_70),
	.q_b_7(q_b_7),
	.q_b_71(q_b_71),
	.q_b_16(q_b_16),
	.q_b_80(q_b_80),
	.q_b_17(q_b_17),
	.q_b_81(q_b_81),
	.q_b_18(q_b_18),
	.q_b_82(q_b_82),
	.q_b_19(q_b_19),
	.q_b_83(q_b_83),
	.q_b_20(q_b_20),
	.q_b_84(q_b_84),
	.q_b_21(q_b_21),
	.q_b_85(q_b_85),
	.q_b_22(q_b_22),
	.q_b_86(q_b_86),
	.q_b_23(q_b_23),
	.q_b_87(q_b_87),
	.q_b_32(q_b_32),
	.q_b_96(q_b_96),
	.q_b_33(q_b_33),
	.q_b_97(q_b_97),
	.q_b_34(q_b_34),
	.q_b_98(q_b_98),
	.q_b_35(q_b_35),
	.q_b_99(q_b_99),
	.q_b_36(q_b_36),
	.q_b_100(q_b_100),
	.q_b_37(q_b_37),
	.q_b_101(q_b_101),
	.q_b_38(q_b_38),
	.q_b_102(q_b_102),
	.q_b_39(q_b_39),
	.q_b_103(q_b_103),
	.q_b_48(q_b_48),
	.q_b_112(q_b_112),
	.q_b_49(q_b_49),
	.q_b_113(q_b_113),
	.q_b_50(q_b_50),
	.q_b_114(q_b_114),
	.q_b_51(q_b_51),
	.q_b_115(q_b_115),
	.q_b_52(q_b_52),
	.q_b_116(q_b_116),
	.q_b_53(q_b_53),
	.q_b_117(q_b_117),
	.q_b_54(q_b_54),
	.q_b_118(q_b_118),
	.q_b_55(q_b_55),
	.q_b_119(q_b_119),
	.q_b_8(q_b_8),
	.q_b_72(q_b_72),
	.q_b_9(q_b_9),
	.q_b_73(q_b_73),
	.q_b_10(q_b_10),
	.q_b_74(q_b_74),
	.q_b_11(q_b_11),
	.q_b_75(q_b_75),
	.q_b_12(q_b_12),
	.q_b_76(q_b_76),
	.q_b_13(q_b_13),
	.q_b_77(q_b_77),
	.q_b_14(q_b_14),
	.q_b_78(q_b_78),
	.q_b_15(q_b_15),
	.q_b_79(q_b_79),
	.q_b_24(q_b_24),
	.q_b_88(q_b_88),
	.q_b_25(q_b_25),
	.q_b_89(q_b_89),
	.q_b_26(q_b_26),
	.q_b_90(q_b_90),
	.q_b_27(q_b_27),
	.q_b_91(q_b_91),
	.q_b_28(q_b_28),
	.q_b_92(q_b_92),
	.q_b_29(q_b_29),
	.q_b_93(q_b_93),
	.q_b_30(q_b_30),
	.q_b_94(q_b_94),
	.q_b_31(q_b_31),
	.q_b_95(q_b_95),
	.q_b_40(q_b_40),
	.q_b_104(q_b_104),
	.q_b_41(q_b_41),
	.q_b_105(q_b_105),
	.q_b_42(q_b_42),
	.q_b_106(q_b_106),
	.q_b_43(q_b_43),
	.q_b_107(q_b_107),
	.q_b_44(q_b_44),
	.q_b_108(q_b_108),
	.q_b_45(q_b_45),
	.q_b_109(q_b_109),
	.q_b_46(q_b_46),
	.q_b_110(q_b_110),
	.q_b_47(q_b_47),
	.q_b_111(q_b_111),
	.q_b_56(q_b_56),
	.q_b_120(q_b_120),
	.q_b_57(q_b_57),
	.q_b_121(q_b_121),
	.q_b_58(q_b_58),
	.q_b_122(q_b_122),
	.q_b_59(q_b_59),
	.q_b_123(q_b_123),
	.q_b_60(q_b_60),
	.q_b_124(q_b_124),
	.q_b_61(q_b_61),
	.q_b_125(q_b_125),
	.q_b_62(q_b_62),
	.q_b_126(q_b_126),
	.q_b_63(q_b_63),
	.q_b_127(q_b_127),
	.clk_0(clk_0),
	.clk_4(\clk|half_rate.pll|altpll_component|auto_generated|clk[4] ),
	.dio_rdata_h_2x_0(\dpio|dio_rdata_h_2x[0]~q ),
	.rd_addr_2x_0(\poa|rd_addr_2x[0]~q ),
	.rd_addr_0(\rdv_pipe|rd_addr[0]~q ),
	.dio_rdata_h_2x_1(\dpio|dio_rdata_h_2x[1]~q ),
	.dio_rdata_h_2x_2(\dpio|dio_rdata_h_2x[2]~q ),
	.dio_rdata_h_2x_3(\dpio|dio_rdata_h_2x[3]~q ),
	.dio_rdata_h_2x_4(\dpio|dio_rdata_h_2x[4]~q ),
	.dio_rdata_h_2x_5(\dpio|dio_rdata_h_2x[5]~q ),
	.dio_rdata_h_2x_6(\dpio|dio_rdata_h_2x[6]~q ),
	.dio_rdata_h_2x_7(\dpio|dio_rdata_h_2x[7]~q ),
	.dio_rdata_h_2x_8(\dpio|dio_rdata_h_2x[8]~q ),
	.dio_rdata_h_2x_9(\dpio|dio_rdata_h_2x[9]~q ),
	.dio_rdata_h_2x_10(\dpio|dio_rdata_h_2x[10]~q ),
	.dio_rdata_h_2x_11(\dpio|dio_rdata_h_2x[11]~q ),
	.dio_rdata_h_2x_12(\dpio|dio_rdata_h_2x[12]~q ),
	.dio_rdata_h_2x_13(\dpio|dio_rdata_h_2x[13]~q ),
	.dio_rdata_h_2x_14(\dpio|dio_rdata_h_2x[14]~q ),
	.dio_rdata_h_2x_15(\dpio|dio_rdata_h_2x[15]~q ),
	.dio_rdata_h_2x_16(\dpio|dio_rdata_h_2x[16]~q ),
	.dio_rdata_h_2x_17(\dpio|dio_rdata_h_2x[17]~q ),
	.dio_rdata_h_2x_18(\dpio|dio_rdata_h_2x[18]~q ),
	.dio_rdata_h_2x_19(\dpio|dio_rdata_h_2x[19]~q ),
	.dio_rdata_h_2x_20(\dpio|dio_rdata_h_2x[20]~q ),
	.dio_rdata_h_2x_21(\dpio|dio_rdata_h_2x[21]~q ),
	.dio_rdata_h_2x_22(\dpio|dio_rdata_h_2x[22]~q ),
	.dio_rdata_h_2x_23(\dpio|dio_rdata_h_2x[23]~q ),
	.dio_rdata_h_2x_24(\dpio|dio_rdata_h_2x[24]~q ),
	.dio_rdata_h_2x_25(\dpio|dio_rdata_h_2x[25]~q ),
	.dio_rdata_h_2x_26(\dpio|dio_rdata_h_2x[26]~q ),
	.dio_rdata_h_2x_27(\dpio|dio_rdata_h_2x[27]~q ),
	.dio_rdata_h_2x_28(\dpio|dio_rdata_h_2x[28]~q ),
	.dio_rdata_h_2x_29(\dpio|dio_rdata_h_2x[29]~q ),
	.dio_rdata_h_2x_30(\dpio|dio_rdata_h_2x[30]~q ),
	.dio_rdata_h_2x_31(\dpio|dio_rdata_h_2x[31]~q ),
	.dio_rdata_l_2x_0(\dpio|dio_rdata_l_2x[0]~q ),
	.dio_rdata_l_2x_1(\dpio|dio_rdata_l_2x[1]~q ),
	.dio_rdata_l_2x_2(\dpio|dio_rdata_l_2x[2]~q ),
	.dio_rdata_l_2x_3(\dpio|dio_rdata_l_2x[3]~q ),
	.dio_rdata_l_2x_4(\dpio|dio_rdata_l_2x[4]~q ),
	.dio_rdata_l_2x_5(\dpio|dio_rdata_l_2x[5]~q ),
	.dio_rdata_l_2x_6(\dpio|dio_rdata_l_2x[6]~q ),
	.dio_rdata_l_2x_7(\dpio|dio_rdata_l_2x[7]~q ),
	.dio_rdata_l_2x_8(\dpio|dio_rdata_l_2x[8]~q ),
	.dio_rdata_l_2x_9(\dpio|dio_rdata_l_2x[9]~q ),
	.dio_rdata_l_2x_10(\dpio|dio_rdata_l_2x[10]~q ),
	.dio_rdata_l_2x_11(\dpio|dio_rdata_l_2x[11]~q ),
	.dio_rdata_l_2x_12(\dpio|dio_rdata_l_2x[12]~q ),
	.dio_rdata_l_2x_13(\dpio|dio_rdata_l_2x[13]~q ),
	.dio_rdata_l_2x_14(\dpio|dio_rdata_l_2x[14]~q ),
	.dio_rdata_l_2x_15(\dpio|dio_rdata_l_2x[15]~q ),
	.dio_rdata_l_2x_16(\dpio|dio_rdata_l_2x[16]~q ),
	.dio_rdata_l_2x_17(\dpio|dio_rdata_l_2x[17]~q ),
	.dio_rdata_l_2x_18(\dpio|dio_rdata_l_2x[18]~q ),
	.dio_rdata_l_2x_19(\dpio|dio_rdata_l_2x[19]~q ),
	.dio_rdata_l_2x_20(\dpio|dio_rdata_l_2x[20]~q ),
	.dio_rdata_l_2x_21(\dpio|dio_rdata_l_2x[21]~q ),
	.dio_rdata_l_2x_22(\dpio|dio_rdata_l_2x[22]~q ),
	.dio_rdata_l_2x_23(\dpio|dio_rdata_l_2x[23]~q ),
	.dio_rdata_l_2x_24(\dpio|dio_rdata_l_2x[24]~q ),
	.dio_rdata_l_2x_25(\dpio|dio_rdata_l_2x[25]~q ),
	.dio_rdata_l_2x_26(\dpio|dio_rdata_l_2x[26]~q ),
	.dio_rdata_l_2x_27(\dpio|dio_rdata_l_2x[27]~q ),
	.dio_rdata_l_2x_28(\dpio|dio_rdata_l_2x[28]~q ),
	.dio_rdata_l_2x_29(\dpio|dio_rdata_l_2x[29]~q ),
	.dio_rdata_l_2x_30(\dpio|dio_rdata_l_2x[30]~q ),
	.dio_rdata_l_2x_31(\dpio|dio_rdata_l_2x[31]~q ),
	.reset_phy_clk_1x_n(\clk|reset_rdp_phy_clk_pipe|ams_pipe[1]~q ),
	.reset_resync_clk_2x_n(\clk|resync_clk_2x_pipe|ams_pipe[1]~q ));

arriaii_lcell_comb \merged_doing_rd[4] (
	.dataa(!ctl_init_success),
	.datab(!do_read_r),
	.datac(!rdwr_data_valid_r),
	.datad(!doing_read),
	.datae(!\seq_wrapper|seq_inst|seq_rdv_doing_rd[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\merged_doing_rd[4]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \merged_doing_rd[4] .extended_lut = "off";
defparam \merged_doing_rd[4] .lut_mask = 64'h0105FFFF0105FFFF;
defparam \merged_doing_rd[4] .shared_arith = "off";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_addr_cmd (
	clk_0,
	clk_3,
	dataout_0,
	dataout_01,
	dataout_02,
	dataout_03,
	dataout_04,
	dataout_05,
	dataout_06,
	dataout_07,
	dataout_08,
	dataout_09,
	dataout_010,
	dataout_011,
	dataout_012,
	dataout_013,
	dataout_014,
	dataout_015,
	dataout_016,
	dataout_017,
	dataout_018,
	dataout_019,
	dataout_020,
	dataout_021,
	dataout_022,
	dataout_023,
	seq_ac_cke_1,
	seq_ac_addr_0,
	seq_ac_addr_14,
	seq_ac_addr_1,
	seq_ac_addr_15,
	seq_ac_addr_16,
	seq_ac_addr_17,
	seq_ac_addr_18,
	seq_ac_addr_5,
	seq_ac_addr_19,
	seq_ac_addr_8,
	seq_ac_addr_22,
	seq_ac_addr_10,
	seq_ac_addr_24,
	seq_ac_addr_12,
	seq_ac_addr_26,
	seq_ac_ba_0,
	seq_ac_ba_3,
	seq_ac_ba_1,
	seq_ac_ba_4,
	seq_ac_rst_n_0,
	ams_pipe_1,
	seq_ac_add_1t_ac_lat_internal,
	seq_ac_cs_n_0,
	seq_ac_sel,
	afi_cs_n_1,
	int_cke_r_0,
	afi_addr_0,
	afi_addr_1,
	afi_addr_2,
	afi_addr_3,
	afi_addr_4,
	afi_addr_5,
	afi_addr_6,
	afi_addr_7,
	afi_addr_8,
	afi_addr_9,
	afi_addr_10,
	afi_addr_11,
	afi_addr_12,
	afi_addr_13,
	afi_ba_0,
	afi_ba_1,
	afi_ba_2,
	afi_ras_n_0,
	afi_cas_n_0,
	afi_we_n_0,
	GND_port,
	seq_ac_cas_n_0,
	seq_ac_cas_n_1,
	seq_ac_cs_n_1,
	seq_ac_ras_n_0,
	seq_ac_ras_n_1,
	seq_ac_we_n_0,
	seq_ac_we_n_1)/* synthesis synthesis_greybox=0 */;
input 	clk_0;
input 	clk_3;
output 	dataout_0;
output 	dataout_01;
output 	dataout_02;
output 	dataout_03;
output 	dataout_04;
output 	dataout_05;
output 	dataout_06;
output 	dataout_07;
output 	dataout_08;
output 	dataout_09;
output 	dataout_010;
output 	dataout_011;
output 	dataout_012;
output 	dataout_013;
output 	dataout_014;
output 	dataout_015;
output 	dataout_016;
output 	dataout_017;
output 	dataout_018;
output 	dataout_019;
output 	dataout_020;
output 	dataout_021;
output 	dataout_022;
output 	dataout_023;
input 	seq_ac_cke_1;
input 	seq_ac_addr_0;
input 	seq_ac_addr_14;
input 	seq_ac_addr_1;
input 	seq_ac_addr_15;
input 	seq_ac_addr_16;
input 	seq_ac_addr_17;
input 	seq_ac_addr_18;
input 	seq_ac_addr_5;
input 	seq_ac_addr_19;
input 	seq_ac_addr_8;
input 	seq_ac_addr_22;
input 	seq_ac_addr_10;
input 	seq_ac_addr_24;
input 	seq_ac_addr_12;
input 	seq_ac_addr_26;
input 	seq_ac_ba_0;
input 	seq_ac_ba_3;
input 	seq_ac_ba_1;
input 	seq_ac_ba_4;
input 	seq_ac_rst_n_0;
input 	ams_pipe_1;
input 	seq_ac_add_1t_ac_lat_internal;
input 	seq_ac_cs_n_0;
input 	seq_ac_sel;
input 	afi_cs_n_1;
input 	int_cke_r_0;
input 	afi_addr_0;
input 	afi_addr_1;
input 	afi_addr_2;
input 	afi_addr_3;
input 	afi_addr_4;
input 	afi_addr_5;
input 	afi_addr_6;
input 	afi_addr_7;
input 	afi_addr_8;
input 	afi_addr_9;
input 	afi_addr_10;
input 	afi_addr_11;
input 	afi_addr_12;
input 	afi_addr_13;
input 	afi_ba_0;
input 	afi_ba_1;
input 	afi_ba_2;
input 	afi_ras_n_0;
input 	afi_cas_n_0;
input 	afi_we_n_0;
input 	GND_port;
input 	seq_ac_cas_n_0;
input 	seq_ac_cas_n_1;
input 	seq_ac_cs_n_1;
input 	seq_ac_ras_n_0;
input 	seq_ac_ras_n_1;
input 	seq_ac_we_n_0;
input 	seq_ac_we_n_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \period_sel_addr[7]~q ;
wire \count_addr_2x[7]~q ;
wire \count_addr_rst_n_2x_r~q ;
wire \period_sel_addr~0_combout ;
wire \count_addr[0]~q ;
wire \count_addr[0]~0_combout ;


ddr3_int_ddr3_int_phy_alt_mem_phy_ac_2 \addr[11].addr_struct (
	.phy_clk_1x(clk_0),
	.clk_3(clk_3),
	.dataout_0(dataout_014),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.period_sel_addr_7(\period_sel_addr[7]~q ),
	.seq_ac_sel(seq_ac_sel),
	.afi_addr_11(afi_addr_11),
	.GND_port(GND_port));

ddr3_int_ddr3_int_phy_alt_mem_phy_ac_3 \addr[12].addr_struct (
	.phy_clk_1x(clk_0),
	.clk_3(clk_3),
	.dataout_0(dataout_015),
	.seq_ac_addr_12(seq_ac_addr_12),
	.seq_ac_addr_26(seq_ac_addr_26),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.period_sel_addr_7(\period_sel_addr[7]~q ),
	.seq_ac_sel(seq_ac_sel),
	.afi_addr_12(afi_addr_12));

ddr3_int_ddr3_int_phy_alt_mem_phy_ac_4 \addr[13].addr_struct (
	.phy_clk_1x(clk_0),
	.clk_3(clk_3),
	.dataout_0(dataout_016),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.period_sel_addr_7(\period_sel_addr[7]~q ),
	.seq_ac_sel(seq_ac_sel),
	.afi_addr_13(afi_addr_13),
	.GND_port(GND_port));

ddr3_int_ddr3_int_phy_alt_mem_phy_ac_14 \ba[0].ba_struct (
	.phy_clk_1x(clk_0),
	.clk_3(clk_3),
	.dataout_0(dataout_017),
	.seq_ac_ba_0(seq_ac_ba_0),
	.seq_ac_ba_3(seq_ac_ba_3),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.period_sel_addr_7(\period_sel_addr[7]~q ),
	.seq_ac_sel(seq_ac_sel),
	.afi_ba_0(afi_ba_0));

ddr3_int_ddr3_int_phy_alt_mem_phy_ac_15 \ba[1].ba_struct (
	.phy_clk_1x(clk_0),
	.clk_3(clk_3),
	.dataout_0(dataout_018),
	.seq_ac_ba_1(seq_ac_ba_1),
	.seq_ac_ba_4(seq_ac_ba_4),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.period_sel_addr_7(\period_sel_addr[7]~q ),
	.seq_ac_sel(seq_ac_sel),
	.afi_ba_1(afi_ba_1));

ddr3_int_ddr3_int_phy_alt_mem_phy_ac_16 \ba[2].ba_struct (
	.phy_clk_1x(clk_0),
	.clk_3(clk_3),
	.dataout_0(dataout_019),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.period_sel_addr_7(\period_sel_addr[7]~q ),
	.seq_ac_sel(seq_ac_sel),
	.afi_ba_2(afi_ba_2),
	.GND_port(GND_port));

ddr3_int_ddr3_int_phy_alt_mem_phy_ac_17 cas_n_struct(
	.phy_clk_1x(clk_0),
	.clk_3(clk_3),
	.dataout_0(dataout_021),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.period_sel_addr_7(\period_sel_addr[7]~q ),
	.seq_ac_sel(seq_ac_sel),
	.afi_cas_n_0(afi_cas_n_0),
	.seq_ac_cas_n_0(seq_ac_cas_n_0),
	.seq_ac_cas_n_1(seq_ac_cas_n_1));

ddr3_int_ddr3_int_phy_alt_mem_phy_ac_18 \cke[0].cke_struct (
	.phy_clk_1x(clk_0),
	.clk_3(clk_3),
	.dataout_0(dataout_02),
	.seq_ac_cke_1(seq_ac_cke_1),
	.ams_pipe_1(ams_pipe_1),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.period_sel_addr_7(\period_sel_addr[7]~q ),
	.seq_ac_sel(seq_ac_sel),
	.int_cke_r_0(int_cke_r_0));

ddr3_int_ddr3_int_phy_alt_mem_phy_ac_19 \cs_n[0].cs_n_struct (
	.phy_clk_1x(clk_0),
	.clk_3(clk_3),
	.dataout_0(dataout_01),
	.ams_pipe_1(ams_pipe_1),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.period_sel_addr_7(\period_sel_addr[7]~q ),
	.seq_ac_cs_n_0(seq_ac_cs_n_0),
	.seq_ac_sel(seq_ac_sel),
	.afi_cs_n_1(afi_cs_n_1),
	.seq_ac_cs_n_1(seq_ac_cs_n_1));

ddr3_int_ddr3_int_phy_alt_mem_phy_ac_21 \gen_odt.odt[0].odt_struct (
	.phy_clk_1x(clk_0),
	.clk_3(clk_3),
	.dataout_0(dataout_0),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.period_sel_addr_7(\period_sel_addr[7]~q ));

ddr3_int_ddr3_int_phy_alt_mem_phy_ac_22 ras_n_struct(
	.phy_clk_1x(clk_0),
	.clk_3(clk_3),
	.dataout_0(dataout_020),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.period_sel_addr_7(\period_sel_addr[7]~q ),
	.seq_ac_sel(seq_ac_sel),
	.afi_ras_n_0(afi_ras_n_0),
	.seq_ac_ras_n_0(seq_ac_ras_n_0),
	.seq_ac_ras_n_1(seq_ac_ras_n_1));

ddr3_int_ddr3_int_phy_alt_mem_phy_ac_23 we_n_struct(
	.phy_clk_1x(clk_0),
	.clk_3(clk_3),
	.dataout_0(dataout_022),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.period_sel_addr_7(\period_sel_addr[7]~q ),
	.seq_ac_sel(seq_ac_sel),
	.afi_we_n_0(afi_we_n_0),
	.seq_ac_we_n_0(seq_ac_we_n_0),
	.seq_ac_we_n_1(seq_ac_we_n_1));

ddr3_int_ddr3_int_phy_alt_mem_phy_ac_20 \ddr3_rst.ddr3_rst_struct (
	.phy_clk_1x(clk_0),
	.clk_3(clk_3),
	.dataout_0(dataout_023),
	.seq_ac_rst_n_0(seq_ac_rst_n_0),
	.ams_pipe_1(ams_pipe_1),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.period_sel_addr_7(\period_sel_addr[7]~q ),
	.seq_ac_sel(seq_ac_sel));

ddr3_int_ddr3_int_phy_alt_mem_phy_ac \addr[0].addr_struct (
	.phy_clk_1x(clk_0),
	.clk_3(clk_3),
	.dataout_0(dataout_03),
	.seq_ac_addr_0(seq_ac_addr_0),
	.seq_ac_addr_14(seq_ac_addr_14),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.period_sel_addr_7(\period_sel_addr[7]~q ),
	.seq_ac_sel(seq_ac_sel),
	.afi_addr_0(afi_addr_0));

ddr3_int_ddr3_int_phy_alt_mem_phy_ac_5 \addr[1].addr_struct (
	.phy_clk_1x(clk_0),
	.clk_3(clk_3),
	.dataout_0(dataout_04),
	.seq_ac_addr_1(seq_ac_addr_1),
	.seq_ac_addr_15(seq_ac_addr_15),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.period_sel_addr_7(\period_sel_addr[7]~q ),
	.seq_ac_sel(seq_ac_sel),
	.afi_addr_1(afi_addr_1));

ddr3_int_ddr3_int_phy_alt_mem_phy_ac_6 \addr[2].addr_struct (
	.phy_clk_1x(clk_0),
	.clk_3(clk_3),
	.dataout_0(dataout_05),
	.seq_ac_addr_16(seq_ac_addr_16),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.period_sel_addr_7(\period_sel_addr[7]~q ),
	.seq_ac_sel(seq_ac_sel),
	.afi_addr_2(afi_addr_2));

ddr3_int_ddr3_int_phy_alt_mem_phy_ac_7 \addr[3].addr_struct (
	.phy_clk_1x(clk_0),
	.clk_3(clk_3),
	.dataout_0(dataout_06),
	.seq_ac_addr_17(seq_ac_addr_17),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.period_sel_addr_7(\period_sel_addr[7]~q ),
	.seq_ac_sel(seq_ac_sel),
	.afi_addr_3(afi_addr_3));

ddr3_int_ddr3_int_phy_alt_mem_phy_ac_8 \addr[4].addr_struct (
	.phy_clk_1x(clk_0),
	.clk_3(clk_3),
	.dataout_0(dataout_07),
	.seq_ac_addr_18(seq_ac_addr_18),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.period_sel_addr_7(\period_sel_addr[7]~q ),
	.seq_ac_sel(seq_ac_sel),
	.afi_addr_4(afi_addr_4));

ddr3_int_ddr3_int_phy_alt_mem_phy_ac_9 \addr[5].addr_struct (
	.phy_clk_1x(clk_0),
	.clk_3(clk_3),
	.dataout_0(dataout_08),
	.seq_ac_addr_5(seq_ac_addr_5),
	.seq_ac_addr_19(seq_ac_addr_19),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.period_sel_addr_7(\period_sel_addr[7]~q ),
	.seq_ac_sel(seq_ac_sel),
	.afi_addr_5(afi_addr_5));

ddr3_int_ddr3_int_phy_alt_mem_phy_ac_10 \addr[6].addr_struct (
	.phy_clk_1x(clk_0),
	.clk_3(clk_3),
	.dataout_0(dataout_09),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.period_sel_addr_7(\period_sel_addr[7]~q ),
	.seq_ac_sel(seq_ac_sel),
	.afi_addr_6(afi_addr_6),
	.GND_port(GND_port));

ddr3_int_ddr3_int_phy_alt_mem_phy_ac_11 \addr[7].addr_struct (
	.phy_clk_1x(clk_0),
	.clk_3(clk_3),
	.dataout_0(dataout_010),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.period_sel_addr_7(\period_sel_addr[7]~q ),
	.seq_ac_sel(seq_ac_sel),
	.afi_addr_7(afi_addr_7),
	.GND_port(GND_port));

ddr3_int_ddr3_int_phy_alt_mem_phy_ac_12 \addr[8].addr_struct (
	.phy_clk_1x(clk_0),
	.clk_3(clk_3),
	.dataout_0(dataout_011),
	.seq_ac_addr_8(seq_ac_addr_8),
	.seq_ac_addr_22(seq_ac_addr_22),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.period_sel_addr_7(\period_sel_addr[7]~q ),
	.seq_ac_sel(seq_ac_sel),
	.afi_addr_8(afi_addr_8));

ddr3_int_ddr3_int_phy_alt_mem_phy_ac_13 \addr[9].addr_struct (
	.phy_clk_1x(clk_0),
	.clk_3(clk_3),
	.dataout_0(dataout_012),
	.seq_ac_addr_0(seq_ac_addr_0),
	.seq_ac_addr_14(seq_ac_addr_14),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.period_sel_addr_7(\period_sel_addr[7]~q ),
	.seq_ac_sel(seq_ac_sel),
	.afi_addr_9(afi_addr_9));

ddr3_int_ddr3_int_phy_alt_mem_phy_ac_1 \addr[10].addr_struct (
	.phy_clk_1x(clk_0),
	.clk_3(clk_3),
	.dataout_0(dataout_013),
	.seq_ac_addr_10(seq_ac_addr_10),
	.seq_ac_addr_24(seq_ac_addr_24),
	.seq_ac_add_1t_ac_lat_internal(seq_ac_add_1t_ac_lat_internal),
	.period_sel_addr_7(\period_sel_addr[7]~q ),
	.seq_ac_sel(seq_ac_sel),
	.afi_addr_10(afi_addr_10));

dffeas \period_sel_addr[7] (
	.clk(clk_3),
	.d(\period_sel_addr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\period_sel_addr[7]~q ),
	.prn(vcc));
defparam \period_sel_addr[7] .is_wysiwyg = "true";
defparam \period_sel_addr[7] .power_up = "low";

dffeas \count_addr_2x[7] (
	.clk(clk_3),
	.d(\count_addr[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\count_addr_2x[7]~q ),
	.prn(vcc));
defparam \count_addr_2x[7] .is_wysiwyg = "true";
defparam \count_addr_2x[7] .power_up = "low";

dffeas count_addr_rst_n_2x_r(
	.clk(clk_3),
	.d(\count_addr_2x[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\count_addr_rst_n_2x_r~q ),
	.prn(vcc));
defparam count_addr_rst_n_2x_r.is_wysiwyg = "true";
defparam count_addr_rst_n_2x_r.power_up = "low";

arriaii_lcell_comb \period_sel_addr~0 (
	.dataa(!\count_addr_2x[7]~q ),
	.datab(!\count_addr_rst_n_2x_r~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\period_sel_addr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \period_sel_addr~0 .extended_lut = "off";
defparam \period_sel_addr~0 .lut_mask = 64'h9999999999999999;
defparam \period_sel_addr~0 .shared_arith = "off";

dffeas \count_addr[0] (
	.clk(clk_0),
	.d(\count_addr[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\count_addr[0]~q ),
	.prn(vcc));
defparam \count_addr[0] .is_wysiwyg = "true";
defparam \count_addr[0] .power_up = "low";

arriaii_lcell_comb \count_addr[0]~0 (
	.dataa(!\count_addr[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count_addr[0]~0 .extended_lut = "off";
defparam \count_addr[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \count_addr[0]~0 .shared_arith = "off";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_ac (
	phy_clk_1x,
	clk_3,
	dataout_0,
	seq_ac_addr_0,
	seq_ac_addr_14,
	seq_ac_add_1t_ac_lat_internal,
	period_sel_addr_7,
	seq_ac_sel,
	afi_addr_0)/* synthesis synthesis_greybox=0 */;
input 	phy_clk_1x;
input 	clk_3;
output 	dataout_0;
input 	seq_ac_addr_0;
input 	seq_ac_addr_14;
input 	seq_ac_add_1t_ac_lat_internal;
input 	period_sel_addr_7;
input 	seq_ac_sel;
input 	afi_addr_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ac_h~q ;
wire \ac_l~q ;
wire \ac_2x_r~q ;
wire \ac_2x_2r~q ;
wire \ac_h_2r~q ;
wire \ac_l_2r~q ;
wire \ac_2x~0_combout ;
wire \ac_1t~q ;
wire \ac_2x_r~0_combout ;
wire \ac_h_r~q ;
wire \ac_l_r~q ;
wire \ac_h_r~0_combout ;
wire \ac_l_r~0_combout ;


ddr3_int_altddio_out_1 \half_rate.addr_pin (
	.outclock(clk_3),
	.dataout({dataout_0}),
	.datain_l({\ac_2x_r~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_h(
	.clk(phy_clk_1x),
	.d(seq_ac_addr_0),
	.asdata(afi_addr_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_h~q ),
	.prn(vcc));
defparam ac_h.is_wysiwyg = "true";
defparam ac_h.power_up = "low";

dffeas ac_l(
	.clk(phy_clk_1x),
	.d(seq_ac_addr_14),
	.asdata(afi_addr_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_l~q ),
	.prn(vcc));
defparam ac_l.is_wysiwyg = "true";
defparam ac_l.power_up = "low";

dffeas ac_2x_r(
	.clk(clk_3),
	.d(\ac_2x_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_r~q ),
	.prn(vcc));
defparam ac_2x_r.is_wysiwyg = "true";
defparam ac_2x_r.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_3),
	.d(\ac_2x_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

dffeas ac_h_2r(
	.clk(clk_3),
	.d(\ac_h_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_2r~q ),
	.prn(vcc));
defparam ac_h_2r.is_wysiwyg = "true";
defparam ac_h_2r.power_up = "low";

dffeas ac_l_2r(
	.clk(clk_3),
	.d(\ac_l_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_2r~q ),
	.prn(vcc));
defparam ac_l_2r.is_wysiwyg = "true";
defparam ac_l_2r.power_up = "low";

arriaii_lcell_comb \ac_2x~0 (
	.dataa(!period_sel_addr_7),
	.datab(!\ac_h_2r~q ),
	.datac(!\ac_l_2r~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x~0 .extended_lut = "off";
defparam \ac_2x~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \ac_2x~0 .shared_arith = "off";

dffeas ac_1t(
	.clk(clk_3),
	.d(\ac_2x~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

arriaii_lcell_comb \ac_2x_r~0 (
	.dataa(!seq_ac_add_1t_ac_lat_internal),
	.datab(!\ac_2x~0_combout ),
	.datac(!\ac_1t~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x_r~0 .extended_lut = "off";
defparam \ac_2x_r~0 .lut_mask = 64'h2727272727272727;
defparam \ac_2x_r~0 .shared_arith = "off";

dffeas ac_h_r(
	.clk(phy_clk_1x),
	.d(\ac_h_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_r~q ),
	.prn(vcc));
defparam ac_h_r.is_wysiwyg = "true";
defparam ac_h_r.power_up = "low";

dffeas ac_l_r(
	.clk(phy_clk_1x),
	.d(\ac_l_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_r~q ),
	.prn(vcc));
defparam ac_l_r.is_wysiwyg = "true";
defparam ac_l_r.power_up = "low";

arriaii_lcell_comb \ac_h_r~0 (
	.dataa(!\ac_h~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_h_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_h_r~0 .extended_lut = "off";
defparam \ac_h_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_h_r~0 .shared_arith = "off";

arriaii_lcell_comb \ac_l_r~0 (
	.dataa(!\ac_l~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_l_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_l_r~0 .extended_lut = "off";
defparam \ac_l_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_l_r~0 .shared_arith = "off";

endmodule

module ddr3_int_altddio_out_1 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
inout 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_ddio_out_6ed auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module ddr3_int_ddio_out_6ed (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



arriaii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_ac_1 (
	phy_clk_1x,
	clk_3,
	dataout_0,
	seq_ac_addr_10,
	seq_ac_addr_24,
	seq_ac_add_1t_ac_lat_internal,
	period_sel_addr_7,
	seq_ac_sel,
	afi_addr_10)/* synthesis synthesis_greybox=0 */;
input 	phy_clk_1x;
input 	clk_3;
output 	dataout_0;
input 	seq_ac_addr_10;
input 	seq_ac_addr_24;
input 	seq_ac_add_1t_ac_lat_internal;
input 	period_sel_addr_7;
input 	seq_ac_sel;
input 	afi_addr_10;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ac_h~q ;
wire \ac_l~q ;
wire \ac_2x_r~q ;
wire \ac_2x_2r~q ;
wire \ac_h_2r~q ;
wire \ac_l_2r~q ;
wire \ac_2x~0_combout ;
wire \ac_1t~q ;
wire \ac_2x_r~0_combout ;
wire \ac_h_r~q ;
wire \ac_l_r~q ;
wire \ac_h_r~0_combout ;
wire \ac_l_r~0_combout ;


ddr3_int_altddio_out_2 \half_rate.addr_pin (
	.outclock(clk_3),
	.dataout({dataout_0}),
	.datain_l({\ac_2x_r~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_h(
	.clk(phy_clk_1x),
	.d(seq_ac_addr_10),
	.asdata(afi_addr_10),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_h~q ),
	.prn(vcc));
defparam ac_h.is_wysiwyg = "true";
defparam ac_h.power_up = "low";

dffeas ac_l(
	.clk(phy_clk_1x),
	.d(seq_ac_addr_24),
	.asdata(afi_addr_10),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_l~q ),
	.prn(vcc));
defparam ac_l.is_wysiwyg = "true";
defparam ac_l.power_up = "low";

dffeas ac_2x_r(
	.clk(clk_3),
	.d(\ac_2x_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_r~q ),
	.prn(vcc));
defparam ac_2x_r.is_wysiwyg = "true";
defparam ac_2x_r.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_3),
	.d(\ac_2x_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

dffeas ac_h_2r(
	.clk(clk_3),
	.d(\ac_h_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_2r~q ),
	.prn(vcc));
defparam ac_h_2r.is_wysiwyg = "true";
defparam ac_h_2r.power_up = "low";

dffeas ac_l_2r(
	.clk(clk_3),
	.d(\ac_l_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_2r~q ),
	.prn(vcc));
defparam ac_l_2r.is_wysiwyg = "true";
defparam ac_l_2r.power_up = "low";

arriaii_lcell_comb \ac_2x~0 (
	.dataa(!period_sel_addr_7),
	.datab(!\ac_h_2r~q ),
	.datac(!\ac_l_2r~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x~0 .extended_lut = "off";
defparam \ac_2x~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \ac_2x~0 .shared_arith = "off";

dffeas ac_1t(
	.clk(clk_3),
	.d(\ac_2x~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

arriaii_lcell_comb \ac_2x_r~0 (
	.dataa(!seq_ac_add_1t_ac_lat_internal),
	.datab(!\ac_2x~0_combout ),
	.datac(!\ac_1t~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x_r~0 .extended_lut = "off";
defparam \ac_2x_r~0 .lut_mask = 64'h2727272727272727;
defparam \ac_2x_r~0 .shared_arith = "off";

dffeas ac_h_r(
	.clk(phy_clk_1x),
	.d(\ac_h_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_r~q ),
	.prn(vcc));
defparam ac_h_r.is_wysiwyg = "true";
defparam ac_h_r.power_up = "low";

dffeas ac_l_r(
	.clk(phy_clk_1x),
	.d(\ac_l_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_r~q ),
	.prn(vcc));
defparam ac_l_r.is_wysiwyg = "true";
defparam ac_l_r.power_up = "low";

arriaii_lcell_comb \ac_h_r~0 (
	.dataa(!\ac_h~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_h_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_h_r~0 .extended_lut = "off";
defparam \ac_h_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_h_r~0 .shared_arith = "off";

arriaii_lcell_comb \ac_l_r~0 (
	.dataa(!\ac_l~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_l_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_l_r~0 .extended_lut = "off";
defparam \ac_l_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_l_r~0 .shared_arith = "off";

endmodule

module ddr3_int_altddio_out_2 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
inout 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_ddio_out_6ed_1 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module ddr3_int_ddio_out_6ed_1 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



arriaii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_ac_2 (
	phy_clk_1x,
	clk_3,
	dataout_0,
	seq_ac_add_1t_ac_lat_internal,
	period_sel_addr_7,
	seq_ac_sel,
	afi_addr_11,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	phy_clk_1x;
input 	clk_3;
output 	dataout_0;
input 	seq_ac_add_1t_ac_lat_internal;
input 	period_sel_addr_7;
input 	seq_ac_sel;
input 	afi_addr_11;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ac_l~q ;
wire \ac_2x_r~q ;
wire \ac_2x_2r~q ;
wire \ac_h_2r~q ;
wire \ac_l_2r~q ;
wire \ac_2x~0_combout ;
wire \ac_1t~q ;
wire \ac_2x_r~0_combout ;
wire \ac_h_r~q ;
wire \ac_l_r~q ;
wire \ac_h_r~0_combout ;
wire \ac_l_r~0_combout ;


ddr3_int_altddio_out_3 \half_rate.addr_pin (
	.outclock(clk_3),
	.dataout({dataout_0}),
	.datain_l({\ac_2x_r~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_l(
	.clk(phy_clk_1x),
	.d(GND_port),
	.asdata(afi_addr_11),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_l~q ),
	.prn(vcc));
defparam ac_l.is_wysiwyg = "true";
defparam ac_l.power_up = "low";

dffeas ac_2x_r(
	.clk(clk_3),
	.d(\ac_2x_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_r~q ),
	.prn(vcc));
defparam ac_2x_r.is_wysiwyg = "true";
defparam ac_2x_r.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_3),
	.d(\ac_2x_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

dffeas ac_h_2r(
	.clk(clk_3),
	.d(\ac_h_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_2r~q ),
	.prn(vcc));
defparam ac_h_2r.is_wysiwyg = "true";
defparam ac_h_2r.power_up = "low";

dffeas ac_l_2r(
	.clk(clk_3),
	.d(\ac_l_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_2r~q ),
	.prn(vcc));
defparam ac_l_2r.is_wysiwyg = "true";
defparam ac_l_2r.power_up = "low";

arriaii_lcell_comb \ac_2x~0 (
	.dataa(!period_sel_addr_7),
	.datab(!\ac_h_2r~q ),
	.datac(!\ac_l_2r~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x~0 .extended_lut = "off";
defparam \ac_2x~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \ac_2x~0 .shared_arith = "off";

dffeas ac_1t(
	.clk(clk_3),
	.d(\ac_2x~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

arriaii_lcell_comb \ac_2x_r~0 (
	.dataa(!seq_ac_add_1t_ac_lat_internal),
	.datab(!\ac_2x~0_combout ),
	.datac(!\ac_1t~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x_r~0 .extended_lut = "off";
defparam \ac_2x_r~0 .lut_mask = 64'h2727272727272727;
defparam \ac_2x_r~0 .shared_arith = "off";

dffeas ac_h_r(
	.clk(phy_clk_1x),
	.d(\ac_h_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_r~q ),
	.prn(vcc));
defparam ac_h_r.is_wysiwyg = "true";
defparam ac_h_r.power_up = "low";

dffeas ac_l_r(
	.clk(phy_clk_1x),
	.d(\ac_l_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_r~q ),
	.prn(vcc));
defparam ac_l_r.is_wysiwyg = "true";
defparam ac_l_r.power_up = "low";

arriaii_lcell_comb \ac_h_r~0 (
	.dataa(!\ac_l~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_h_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_h_r~0 .extended_lut = "off";
defparam \ac_h_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_h_r~0 .shared_arith = "off";

arriaii_lcell_comb \ac_l_r~0 (
	.dataa(!\ac_l~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_l_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_l_r~0 .extended_lut = "off";
defparam \ac_l_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_l_r~0 .shared_arith = "off";

endmodule

module ddr3_int_altddio_out_3 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
inout 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_ddio_out_6ed_2 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module ddr3_int_ddio_out_6ed_2 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



arriaii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_ac_3 (
	phy_clk_1x,
	clk_3,
	dataout_0,
	seq_ac_addr_12,
	seq_ac_addr_26,
	seq_ac_add_1t_ac_lat_internal,
	period_sel_addr_7,
	seq_ac_sel,
	afi_addr_12)/* synthesis synthesis_greybox=0 */;
input 	phy_clk_1x;
input 	clk_3;
output 	dataout_0;
input 	seq_ac_addr_12;
input 	seq_ac_addr_26;
input 	seq_ac_add_1t_ac_lat_internal;
input 	period_sel_addr_7;
input 	seq_ac_sel;
input 	afi_addr_12;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ac_h~q ;
wire \ac_l~q ;
wire \ac_2x_r~q ;
wire \ac_2x_2r~q ;
wire \ac_h_2r~q ;
wire \ac_l_2r~q ;
wire \ac_2x~0_combout ;
wire \ac_1t~q ;
wire \ac_2x_r~0_combout ;
wire \ac_h_r~q ;
wire \ac_l_r~q ;
wire \ac_h_r~0_combout ;
wire \ac_l_r~0_combout ;


ddr3_int_altddio_out_4 \half_rate.addr_pin (
	.outclock(clk_3),
	.dataout({dataout_0}),
	.datain_l({\ac_2x_r~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_h(
	.clk(phy_clk_1x),
	.d(seq_ac_addr_12),
	.asdata(afi_addr_12),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_h~q ),
	.prn(vcc));
defparam ac_h.is_wysiwyg = "true";
defparam ac_h.power_up = "low";

dffeas ac_l(
	.clk(phy_clk_1x),
	.d(seq_ac_addr_26),
	.asdata(afi_addr_12),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_l~q ),
	.prn(vcc));
defparam ac_l.is_wysiwyg = "true";
defparam ac_l.power_up = "low";

dffeas ac_2x_r(
	.clk(clk_3),
	.d(\ac_2x_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_r~q ),
	.prn(vcc));
defparam ac_2x_r.is_wysiwyg = "true";
defparam ac_2x_r.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_3),
	.d(\ac_2x_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

dffeas ac_h_2r(
	.clk(clk_3),
	.d(\ac_h_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_2r~q ),
	.prn(vcc));
defparam ac_h_2r.is_wysiwyg = "true";
defparam ac_h_2r.power_up = "low";

dffeas ac_l_2r(
	.clk(clk_3),
	.d(\ac_l_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_2r~q ),
	.prn(vcc));
defparam ac_l_2r.is_wysiwyg = "true";
defparam ac_l_2r.power_up = "low";

arriaii_lcell_comb \ac_2x~0 (
	.dataa(!period_sel_addr_7),
	.datab(!\ac_h_2r~q ),
	.datac(!\ac_l_2r~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x~0 .extended_lut = "off";
defparam \ac_2x~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \ac_2x~0 .shared_arith = "off";

dffeas ac_1t(
	.clk(clk_3),
	.d(\ac_2x~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

arriaii_lcell_comb \ac_2x_r~0 (
	.dataa(!seq_ac_add_1t_ac_lat_internal),
	.datab(!\ac_2x~0_combout ),
	.datac(!\ac_1t~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x_r~0 .extended_lut = "off";
defparam \ac_2x_r~0 .lut_mask = 64'h2727272727272727;
defparam \ac_2x_r~0 .shared_arith = "off";

dffeas ac_h_r(
	.clk(phy_clk_1x),
	.d(\ac_h_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_r~q ),
	.prn(vcc));
defparam ac_h_r.is_wysiwyg = "true";
defparam ac_h_r.power_up = "low";

dffeas ac_l_r(
	.clk(phy_clk_1x),
	.d(\ac_l_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_r~q ),
	.prn(vcc));
defparam ac_l_r.is_wysiwyg = "true";
defparam ac_l_r.power_up = "low";

arriaii_lcell_comb \ac_h_r~0 (
	.dataa(!\ac_h~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_h_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_h_r~0 .extended_lut = "off";
defparam \ac_h_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_h_r~0 .shared_arith = "off";

arriaii_lcell_comb \ac_l_r~0 (
	.dataa(!\ac_l~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_l_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_l_r~0 .extended_lut = "off";
defparam \ac_l_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_l_r~0 .shared_arith = "off";

endmodule

module ddr3_int_altddio_out_4 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
inout 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_ddio_out_6ed_3 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module ddr3_int_ddio_out_6ed_3 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



arriaii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_ac_4 (
	phy_clk_1x,
	clk_3,
	dataout_0,
	seq_ac_add_1t_ac_lat_internal,
	period_sel_addr_7,
	seq_ac_sel,
	afi_addr_13,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	phy_clk_1x;
input 	clk_3;
output 	dataout_0;
input 	seq_ac_add_1t_ac_lat_internal;
input 	period_sel_addr_7;
input 	seq_ac_sel;
input 	afi_addr_13;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ac_l~q ;
wire \ac_2x_r~q ;
wire \ac_2x_2r~q ;
wire \ac_h_2r~q ;
wire \ac_l_2r~q ;
wire \ac_2x~0_combout ;
wire \ac_1t~q ;
wire \ac_2x_r~0_combout ;
wire \ac_h_r~q ;
wire \ac_l_r~q ;
wire \ac_h_r~0_combout ;
wire \ac_l_r~0_combout ;


ddr3_int_altddio_out_5 \half_rate.addr_pin (
	.outclock(clk_3),
	.dataout({dataout_0}),
	.datain_l({\ac_2x_r~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_l(
	.clk(phy_clk_1x),
	.d(GND_port),
	.asdata(afi_addr_13),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_l~q ),
	.prn(vcc));
defparam ac_l.is_wysiwyg = "true";
defparam ac_l.power_up = "low";

dffeas ac_2x_r(
	.clk(clk_3),
	.d(\ac_2x_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_r~q ),
	.prn(vcc));
defparam ac_2x_r.is_wysiwyg = "true";
defparam ac_2x_r.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_3),
	.d(\ac_2x_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

dffeas ac_h_2r(
	.clk(clk_3),
	.d(\ac_h_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_2r~q ),
	.prn(vcc));
defparam ac_h_2r.is_wysiwyg = "true";
defparam ac_h_2r.power_up = "low";

dffeas ac_l_2r(
	.clk(clk_3),
	.d(\ac_l_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_2r~q ),
	.prn(vcc));
defparam ac_l_2r.is_wysiwyg = "true";
defparam ac_l_2r.power_up = "low";

arriaii_lcell_comb \ac_2x~0 (
	.dataa(!period_sel_addr_7),
	.datab(!\ac_h_2r~q ),
	.datac(!\ac_l_2r~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x~0 .extended_lut = "off";
defparam \ac_2x~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \ac_2x~0 .shared_arith = "off";

dffeas ac_1t(
	.clk(clk_3),
	.d(\ac_2x~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

arriaii_lcell_comb \ac_2x_r~0 (
	.dataa(!seq_ac_add_1t_ac_lat_internal),
	.datab(!\ac_2x~0_combout ),
	.datac(!\ac_1t~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x_r~0 .extended_lut = "off";
defparam \ac_2x_r~0 .lut_mask = 64'h2727272727272727;
defparam \ac_2x_r~0 .shared_arith = "off";

dffeas ac_h_r(
	.clk(phy_clk_1x),
	.d(\ac_h_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_r~q ),
	.prn(vcc));
defparam ac_h_r.is_wysiwyg = "true";
defparam ac_h_r.power_up = "low";

dffeas ac_l_r(
	.clk(phy_clk_1x),
	.d(\ac_l_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_r~q ),
	.prn(vcc));
defparam ac_l_r.is_wysiwyg = "true";
defparam ac_l_r.power_up = "low";

arriaii_lcell_comb \ac_h_r~0 (
	.dataa(!\ac_l~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_h_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_h_r~0 .extended_lut = "off";
defparam \ac_h_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_h_r~0 .shared_arith = "off";

arriaii_lcell_comb \ac_l_r~0 (
	.dataa(!\ac_l~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_l_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_l_r~0 .extended_lut = "off";
defparam \ac_l_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_l_r~0 .shared_arith = "off";

endmodule

module ddr3_int_altddio_out_5 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
inout 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_ddio_out_6ed_4 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module ddr3_int_ddio_out_6ed_4 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



arriaii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_ac_5 (
	phy_clk_1x,
	clk_3,
	dataout_0,
	seq_ac_addr_1,
	seq_ac_addr_15,
	seq_ac_add_1t_ac_lat_internal,
	period_sel_addr_7,
	seq_ac_sel,
	afi_addr_1)/* synthesis synthesis_greybox=0 */;
input 	phy_clk_1x;
input 	clk_3;
output 	dataout_0;
input 	seq_ac_addr_1;
input 	seq_ac_addr_15;
input 	seq_ac_add_1t_ac_lat_internal;
input 	period_sel_addr_7;
input 	seq_ac_sel;
input 	afi_addr_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ac_h~q ;
wire \ac_l~q ;
wire \ac_2x_r~q ;
wire \ac_2x_2r~q ;
wire \ac_h_2r~q ;
wire \ac_l_2r~q ;
wire \ac_2x~0_combout ;
wire \ac_1t~q ;
wire \ac_2x_r~0_combout ;
wire \ac_h_r~q ;
wire \ac_l_r~q ;
wire \ac_h_r~0_combout ;
wire \ac_l_r~0_combout ;


ddr3_int_altddio_out_6 \half_rate.addr_pin (
	.outclock(clk_3),
	.dataout({dataout_0}),
	.datain_l({\ac_2x_r~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_h(
	.clk(phy_clk_1x),
	.d(seq_ac_addr_1),
	.asdata(afi_addr_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_h~q ),
	.prn(vcc));
defparam ac_h.is_wysiwyg = "true";
defparam ac_h.power_up = "low";

dffeas ac_l(
	.clk(phy_clk_1x),
	.d(seq_ac_addr_15),
	.asdata(afi_addr_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_l~q ),
	.prn(vcc));
defparam ac_l.is_wysiwyg = "true";
defparam ac_l.power_up = "low";

dffeas ac_2x_r(
	.clk(clk_3),
	.d(\ac_2x_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_r~q ),
	.prn(vcc));
defparam ac_2x_r.is_wysiwyg = "true";
defparam ac_2x_r.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_3),
	.d(\ac_2x_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

dffeas ac_h_2r(
	.clk(clk_3),
	.d(\ac_h_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_2r~q ),
	.prn(vcc));
defparam ac_h_2r.is_wysiwyg = "true";
defparam ac_h_2r.power_up = "low";

dffeas ac_l_2r(
	.clk(clk_3),
	.d(\ac_l_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_2r~q ),
	.prn(vcc));
defparam ac_l_2r.is_wysiwyg = "true";
defparam ac_l_2r.power_up = "low";

arriaii_lcell_comb \ac_2x~0 (
	.dataa(!period_sel_addr_7),
	.datab(!\ac_h_2r~q ),
	.datac(!\ac_l_2r~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x~0 .extended_lut = "off";
defparam \ac_2x~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \ac_2x~0 .shared_arith = "off";

dffeas ac_1t(
	.clk(clk_3),
	.d(\ac_2x~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

arriaii_lcell_comb \ac_2x_r~0 (
	.dataa(!seq_ac_add_1t_ac_lat_internal),
	.datab(!\ac_2x~0_combout ),
	.datac(!\ac_1t~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x_r~0 .extended_lut = "off";
defparam \ac_2x_r~0 .lut_mask = 64'h2727272727272727;
defparam \ac_2x_r~0 .shared_arith = "off";

dffeas ac_h_r(
	.clk(phy_clk_1x),
	.d(\ac_h_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_r~q ),
	.prn(vcc));
defparam ac_h_r.is_wysiwyg = "true";
defparam ac_h_r.power_up = "low";

dffeas ac_l_r(
	.clk(phy_clk_1x),
	.d(\ac_l_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_r~q ),
	.prn(vcc));
defparam ac_l_r.is_wysiwyg = "true";
defparam ac_l_r.power_up = "low";

arriaii_lcell_comb \ac_h_r~0 (
	.dataa(!\ac_h~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_h_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_h_r~0 .extended_lut = "off";
defparam \ac_h_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_h_r~0 .shared_arith = "off";

arriaii_lcell_comb \ac_l_r~0 (
	.dataa(!\ac_l~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_l_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_l_r~0 .extended_lut = "off";
defparam \ac_l_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_l_r~0 .shared_arith = "off";

endmodule

module ddr3_int_altddio_out_6 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
inout 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_ddio_out_6ed_5 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module ddr3_int_ddio_out_6ed_5 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



arriaii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_ac_6 (
	phy_clk_1x,
	clk_3,
	dataout_0,
	seq_ac_addr_16,
	seq_ac_add_1t_ac_lat_internal,
	period_sel_addr_7,
	seq_ac_sel,
	afi_addr_2)/* synthesis synthesis_greybox=0 */;
input 	phy_clk_1x;
input 	clk_3;
output 	dataout_0;
input 	seq_ac_addr_16;
input 	seq_ac_add_1t_ac_lat_internal;
input 	period_sel_addr_7;
input 	seq_ac_sel;
input 	afi_addr_2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ac_l~q ;
wire \ac_2x_r~q ;
wire \ac_2x_2r~q ;
wire \ac_h_2r~q ;
wire \ac_l_2r~q ;
wire \ac_2x~0_combout ;
wire \ac_1t~q ;
wire \ac_2x_r~0_combout ;
wire \ac_h_r~q ;
wire \ac_l_r~q ;
wire \ac_h_r~0_combout ;
wire \ac_l_r~0_combout ;


ddr3_int_altddio_out_7 \half_rate.addr_pin (
	.outclock(clk_3),
	.dataout({dataout_0}),
	.datain_l({\ac_2x_r~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_l(
	.clk(phy_clk_1x),
	.d(seq_ac_addr_16),
	.asdata(afi_addr_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_l~q ),
	.prn(vcc));
defparam ac_l.is_wysiwyg = "true";
defparam ac_l.power_up = "low";

dffeas ac_2x_r(
	.clk(clk_3),
	.d(\ac_2x_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_r~q ),
	.prn(vcc));
defparam ac_2x_r.is_wysiwyg = "true";
defparam ac_2x_r.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_3),
	.d(\ac_2x_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

dffeas ac_h_2r(
	.clk(clk_3),
	.d(\ac_h_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_2r~q ),
	.prn(vcc));
defparam ac_h_2r.is_wysiwyg = "true";
defparam ac_h_2r.power_up = "low";

dffeas ac_l_2r(
	.clk(clk_3),
	.d(\ac_l_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_2r~q ),
	.prn(vcc));
defparam ac_l_2r.is_wysiwyg = "true";
defparam ac_l_2r.power_up = "low";

arriaii_lcell_comb \ac_2x~0 (
	.dataa(!period_sel_addr_7),
	.datab(!\ac_h_2r~q ),
	.datac(!\ac_l_2r~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x~0 .extended_lut = "off";
defparam \ac_2x~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \ac_2x~0 .shared_arith = "off";

dffeas ac_1t(
	.clk(clk_3),
	.d(\ac_2x~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

arriaii_lcell_comb \ac_2x_r~0 (
	.dataa(!seq_ac_add_1t_ac_lat_internal),
	.datab(!\ac_2x~0_combout ),
	.datac(!\ac_1t~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x_r~0 .extended_lut = "off";
defparam \ac_2x_r~0 .lut_mask = 64'h2727272727272727;
defparam \ac_2x_r~0 .shared_arith = "off";

dffeas ac_h_r(
	.clk(phy_clk_1x),
	.d(\ac_h_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_r~q ),
	.prn(vcc));
defparam ac_h_r.is_wysiwyg = "true";
defparam ac_h_r.power_up = "low";

dffeas ac_l_r(
	.clk(phy_clk_1x),
	.d(\ac_l_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_r~q ),
	.prn(vcc));
defparam ac_l_r.is_wysiwyg = "true";
defparam ac_l_r.power_up = "low";

arriaii_lcell_comb \ac_h_r~0 (
	.dataa(!\ac_l~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_h_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_h_r~0 .extended_lut = "off";
defparam \ac_h_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_h_r~0 .shared_arith = "off";

arriaii_lcell_comb \ac_l_r~0 (
	.dataa(!\ac_l~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_l_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_l_r~0 .extended_lut = "off";
defparam \ac_l_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_l_r~0 .shared_arith = "off";

endmodule

module ddr3_int_altddio_out_7 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
inout 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_ddio_out_6ed_6 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module ddr3_int_ddio_out_6ed_6 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



arriaii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_ac_7 (
	phy_clk_1x,
	clk_3,
	dataout_0,
	seq_ac_addr_17,
	seq_ac_add_1t_ac_lat_internal,
	period_sel_addr_7,
	seq_ac_sel,
	afi_addr_3)/* synthesis synthesis_greybox=0 */;
input 	phy_clk_1x;
input 	clk_3;
output 	dataout_0;
input 	seq_ac_addr_17;
input 	seq_ac_add_1t_ac_lat_internal;
input 	period_sel_addr_7;
input 	seq_ac_sel;
input 	afi_addr_3;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ac_l~q ;
wire \ac_2x_r~q ;
wire \ac_2x_2r~q ;
wire \ac_h_2r~q ;
wire \ac_l_2r~q ;
wire \ac_2x~0_combout ;
wire \ac_1t~q ;
wire \ac_2x_r~0_combout ;
wire \ac_h_r~q ;
wire \ac_l_r~q ;
wire \ac_h_r~0_combout ;
wire \ac_l_r~0_combout ;


ddr3_int_altddio_out_8 \half_rate.addr_pin (
	.outclock(clk_3),
	.dataout({dataout_0}),
	.datain_l({\ac_2x_r~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_l(
	.clk(phy_clk_1x),
	.d(seq_ac_addr_17),
	.asdata(afi_addr_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_l~q ),
	.prn(vcc));
defparam ac_l.is_wysiwyg = "true";
defparam ac_l.power_up = "low";

dffeas ac_2x_r(
	.clk(clk_3),
	.d(\ac_2x_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_r~q ),
	.prn(vcc));
defparam ac_2x_r.is_wysiwyg = "true";
defparam ac_2x_r.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_3),
	.d(\ac_2x_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

dffeas ac_h_2r(
	.clk(clk_3),
	.d(\ac_h_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_2r~q ),
	.prn(vcc));
defparam ac_h_2r.is_wysiwyg = "true";
defparam ac_h_2r.power_up = "low";

dffeas ac_l_2r(
	.clk(clk_3),
	.d(\ac_l_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_2r~q ),
	.prn(vcc));
defparam ac_l_2r.is_wysiwyg = "true";
defparam ac_l_2r.power_up = "low";

arriaii_lcell_comb \ac_2x~0 (
	.dataa(!period_sel_addr_7),
	.datab(!\ac_h_2r~q ),
	.datac(!\ac_l_2r~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x~0 .extended_lut = "off";
defparam \ac_2x~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \ac_2x~0 .shared_arith = "off";

dffeas ac_1t(
	.clk(clk_3),
	.d(\ac_2x~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

arriaii_lcell_comb \ac_2x_r~0 (
	.dataa(!seq_ac_add_1t_ac_lat_internal),
	.datab(!\ac_2x~0_combout ),
	.datac(!\ac_1t~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x_r~0 .extended_lut = "off";
defparam \ac_2x_r~0 .lut_mask = 64'h2727272727272727;
defparam \ac_2x_r~0 .shared_arith = "off";

dffeas ac_h_r(
	.clk(phy_clk_1x),
	.d(\ac_h_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_r~q ),
	.prn(vcc));
defparam ac_h_r.is_wysiwyg = "true";
defparam ac_h_r.power_up = "low";

dffeas ac_l_r(
	.clk(phy_clk_1x),
	.d(\ac_l_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_r~q ),
	.prn(vcc));
defparam ac_l_r.is_wysiwyg = "true";
defparam ac_l_r.power_up = "low";

arriaii_lcell_comb \ac_h_r~0 (
	.dataa(!\ac_l~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_h_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_h_r~0 .extended_lut = "off";
defparam \ac_h_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_h_r~0 .shared_arith = "off";

arriaii_lcell_comb \ac_l_r~0 (
	.dataa(!\ac_l~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_l_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_l_r~0 .extended_lut = "off";
defparam \ac_l_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_l_r~0 .shared_arith = "off";

endmodule

module ddr3_int_altddio_out_8 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
inout 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_ddio_out_6ed_7 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module ddr3_int_ddio_out_6ed_7 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



arriaii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_ac_8 (
	phy_clk_1x,
	clk_3,
	dataout_0,
	seq_ac_addr_18,
	seq_ac_add_1t_ac_lat_internal,
	period_sel_addr_7,
	seq_ac_sel,
	afi_addr_4)/* synthesis synthesis_greybox=0 */;
input 	phy_clk_1x;
input 	clk_3;
output 	dataout_0;
input 	seq_ac_addr_18;
input 	seq_ac_add_1t_ac_lat_internal;
input 	period_sel_addr_7;
input 	seq_ac_sel;
input 	afi_addr_4;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ac_l~q ;
wire \ac_2x_r~q ;
wire \ac_2x_2r~q ;
wire \ac_h_2r~q ;
wire \ac_l_2r~q ;
wire \ac_2x~0_combout ;
wire \ac_1t~q ;
wire \ac_2x_r~0_combout ;
wire \ac_h_r~q ;
wire \ac_l_r~q ;
wire \ac_h_r~0_combout ;
wire \ac_l_r~0_combout ;


ddr3_int_altddio_out_9 \half_rate.addr_pin (
	.outclock(clk_3),
	.dataout({dataout_0}),
	.datain_l({\ac_2x_r~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_l(
	.clk(phy_clk_1x),
	.d(seq_ac_addr_18),
	.asdata(afi_addr_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_l~q ),
	.prn(vcc));
defparam ac_l.is_wysiwyg = "true";
defparam ac_l.power_up = "low";

dffeas ac_2x_r(
	.clk(clk_3),
	.d(\ac_2x_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_r~q ),
	.prn(vcc));
defparam ac_2x_r.is_wysiwyg = "true";
defparam ac_2x_r.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_3),
	.d(\ac_2x_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

dffeas ac_h_2r(
	.clk(clk_3),
	.d(\ac_h_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_2r~q ),
	.prn(vcc));
defparam ac_h_2r.is_wysiwyg = "true";
defparam ac_h_2r.power_up = "low";

dffeas ac_l_2r(
	.clk(clk_3),
	.d(\ac_l_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_2r~q ),
	.prn(vcc));
defparam ac_l_2r.is_wysiwyg = "true";
defparam ac_l_2r.power_up = "low";

arriaii_lcell_comb \ac_2x~0 (
	.dataa(!period_sel_addr_7),
	.datab(!\ac_h_2r~q ),
	.datac(!\ac_l_2r~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x~0 .extended_lut = "off";
defparam \ac_2x~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \ac_2x~0 .shared_arith = "off";

dffeas ac_1t(
	.clk(clk_3),
	.d(\ac_2x~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

arriaii_lcell_comb \ac_2x_r~0 (
	.dataa(!seq_ac_add_1t_ac_lat_internal),
	.datab(!\ac_2x~0_combout ),
	.datac(!\ac_1t~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x_r~0 .extended_lut = "off";
defparam \ac_2x_r~0 .lut_mask = 64'h2727272727272727;
defparam \ac_2x_r~0 .shared_arith = "off";

dffeas ac_h_r(
	.clk(phy_clk_1x),
	.d(\ac_h_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_r~q ),
	.prn(vcc));
defparam ac_h_r.is_wysiwyg = "true";
defparam ac_h_r.power_up = "low";

dffeas ac_l_r(
	.clk(phy_clk_1x),
	.d(\ac_l_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_r~q ),
	.prn(vcc));
defparam ac_l_r.is_wysiwyg = "true";
defparam ac_l_r.power_up = "low";

arriaii_lcell_comb \ac_h_r~0 (
	.dataa(!\ac_l~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_h_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_h_r~0 .extended_lut = "off";
defparam \ac_h_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_h_r~0 .shared_arith = "off";

arriaii_lcell_comb \ac_l_r~0 (
	.dataa(!\ac_l~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_l_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_l_r~0 .extended_lut = "off";
defparam \ac_l_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_l_r~0 .shared_arith = "off";

endmodule

module ddr3_int_altddio_out_9 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
inout 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_ddio_out_6ed_8 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module ddr3_int_ddio_out_6ed_8 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



arriaii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_ac_9 (
	phy_clk_1x,
	clk_3,
	dataout_0,
	seq_ac_addr_5,
	seq_ac_addr_19,
	seq_ac_add_1t_ac_lat_internal,
	period_sel_addr_7,
	seq_ac_sel,
	afi_addr_5)/* synthesis synthesis_greybox=0 */;
input 	phy_clk_1x;
input 	clk_3;
output 	dataout_0;
input 	seq_ac_addr_5;
input 	seq_ac_addr_19;
input 	seq_ac_add_1t_ac_lat_internal;
input 	period_sel_addr_7;
input 	seq_ac_sel;
input 	afi_addr_5;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ac_h~q ;
wire \ac_l~q ;
wire \ac_2x_r~q ;
wire \ac_2x_2r~q ;
wire \ac_h_2r~q ;
wire \ac_l_2r~q ;
wire \ac_2x~0_combout ;
wire \ac_1t~q ;
wire \ac_2x_r~0_combout ;
wire \ac_h_r~q ;
wire \ac_l_r~q ;
wire \ac_h_r~0_combout ;
wire \ac_l_r~0_combout ;


ddr3_int_altddio_out_10 \half_rate.addr_pin (
	.outclock(clk_3),
	.dataout({dataout_0}),
	.datain_l({\ac_2x_r~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_h(
	.clk(phy_clk_1x),
	.d(seq_ac_addr_5),
	.asdata(afi_addr_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_h~q ),
	.prn(vcc));
defparam ac_h.is_wysiwyg = "true";
defparam ac_h.power_up = "low";

dffeas ac_l(
	.clk(phy_clk_1x),
	.d(seq_ac_addr_19),
	.asdata(afi_addr_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_l~q ),
	.prn(vcc));
defparam ac_l.is_wysiwyg = "true";
defparam ac_l.power_up = "low";

dffeas ac_2x_r(
	.clk(clk_3),
	.d(\ac_2x_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_r~q ),
	.prn(vcc));
defparam ac_2x_r.is_wysiwyg = "true";
defparam ac_2x_r.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_3),
	.d(\ac_2x_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

dffeas ac_h_2r(
	.clk(clk_3),
	.d(\ac_h_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_2r~q ),
	.prn(vcc));
defparam ac_h_2r.is_wysiwyg = "true";
defparam ac_h_2r.power_up = "low";

dffeas ac_l_2r(
	.clk(clk_3),
	.d(\ac_l_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_2r~q ),
	.prn(vcc));
defparam ac_l_2r.is_wysiwyg = "true";
defparam ac_l_2r.power_up = "low";

arriaii_lcell_comb \ac_2x~0 (
	.dataa(!period_sel_addr_7),
	.datab(!\ac_h_2r~q ),
	.datac(!\ac_l_2r~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x~0 .extended_lut = "off";
defparam \ac_2x~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \ac_2x~0 .shared_arith = "off";

dffeas ac_1t(
	.clk(clk_3),
	.d(\ac_2x~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

arriaii_lcell_comb \ac_2x_r~0 (
	.dataa(!seq_ac_add_1t_ac_lat_internal),
	.datab(!\ac_2x~0_combout ),
	.datac(!\ac_1t~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x_r~0 .extended_lut = "off";
defparam \ac_2x_r~0 .lut_mask = 64'h2727272727272727;
defparam \ac_2x_r~0 .shared_arith = "off";

dffeas ac_h_r(
	.clk(phy_clk_1x),
	.d(\ac_h_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_r~q ),
	.prn(vcc));
defparam ac_h_r.is_wysiwyg = "true";
defparam ac_h_r.power_up = "low";

dffeas ac_l_r(
	.clk(phy_clk_1x),
	.d(\ac_l_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_r~q ),
	.prn(vcc));
defparam ac_l_r.is_wysiwyg = "true";
defparam ac_l_r.power_up = "low";

arriaii_lcell_comb \ac_h_r~0 (
	.dataa(!\ac_h~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_h_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_h_r~0 .extended_lut = "off";
defparam \ac_h_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_h_r~0 .shared_arith = "off";

arriaii_lcell_comb \ac_l_r~0 (
	.dataa(!\ac_l~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_l_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_l_r~0 .extended_lut = "off";
defparam \ac_l_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_l_r~0 .shared_arith = "off";

endmodule

module ddr3_int_altddio_out_10 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
inout 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_ddio_out_6ed_9 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module ddr3_int_ddio_out_6ed_9 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



arriaii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_ac_10 (
	phy_clk_1x,
	clk_3,
	dataout_0,
	seq_ac_add_1t_ac_lat_internal,
	period_sel_addr_7,
	seq_ac_sel,
	afi_addr_6,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	phy_clk_1x;
input 	clk_3;
output 	dataout_0;
input 	seq_ac_add_1t_ac_lat_internal;
input 	period_sel_addr_7;
input 	seq_ac_sel;
input 	afi_addr_6;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ac_l~q ;
wire \ac_2x_r~q ;
wire \ac_2x_2r~q ;
wire \ac_h_2r~q ;
wire \ac_l_2r~q ;
wire \ac_2x~0_combout ;
wire \ac_1t~q ;
wire \ac_2x_r~0_combout ;
wire \ac_h_r~q ;
wire \ac_l_r~q ;
wire \ac_h_r~0_combout ;
wire \ac_l_r~0_combout ;


ddr3_int_altddio_out_11 \half_rate.addr_pin (
	.outclock(clk_3),
	.dataout({dataout_0}),
	.datain_l({\ac_2x_r~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_l(
	.clk(phy_clk_1x),
	.d(GND_port),
	.asdata(afi_addr_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_l~q ),
	.prn(vcc));
defparam ac_l.is_wysiwyg = "true";
defparam ac_l.power_up = "low";

dffeas ac_2x_r(
	.clk(clk_3),
	.d(\ac_2x_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_r~q ),
	.prn(vcc));
defparam ac_2x_r.is_wysiwyg = "true";
defparam ac_2x_r.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_3),
	.d(\ac_2x_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

dffeas ac_h_2r(
	.clk(clk_3),
	.d(\ac_h_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_2r~q ),
	.prn(vcc));
defparam ac_h_2r.is_wysiwyg = "true";
defparam ac_h_2r.power_up = "low";

dffeas ac_l_2r(
	.clk(clk_3),
	.d(\ac_l_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_2r~q ),
	.prn(vcc));
defparam ac_l_2r.is_wysiwyg = "true";
defparam ac_l_2r.power_up = "low";

arriaii_lcell_comb \ac_2x~0 (
	.dataa(!period_sel_addr_7),
	.datab(!\ac_h_2r~q ),
	.datac(!\ac_l_2r~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x~0 .extended_lut = "off";
defparam \ac_2x~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \ac_2x~0 .shared_arith = "off";

dffeas ac_1t(
	.clk(clk_3),
	.d(\ac_2x~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

arriaii_lcell_comb \ac_2x_r~0 (
	.dataa(!seq_ac_add_1t_ac_lat_internal),
	.datab(!\ac_2x~0_combout ),
	.datac(!\ac_1t~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x_r~0 .extended_lut = "off";
defparam \ac_2x_r~0 .lut_mask = 64'h2727272727272727;
defparam \ac_2x_r~0 .shared_arith = "off";

dffeas ac_h_r(
	.clk(phy_clk_1x),
	.d(\ac_h_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_r~q ),
	.prn(vcc));
defparam ac_h_r.is_wysiwyg = "true";
defparam ac_h_r.power_up = "low";

dffeas ac_l_r(
	.clk(phy_clk_1x),
	.d(\ac_l_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_r~q ),
	.prn(vcc));
defparam ac_l_r.is_wysiwyg = "true";
defparam ac_l_r.power_up = "low";

arriaii_lcell_comb \ac_h_r~0 (
	.dataa(!\ac_l~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_h_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_h_r~0 .extended_lut = "off";
defparam \ac_h_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_h_r~0 .shared_arith = "off";

arriaii_lcell_comb \ac_l_r~0 (
	.dataa(!\ac_l~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_l_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_l_r~0 .extended_lut = "off";
defparam \ac_l_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_l_r~0 .shared_arith = "off";

endmodule

module ddr3_int_altddio_out_11 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
inout 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_ddio_out_6ed_10 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module ddr3_int_ddio_out_6ed_10 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



arriaii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_ac_11 (
	phy_clk_1x,
	clk_3,
	dataout_0,
	seq_ac_add_1t_ac_lat_internal,
	period_sel_addr_7,
	seq_ac_sel,
	afi_addr_7,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	phy_clk_1x;
input 	clk_3;
output 	dataout_0;
input 	seq_ac_add_1t_ac_lat_internal;
input 	period_sel_addr_7;
input 	seq_ac_sel;
input 	afi_addr_7;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ac_l~q ;
wire \ac_2x_r~q ;
wire \ac_2x_2r~q ;
wire \ac_h_2r~q ;
wire \ac_l_2r~q ;
wire \ac_2x~0_combout ;
wire \ac_1t~q ;
wire \ac_2x_r~0_combout ;
wire \ac_h_r~q ;
wire \ac_l_r~q ;
wire \ac_h_r~0_combout ;
wire \ac_l_r~0_combout ;


ddr3_int_altddio_out_12 \half_rate.addr_pin (
	.outclock(clk_3),
	.dataout({dataout_0}),
	.datain_l({\ac_2x_r~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_l(
	.clk(phy_clk_1x),
	.d(GND_port),
	.asdata(afi_addr_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_l~q ),
	.prn(vcc));
defparam ac_l.is_wysiwyg = "true";
defparam ac_l.power_up = "low";

dffeas ac_2x_r(
	.clk(clk_3),
	.d(\ac_2x_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_r~q ),
	.prn(vcc));
defparam ac_2x_r.is_wysiwyg = "true";
defparam ac_2x_r.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_3),
	.d(\ac_2x_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

dffeas ac_h_2r(
	.clk(clk_3),
	.d(\ac_h_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_2r~q ),
	.prn(vcc));
defparam ac_h_2r.is_wysiwyg = "true";
defparam ac_h_2r.power_up = "low";

dffeas ac_l_2r(
	.clk(clk_3),
	.d(\ac_l_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_2r~q ),
	.prn(vcc));
defparam ac_l_2r.is_wysiwyg = "true";
defparam ac_l_2r.power_up = "low";

arriaii_lcell_comb \ac_2x~0 (
	.dataa(!period_sel_addr_7),
	.datab(!\ac_h_2r~q ),
	.datac(!\ac_l_2r~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x~0 .extended_lut = "off";
defparam \ac_2x~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \ac_2x~0 .shared_arith = "off";

dffeas ac_1t(
	.clk(clk_3),
	.d(\ac_2x~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

arriaii_lcell_comb \ac_2x_r~0 (
	.dataa(!seq_ac_add_1t_ac_lat_internal),
	.datab(!\ac_2x~0_combout ),
	.datac(!\ac_1t~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x_r~0 .extended_lut = "off";
defparam \ac_2x_r~0 .lut_mask = 64'h2727272727272727;
defparam \ac_2x_r~0 .shared_arith = "off";

dffeas ac_h_r(
	.clk(phy_clk_1x),
	.d(\ac_h_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_r~q ),
	.prn(vcc));
defparam ac_h_r.is_wysiwyg = "true";
defparam ac_h_r.power_up = "low";

dffeas ac_l_r(
	.clk(phy_clk_1x),
	.d(\ac_l_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_r~q ),
	.prn(vcc));
defparam ac_l_r.is_wysiwyg = "true";
defparam ac_l_r.power_up = "low";

arriaii_lcell_comb \ac_h_r~0 (
	.dataa(!\ac_l~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_h_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_h_r~0 .extended_lut = "off";
defparam \ac_h_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_h_r~0 .shared_arith = "off";

arriaii_lcell_comb \ac_l_r~0 (
	.dataa(!\ac_l~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_l_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_l_r~0 .extended_lut = "off";
defparam \ac_l_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_l_r~0 .shared_arith = "off";

endmodule

module ddr3_int_altddio_out_12 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
inout 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_ddio_out_6ed_11 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module ddr3_int_ddio_out_6ed_11 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



arriaii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_ac_12 (
	phy_clk_1x,
	clk_3,
	dataout_0,
	seq_ac_addr_8,
	seq_ac_addr_22,
	seq_ac_add_1t_ac_lat_internal,
	period_sel_addr_7,
	seq_ac_sel,
	afi_addr_8)/* synthesis synthesis_greybox=0 */;
input 	phy_clk_1x;
input 	clk_3;
output 	dataout_0;
input 	seq_ac_addr_8;
input 	seq_ac_addr_22;
input 	seq_ac_add_1t_ac_lat_internal;
input 	period_sel_addr_7;
input 	seq_ac_sel;
input 	afi_addr_8;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ac_h~q ;
wire \ac_l~q ;
wire \ac_2x_r~q ;
wire \ac_2x_2r~q ;
wire \ac_h_2r~q ;
wire \ac_l_2r~q ;
wire \ac_2x~0_combout ;
wire \ac_1t~q ;
wire \ac_2x_r~0_combout ;
wire \ac_h_r~q ;
wire \ac_l_r~q ;
wire \ac_h_r~0_combout ;
wire \ac_l_r~0_combout ;


ddr3_int_altddio_out_13 \half_rate.addr_pin (
	.outclock(clk_3),
	.dataout({dataout_0}),
	.datain_l({\ac_2x_r~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_h(
	.clk(phy_clk_1x),
	.d(seq_ac_addr_8),
	.asdata(afi_addr_8),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_h~q ),
	.prn(vcc));
defparam ac_h.is_wysiwyg = "true";
defparam ac_h.power_up = "low";

dffeas ac_l(
	.clk(phy_clk_1x),
	.d(seq_ac_addr_22),
	.asdata(afi_addr_8),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_l~q ),
	.prn(vcc));
defparam ac_l.is_wysiwyg = "true";
defparam ac_l.power_up = "low";

dffeas ac_2x_r(
	.clk(clk_3),
	.d(\ac_2x_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_r~q ),
	.prn(vcc));
defparam ac_2x_r.is_wysiwyg = "true";
defparam ac_2x_r.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_3),
	.d(\ac_2x_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

dffeas ac_h_2r(
	.clk(clk_3),
	.d(\ac_h_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_2r~q ),
	.prn(vcc));
defparam ac_h_2r.is_wysiwyg = "true";
defparam ac_h_2r.power_up = "low";

dffeas ac_l_2r(
	.clk(clk_3),
	.d(\ac_l_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_2r~q ),
	.prn(vcc));
defparam ac_l_2r.is_wysiwyg = "true";
defparam ac_l_2r.power_up = "low";

arriaii_lcell_comb \ac_2x~0 (
	.dataa(!period_sel_addr_7),
	.datab(!\ac_h_2r~q ),
	.datac(!\ac_l_2r~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x~0 .extended_lut = "off";
defparam \ac_2x~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \ac_2x~0 .shared_arith = "off";

dffeas ac_1t(
	.clk(clk_3),
	.d(\ac_2x~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

arriaii_lcell_comb \ac_2x_r~0 (
	.dataa(!seq_ac_add_1t_ac_lat_internal),
	.datab(!\ac_2x~0_combout ),
	.datac(!\ac_1t~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x_r~0 .extended_lut = "off";
defparam \ac_2x_r~0 .lut_mask = 64'h2727272727272727;
defparam \ac_2x_r~0 .shared_arith = "off";

dffeas ac_h_r(
	.clk(phy_clk_1x),
	.d(\ac_h_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_r~q ),
	.prn(vcc));
defparam ac_h_r.is_wysiwyg = "true";
defparam ac_h_r.power_up = "low";

dffeas ac_l_r(
	.clk(phy_clk_1x),
	.d(\ac_l_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_r~q ),
	.prn(vcc));
defparam ac_l_r.is_wysiwyg = "true";
defparam ac_l_r.power_up = "low";

arriaii_lcell_comb \ac_h_r~0 (
	.dataa(!\ac_h~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_h_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_h_r~0 .extended_lut = "off";
defparam \ac_h_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_h_r~0 .shared_arith = "off";

arriaii_lcell_comb \ac_l_r~0 (
	.dataa(!\ac_l~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_l_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_l_r~0 .extended_lut = "off";
defparam \ac_l_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_l_r~0 .shared_arith = "off";

endmodule

module ddr3_int_altddio_out_13 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
inout 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_ddio_out_6ed_12 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module ddr3_int_ddio_out_6ed_12 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



arriaii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_ac_13 (
	phy_clk_1x,
	clk_3,
	dataout_0,
	seq_ac_addr_0,
	seq_ac_addr_14,
	seq_ac_add_1t_ac_lat_internal,
	period_sel_addr_7,
	seq_ac_sel,
	afi_addr_9)/* synthesis synthesis_greybox=0 */;
input 	phy_clk_1x;
input 	clk_3;
output 	dataout_0;
input 	seq_ac_addr_0;
input 	seq_ac_addr_14;
input 	seq_ac_add_1t_ac_lat_internal;
input 	period_sel_addr_7;
input 	seq_ac_sel;
input 	afi_addr_9;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ac_h~q ;
wire \ac_l~q ;
wire \ac_2x_r~q ;
wire \ac_2x_2r~q ;
wire \ac_h_2r~q ;
wire \ac_l_2r~q ;
wire \ac_2x~0_combout ;
wire \ac_1t~q ;
wire \ac_2x_r~0_combout ;
wire \ac_h_r~q ;
wire \ac_l_r~q ;
wire \ac_h_r~0_combout ;
wire \ac_l_r~0_combout ;


ddr3_int_altddio_out_14 \half_rate.addr_pin (
	.outclock(clk_3),
	.dataout({dataout_0}),
	.datain_l({\ac_2x_r~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_h(
	.clk(phy_clk_1x),
	.d(seq_ac_addr_0),
	.asdata(afi_addr_9),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_h~q ),
	.prn(vcc));
defparam ac_h.is_wysiwyg = "true";
defparam ac_h.power_up = "low";

dffeas ac_l(
	.clk(phy_clk_1x),
	.d(seq_ac_addr_14),
	.asdata(afi_addr_9),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_l~q ),
	.prn(vcc));
defparam ac_l.is_wysiwyg = "true";
defparam ac_l.power_up = "low";

dffeas ac_2x_r(
	.clk(clk_3),
	.d(\ac_2x_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_r~q ),
	.prn(vcc));
defparam ac_2x_r.is_wysiwyg = "true";
defparam ac_2x_r.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_3),
	.d(\ac_2x_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

dffeas ac_h_2r(
	.clk(clk_3),
	.d(\ac_h_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_2r~q ),
	.prn(vcc));
defparam ac_h_2r.is_wysiwyg = "true";
defparam ac_h_2r.power_up = "low";

dffeas ac_l_2r(
	.clk(clk_3),
	.d(\ac_l_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_2r~q ),
	.prn(vcc));
defparam ac_l_2r.is_wysiwyg = "true";
defparam ac_l_2r.power_up = "low";

arriaii_lcell_comb \ac_2x~0 (
	.dataa(!period_sel_addr_7),
	.datab(!\ac_h_2r~q ),
	.datac(!\ac_l_2r~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x~0 .extended_lut = "off";
defparam \ac_2x~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \ac_2x~0 .shared_arith = "off";

dffeas ac_1t(
	.clk(clk_3),
	.d(\ac_2x~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

arriaii_lcell_comb \ac_2x_r~0 (
	.dataa(!seq_ac_add_1t_ac_lat_internal),
	.datab(!\ac_2x~0_combout ),
	.datac(!\ac_1t~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x_r~0 .extended_lut = "off";
defparam \ac_2x_r~0 .lut_mask = 64'h2727272727272727;
defparam \ac_2x_r~0 .shared_arith = "off";

dffeas ac_h_r(
	.clk(phy_clk_1x),
	.d(\ac_h_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_r~q ),
	.prn(vcc));
defparam ac_h_r.is_wysiwyg = "true";
defparam ac_h_r.power_up = "low";

dffeas ac_l_r(
	.clk(phy_clk_1x),
	.d(\ac_l_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_r~q ),
	.prn(vcc));
defparam ac_l_r.is_wysiwyg = "true";
defparam ac_l_r.power_up = "low";

arriaii_lcell_comb \ac_h_r~0 (
	.dataa(!\ac_h~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_h_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_h_r~0 .extended_lut = "off";
defparam \ac_h_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_h_r~0 .shared_arith = "off";

arriaii_lcell_comb \ac_l_r~0 (
	.dataa(!\ac_l~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_l_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_l_r~0 .extended_lut = "off";
defparam \ac_l_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_l_r~0 .shared_arith = "off";

endmodule

module ddr3_int_altddio_out_14 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
inout 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_ddio_out_6ed_13 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module ddr3_int_ddio_out_6ed_13 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



arriaii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_ac_14 (
	phy_clk_1x,
	clk_3,
	dataout_0,
	seq_ac_ba_0,
	seq_ac_ba_3,
	seq_ac_add_1t_ac_lat_internal,
	period_sel_addr_7,
	seq_ac_sel,
	afi_ba_0)/* synthesis synthesis_greybox=0 */;
input 	phy_clk_1x;
input 	clk_3;
output 	dataout_0;
input 	seq_ac_ba_0;
input 	seq_ac_ba_3;
input 	seq_ac_add_1t_ac_lat_internal;
input 	period_sel_addr_7;
input 	seq_ac_sel;
input 	afi_ba_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ac_h~q ;
wire \ac_l~q ;
wire \ac_2x_r~q ;
wire \ac_2x_2r~q ;
wire \ac_h_2r~q ;
wire \ac_l_2r~q ;
wire \ac_2x~0_combout ;
wire \ac_1t~q ;
wire \ac_2x_r~0_combout ;
wire \ac_h_r~q ;
wire \ac_l_r~q ;


ddr3_int_altddio_out_15 \half_rate.addr_pin (
	.outclock(clk_3),
	.dataout({dataout_0}),
	.datain_l({\ac_2x_r~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_h(
	.clk(phy_clk_1x),
	.d(seq_ac_ba_0),
	.asdata(afi_ba_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_h~q ),
	.prn(vcc));
defparam ac_h.is_wysiwyg = "true";
defparam ac_h.power_up = "low";

dffeas ac_l(
	.clk(phy_clk_1x),
	.d(seq_ac_ba_3),
	.asdata(afi_ba_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_l~q ),
	.prn(vcc));
defparam ac_l.is_wysiwyg = "true";
defparam ac_l.power_up = "low";

dffeas ac_2x_r(
	.clk(clk_3),
	.d(\ac_2x_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_r~q ),
	.prn(vcc));
defparam ac_2x_r.is_wysiwyg = "true";
defparam ac_2x_r.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_3),
	.d(\ac_2x_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

dffeas ac_h_2r(
	.clk(clk_3),
	.d(\ac_h_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_2r~q ),
	.prn(vcc));
defparam ac_h_2r.is_wysiwyg = "true";
defparam ac_h_2r.power_up = "low";

dffeas ac_l_2r(
	.clk(clk_3),
	.d(\ac_l_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_2r~q ),
	.prn(vcc));
defparam ac_l_2r.is_wysiwyg = "true";
defparam ac_l_2r.power_up = "low";

arriaii_lcell_comb \ac_2x~0 (
	.dataa(!period_sel_addr_7),
	.datab(!\ac_h_2r~q ),
	.datac(!\ac_l_2r~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x~0 .extended_lut = "off";
defparam \ac_2x~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \ac_2x~0 .shared_arith = "off";

dffeas ac_1t(
	.clk(clk_3),
	.d(\ac_2x~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

arriaii_lcell_comb \ac_2x_r~0 (
	.dataa(!seq_ac_add_1t_ac_lat_internal),
	.datab(!\ac_2x~0_combout ),
	.datac(!\ac_1t~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x_r~0 .extended_lut = "off";
defparam \ac_2x_r~0 .lut_mask = 64'h2727272727272727;
defparam \ac_2x_r~0 .shared_arith = "off";

dffeas ac_h_r(
	.clk(phy_clk_1x),
	.d(\ac_h~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_r~q ),
	.prn(vcc));
defparam ac_h_r.is_wysiwyg = "true";
defparam ac_h_r.power_up = "low";

dffeas ac_l_r(
	.clk(phy_clk_1x),
	.d(\ac_l~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_r~q ),
	.prn(vcc));
defparam ac_l_r.is_wysiwyg = "true";
defparam ac_l_r.power_up = "low";

endmodule

module ddr3_int_altddio_out_15 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
inout 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_ddio_out_pgd auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module ddr3_int_ddio_out_pgd (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



arriaii_ddio_out \ddio_outa[0] (
	.datainlo(datain_l[0]),
	.datainhi(datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "clear";
defparam \ddio_outa[0] .power_up = "low";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_ac_15 (
	phy_clk_1x,
	clk_3,
	dataout_0,
	seq_ac_ba_1,
	seq_ac_ba_4,
	seq_ac_add_1t_ac_lat_internal,
	period_sel_addr_7,
	seq_ac_sel,
	afi_ba_1)/* synthesis synthesis_greybox=0 */;
input 	phy_clk_1x;
input 	clk_3;
output 	dataout_0;
input 	seq_ac_ba_1;
input 	seq_ac_ba_4;
input 	seq_ac_add_1t_ac_lat_internal;
input 	period_sel_addr_7;
input 	seq_ac_sel;
input 	afi_ba_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ac_h~q ;
wire \ac_l~q ;
wire \ac_2x_r~q ;
wire \ac_2x_2r~q ;
wire \ac_h_2r~q ;
wire \ac_l_2r~q ;
wire \ac_2x~0_combout ;
wire \ac_1t~q ;
wire \ac_2x_r~0_combout ;
wire \ac_h_r~q ;
wire \ac_l_r~q ;


ddr3_int_altddio_out_16 \half_rate.addr_pin (
	.outclock(clk_3),
	.dataout({dataout_0}),
	.datain_l({\ac_2x_r~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_h(
	.clk(phy_clk_1x),
	.d(seq_ac_ba_1),
	.asdata(afi_ba_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_h~q ),
	.prn(vcc));
defparam ac_h.is_wysiwyg = "true";
defparam ac_h.power_up = "low";

dffeas ac_l(
	.clk(phy_clk_1x),
	.d(seq_ac_ba_4),
	.asdata(afi_ba_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_l~q ),
	.prn(vcc));
defparam ac_l.is_wysiwyg = "true";
defparam ac_l.power_up = "low";

dffeas ac_2x_r(
	.clk(clk_3),
	.d(\ac_2x_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_r~q ),
	.prn(vcc));
defparam ac_2x_r.is_wysiwyg = "true";
defparam ac_2x_r.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_3),
	.d(\ac_2x_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

dffeas ac_h_2r(
	.clk(clk_3),
	.d(\ac_h_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_2r~q ),
	.prn(vcc));
defparam ac_h_2r.is_wysiwyg = "true";
defparam ac_h_2r.power_up = "low";

dffeas ac_l_2r(
	.clk(clk_3),
	.d(\ac_l_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_2r~q ),
	.prn(vcc));
defparam ac_l_2r.is_wysiwyg = "true";
defparam ac_l_2r.power_up = "low";

arriaii_lcell_comb \ac_2x~0 (
	.dataa(!period_sel_addr_7),
	.datab(!\ac_h_2r~q ),
	.datac(!\ac_l_2r~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x~0 .extended_lut = "off";
defparam \ac_2x~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \ac_2x~0 .shared_arith = "off";

dffeas ac_1t(
	.clk(clk_3),
	.d(\ac_2x~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

arriaii_lcell_comb \ac_2x_r~0 (
	.dataa(!seq_ac_add_1t_ac_lat_internal),
	.datab(!\ac_2x~0_combout ),
	.datac(!\ac_1t~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x_r~0 .extended_lut = "off";
defparam \ac_2x_r~0 .lut_mask = 64'h2727272727272727;
defparam \ac_2x_r~0 .shared_arith = "off";

dffeas ac_h_r(
	.clk(phy_clk_1x),
	.d(\ac_h~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_r~q ),
	.prn(vcc));
defparam ac_h_r.is_wysiwyg = "true";
defparam ac_h_r.power_up = "low";

dffeas ac_l_r(
	.clk(phy_clk_1x),
	.d(\ac_l~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_r~q ),
	.prn(vcc));
defparam ac_l_r.is_wysiwyg = "true";
defparam ac_l_r.power_up = "low";

endmodule

module ddr3_int_altddio_out_16 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
inout 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_ddio_out_pgd_1 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module ddr3_int_ddio_out_pgd_1 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



arriaii_ddio_out \ddio_outa[0] (
	.datainlo(datain_l[0]),
	.datainhi(datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "clear";
defparam \ddio_outa[0] .power_up = "low";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_ac_16 (
	phy_clk_1x,
	clk_3,
	dataout_0,
	seq_ac_add_1t_ac_lat_internal,
	period_sel_addr_7,
	seq_ac_sel,
	afi_ba_2,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	phy_clk_1x;
input 	clk_3;
output 	dataout_0;
input 	seq_ac_add_1t_ac_lat_internal;
input 	period_sel_addr_7;
input 	seq_ac_sel;
input 	afi_ba_2;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ac_l~q ;
wire \ac_2x_r~q ;
wire \ac_2x_2r~q ;
wire \ac_h_2r~q ;
wire \ac_l_2r~q ;
wire \ac_2x~0_combout ;
wire \ac_1t~q ;
wire \ac_2x_r~0_combout ;
wire \ac_h_r~q ;
wire \ac_l_r~q ;


ddr3_int_altddio_out_17 \half_rate.addr_pin (
	.outclock(clk_3),
	.dataout({dataout_0}),
	.datain_l({\ac_2x_r~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_l(
	.clk(phy_clk_1x),
	.d(GND_port),
	.asdata(afi_ba_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_l~q ),
	.prn(vcc));
defparam ac_l.is_wysiwyg = "true";
defparam ac_l.power_up = "low";

dffeas ac_2x_r(
	.clk(clk_3),
	.d(\ac_2x_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_r~q ),
	.prn(vcc));
defparam ac_2x_r.is_wysiwyg = "true";
defparam ac_2x_r.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_3),
	.d(\ac_2x_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

dffeas ac_h_2r(
	.clk(clk_3),
	.d(\ac_h_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_2r~q ),
	.prn(vcc));
defparam ac_h_2r.is_wysiwyg = "true";
defparam ac_h_2r.power_up = "low";

dffeas ac_l_2r(
	.clk(clk_3),
	.d(\ac_l_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_2r~q ),
	.prn(vcc));
defparam ac_l_2r.is_wysiwyg = "true";
defparam ac_l_2r.power_up = "low";

arriaii_lcell_comb \ac_2x~0 (
	.dataa(!period_sel_addr_7),
	.datab(!\ac_h_2r~q ),
	.datac(!\ac_l_2r~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x~0 .extended_lut = "off";
defparam \ac_2x~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \ac_2x~0 .shared_arith = "off";

dffeas ac_1t(
	.clk(clk_3),
	.d(\ac_2x~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

arriaii_lcell_comb \ac_2x_r~0 (
	.dataa(!seq_ac_add_1t_ac_lat_internal),
	.datab(!\ac_2x~0_combout ),
	.datac(!\ac_1t~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x_r~0 .extended_lut = "off";
defparam \ac_2x_r~0 .lut_mask = 64'h2727272727272727;
defparam \ac_2x_r~0 .shared_arith = "off";

dffeas ac_h_r(
	.clk(phy_clk_1x),
	.d(\ac_l~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_r~q ),
	.prn(vcc));
defparam ac_h_r.is_wysiwyg = "true";
defparam ac_h_r.power_up = "low";

dffeas ac_l_r(
	.clk(phy_clk_1x),
	.d(\ac_l~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_r~q ),
	.prn(vcc));
defparam ac_l_r.is_wysiwyg = "true";
defparam ac_l_r.power_up = "low";

endmodule

module ddr3_int_altddio_out_17 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
inout 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_ddio_out_pgd_2 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module ddr3_int_ddio_out_pgd_2 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



arriaii_ddio_out \ddio_outa[0] (
	.datainlo(datain_l[0]),
	.datainhi(datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "clear";
defparam \ddio_outa[0] .power_up = "low";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_ac_17 (
	phy_clk_1x,
	clk_3,
	dataout_0,
	seq_ac_add_1t_ac_lat_internal,
	period_sel_addr_7,
	seq_ac_sel,
	afi_cas_n_0,
	seq_ac_cas_n_0,
	seq_ac_cas_n_1)/* synthesis synthesis_greybox=0 */;
input 	phy_clk_1x;
input 	clk_3;
output 	dataout_0;
input 	seq_ac_add_1t_ac_lat_internal;
input 	period_sel_addr_7;
input 	seq_ac_sel;
input 	afi_cas_n_0;
input 	seq_ac_cas_n_0;
input 	seq_ac_cas_n_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ac_h~q ;
wire \ac_l~q ;
wire \ac_2x_r~q ;
wire \ac_2x_2r~q ;
wire \ac_h_2r~q ;
wire \ac_l_2r~q ;
wire \ac_2x~0_combout ;
wire \ac_1t~q ;
wire \ac_2x_r~0_combout ;
wire \ac_h_r~q ;
wire \ac_l_r~q ;
wire \ac_h_r~0_combout ;
wire \ac_l_r~0_combout ;


ddr3_int_altddio_out_18 \half_rate.addr_pin (
	.outclock(clk_3),
	.dataout({dataout_0}),
	.datain_l({\ac_2x_r~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_h(
	.clk(phy_clk_1x),
	.d(seq_ac_cas_n_0),
	.asdata(afi_cas_n_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_h~q ),
	.prn(vcc));
defparam ac_h.is_wysiwyg = "true";
defparam ac_h.power_up = "low";

dffeas ac_l(
	.clk(phy_clk_1x),
	.d(seq_ac_cas_n_1),
	.asdata(afi_cas_n_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_l~q ),
	.prn(vcc));
defparam ac_l.is_wysiwyg = "true";
defparam ac_l.power_up = "low";

dffeas ac_2x_r(
	.clk(clk_3),
	.d(\ac_2x_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_r~q ),
	.prn(vcc));
defparam ac_2x_r.is_wysiwyg = "true";
defparam ac_2x_r.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_3),
	.d(\ac_2x_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

dffeas ac_h_2r(
	.clk(clk_3),
	.d(\ac_h_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_2r~q ),
	.prn(vcc));
defparam ac_h_2r.is_wysiwyg = "true";
defparam ac_h_2r.power_up = "low";

dffeas ac_l_2r(
	.clk(clk_3),
	.d(\ac_l_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_2r~q ),
	.prn(vcc));
defparam ac_l_2r.is_wysiwyg = "true";
defparam ac_l_2r.power_up = "low";

arriaii_lcell_comb \ac_2x~0 (
	.dataa(!period_sel_addr_7),
	.datab(!\ac_h_2r~q ),
	.datac(!\ac_l_2r~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x~0 .extended_lut = "off";
defparam \ac_2x~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \ac_2x~0 .shared_arith = "off";

dffeas ac_1t(
	.clk(clk_3),
	.d(\ac_2x~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

arriaii_lcell_comb \ac_2x_r~0 (
	.dataa(!seq_ac_add_1t_ac_lat_internal),
	.datab(!\ac_2x~0_combout ),
	.datac(!\ac_1t~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x_r~0 .extended_lut = "off";
defparam \ac_2x_r~0 .lut_mask = 64'h2727272727272727;
defparam \ac_2x_r~0 .shared_arith = "off";

dffeas ac_h_r(
	.clk(phy_clk_1x),
	.d(\ac_h_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_r~q ),
	.prn(vcc));
defparam ac_h_r.is_wysiwyg = "true";
defparam ac_h_r.power_up = "low";

dffeas ac_l_r(
	.clk(phy_clk_1x),
	.d(\ac_l_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_r~q ),
	.prn(vcc));
defparam ac_l_r.is_wysiwyg = "true";
defparam ac_l_r.power_up = "low";

arriaii_lcell_comb \ac_h_r~0 (
	.dataa(!\ac_h~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_h_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_h_r~0 .extended_lut = "off";
defparam \ac_h_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_h_r~0 .shared_arith = "off";

arriaii_lcell_comb \ac_l_r~0 (
	.dataa(!\ac_l~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_l_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_l_r~0 .extended_lut = "off";
defparam \ac_l_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_l_r~0 .shared_arith = "off";

endmodule

module ddr3_int_altddio_out_18 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
inout 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_ddio_out_6ed_14 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module ddr3_int_ddio_out_6ed_14 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



arriaii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_ac_18 (
	phy_clk_1x,
	clk_3,
	dataout_0,
	seq_ac_cke_1,
	ams_pipe_1,
	seq_ac_add_1t_ac_lat_internal,
	period_sel_addr_7,
	seq_ac_sel,
	int_cke_r_0)/* synthesis synthesis_greybox=0 */;
input 	phy_clk_1x;
input 	clk_3;
output 	dataout_0;
input 	seq_ac_cke_1;
input 	ams_pipe_1;
input 	seq_ac_add_1t_ac_lat_internal;
input 	period_sel_addr_7;
input 	seq_ac_sel;
input 	int_cke_r_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ac_h~q ;
wire \ac_l~q ;
wire \ac_2x_r~q ;
wire \ac_2x_2r~q ;
wire \ac_h_2r~q ;
wire \ac_l_2r~q ;
wire \ac_2x~0_combout ;
wire \ac_1t~q ;
wire \ac_2x_r~0_combout ;
wire \ac_h_r~q ;
wire \ac_l_r~q ;


ddr3_int_altddio_out_19 \half_rate.addr_pin (
	.outclock(clk_3),
	.dataout({dataout_0}),
	.aclr(ams_pipe_1),
	.datain_l({\ac_2x_r~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_h(
	.clk(phy_clk_1x),
	.d(seq_ac_cke_1),
	.asdata(int_cke_r_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_h~q ),
	.prn(vcc));
defparam ac_h.is_wysiwyg = "true";
defparam ac_h.power_up = "low";

dffeas ac_l(
	.clk(phy_clk_1x),
	.d(seq_ac_cke_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_l~q ),
	.prn(vcc));
defparam ac_l.is_wysiwyg = "true";
defparam ac_l.power_up = "low";

dffeas ac_2x_r(
	.clk(clk_3),
	.d(\ac_2x_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_r~q ),
	.prn(vcc));
defparam ac_2x_r.is_wysiwyg = "true";
defparam ac_2x_r.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_3),
	.d(\ac_2x_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

dffeas ac_h_2r(
	.clk(clk_3),
	.d(\ac_h_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_2r~q ),
	.prn(vcc));
defparam ac_h_2r.is_wysiwyg = "true";
defparam ac_h_2r.power_up = "low";

dffeas ac_l_2r(
	.clk(clk_3),
	.d(\ac_l_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_2r~q ),
	.prn(vcc));
defparam ac_l_2r.is_wysiwyg = "true";
defparam ac_l_2r.power_up = "low";

arriaii_lcell_comb \ac_2x~0 (
	.dataa(!period_sel_addr_7),
	.datab(!\ac_h_2r~q ),
	.datac(!\ac_l_2r~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x~0 .extended_lut = "off";
defparam \ac_2x~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \ac_2x~0 .shared_arith = "off";

dffeas ac_1t(
	.clk(clk_3),
	.d(\ac_2x~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

arriaii_lcell_comb \ac_2x_r~0 (
	.dataa(!seq_ac_add_1t_ac_lat_internal),
	.datab(!\ac_2x~0_combout ),
	.datac(!\ac_1t~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x_r~0 .extended_lut = "off";
defparam \ac_2x_r~0 .lut_mask = 64'h2727272727272727;
defparam \ac_2x_r~0 .shared_arith = "off";

dffeas ac_h_r(
	.clk(phy_clk_1x),
	.d(\ac_h~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_r~q ),
	.prn(vcc));
defparam ac_h_r.is_wysiwyg = "true";
defparam ac_h_r.power_up = "low";

dffeas ac_l_r(
	.clk(phy_clk_1x),
	.d(\ac_l~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_r~q ),
	.prn(vcc));
defparam ac_l_r.is_wysiwyg = "true";
defparam ac_l_r.power_up = "low";

endmodule

module ddr3_int_altddio_out_19 (
	outclock,
	dataout,
	aclr,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
inout 	[0:0] dataout;
input 	aclr;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_ddio_out_pgd_3 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.aclr(aclr),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module ddr3_int_ddio_out_pgd_3 (
	outclock,
	dataout,
	aclr,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
output 	[0:0] dataout;
input 	aclr;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



arriaii_ddio_out \ddio_outa[0] (
	.datainlo(datain_l[0]),
	.datainhi(datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(!aclr),
	.sreset(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "clear";
defparam \ddio_outa[0] .power_up = "low";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_ac_19 (
	phy_clk_1x,
	clk_3,
	dataout_0,
	ams_pipe_1,
	seq_ac_add_1t_ac_lat_internal,
	period_sel_addr_7,
	seq_ac_cs_n_0,
	seq_ac_sel,
	afi_cs_n_1,
	seq_ac_cs_n_1)/* synthesis synthesis_greybox=0 */;
input 	phy_clk_1x;
input 	clk_3;
output 	dataout_0;
input 	ams_pipe_1;
input 	seq_ac_add_1t_ac_lat_internal;
input 	period_sel_addr_7;
input 	seq_ac_cs_n_0;
input 	seq_ac_sel;
input 	afi_cs_n_1;
input 	seq_ac_cs_n_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ac_l~q ;
wire \ac_2x_r~q ;
wire \ac_2x_2r~q ;
wire \ac_h_2r~q ;
wire \ac_l_2r~q ;
wire \ac_2x~0_combout ;
wire \ac_1t~q ;
wire \ac_2x_r~0_combout ;
wire \ac_h_r~q ;
wire \ac_l_r~q ;
wire \ac_h~q ;
wire \ac_h~0_combout ;
wire \ac_h_r~0_combout ;
wire \ac_l_r~0_combout ;


ddr3_int_altddio_out_20 \half_rate.addr_pin (
	.outclock(clk_3),
	.dataout({dataout_0}),
	.datain_l({\ac_2x_r~q }),
	.datain_h({\ac_2x_2r~q }),
	.aset(ams_pipe_1));

dffeas ac_l(
	.clk(phy_clk_1x),
	.d(afi_cs_n_1),
	.asdata(seq_ac_cs_n_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!seq_ac_sel),
	.ena(vcc),
	.q(\ac_l~q ),
	.prn(vcc));
defparam ac_l.is_wysiwyg = "true";
defparam ac_l.power_up = "low";

dffeas ac_2x_r(
	.clk(clk_3),
	.d(\ac_2x_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_r~q ),
	.prn(vcc));
defparam ac_2x_r.is_wysiwyg = "true";
defparam ac_2x_r.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_3),
	.d(\ac_2x_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

dffeas ac_h_2r(
	.clk(clk_3),
	.d(\ac_h_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_2r~q ),
	.prn(vcc));
defparam ac_h_2r.is_wysiwyg = "true";
defparam ac_h_2r.power_up = "low";

dffeas ac_l_2r(
	.clk(clk_3),
	.d(\ac_l_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_2r~q ),
	.prn(vcc));
defparam ac_l_2r.is_wysiwyg = "true";
defparam ac_l_2r.power_up = "low";

arriaii_lcell_comb \ac_2x~0 (
	.dataa(!period_sel_addr_7),
	.datab(!\ac_h_2r~q ),
	.datac(!\ac_l_2r~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x~0 .extended_lut = "off";
defparam \ac_2x~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \ac_2x~0 .shared_arith = "off";

dffeas ac_1t(
	.clk(clk_3),
	.d(\ac_2x~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

arriaii_lcell_comb \ac_2x_r~0 (
	.dataa(!seq_ac_add_1t_ac_lat_internal),
	.datab(!\ac_2x~0_combout ),
	.datac(!\ac_1t~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x_r~0 .extended_lut = "off";
defparam \ac_2x_r~0 .lut_mask = 64'h2727272727272727;
defparam \ac_2x_r~0 .shared_arith = "off";

dffeas ac_h_r(
	.clk(phy_clk_1x),
	.d(\ac_h_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_r~q ),
	.prn(vcc));
defparam ac_h_r.is_wysiwyg = "true";
defparam ac_h_r.power_up = "low";

dffeas ac_l_r(
	.clk(phy_clk_1x),
	.d(\ac_l_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_r~q ),
	.prn(vcc));
defparam ac_l_r.is_wysiwyg = "true";
defparam ac_l_r.power_up = "low";

dffeas ac_h(
	.clk(phy_clk_1x),
	.d(\ac_h~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h~q ),
	.prn(vcc));
defparam ac_h.is_wysiwyg = "true";
defparam ac_h.power_up = "low";

arriaii_lcell_comb \ac_h~0 (
	.dataa(!seq_ac_cs_n_0),
	.datab(!seq_ac_sel),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_h~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_h~0 .extended_lut = "off";
defparam \ac_h~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \ac_h~0 .shared_arith = "off";

arriaii_lcell_comb \ac_h_r~0 (
	.dataa(!\ac_h~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_h_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_h_r~0 .extended_lut = "off";
defparam \ac_h_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_h_r~0 .shared_arith = "off";

arriaii_lcell_comb \ac_l_r~0 (
	.dataa(!\ac_l~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_l_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_l_r~0 .extended_lut = "off";
defparam \ac_l_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_l_r~0 .shared_arith = "off";

endmodule

module ddr3_int_altddio_out_20 (
	outclock,
	dataout,
	datain_l,
	datain_h,
	aset)/* synthesis synthesis_greybox=0 */;
input 	outclock;
inout 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;
input 	aset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_ddio_out_6ed_15 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}),
	.aset(aset));

endmodule

module ddr3_int_ddio_out_6ed_15 (
	outclock,
	dataout,
	datain_l,
	datain_h,
	aset)/* synthesis synthesis_greybox=0 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;
input 	aset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



arriaii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(!aset),
	.sreset(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_ac_20 (
	phy_clk_1x,
	clk_3,
	dataout_0,
	seq_ac_rst_n_0,
	ams_pipe_1,
	seq_ac_add_1t_ac_lat_internal,
	period_sel_addr_7,
	seq_ac_sel)/* synthesis synthesis_greybox=0 */;
input 	phy_clk_1x;
input 	clk_3;
output 	dataout_0;
input 	seq_ac_rst_n_0;
input 	ams_pipe_1;
input 	seq_ac_add_1t_ac_lat_internal;
input 	period_sel_addr_7;
input 	seq_ac_sel;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ac_2x_r~q ;
wire \ac_2x_2r~q ;
wire \ac_h_2r~q ;
wire \ac_l_2r~q ;
wire \ac_2x~0_combout ;
wire \ac_1t~q ;
wire \ac_2x_r~0_combout ;
wire \ac_h_r~q ;
wire \ac_l_r~q ;
wire \ac_h~q ;
wire \ac_h~0_combout ;


ddr3_int_altddio_out_21 \half_rate.addr_pin (
	.outclock(clk_3),
	.dataout({dataout_0}),
	.aclr(ams_pipe_1),
	.datain_l({\ac_2x_r~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_2x_r(
	.clk(clk_3),
	.d(\ac_2x_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_r~q ),
	.prn(vcc));
defparam ac_2x_r.is_wysiwyg = "true";
defparam ac_2x_r.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_3),
	.d(\ac_2x_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

dffeas ac_h_2r(
	.clk(clk_3),
	.d(\ac_h_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_2r~q ),
	.prn(vcc));
defparam ac_h_2r.is_wysiwyg = "true";
defparam ac_h_2r.power_up = "low";

dffeas ac_l_2r(
	.clk(clk_3),
	.d(\ac_l_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_2r~q ),
	.prn(vcc));
defparam ac_l_2r.is_wysiwyg = "true";
defparam ac_l_2r.power_up = "low";

arriaii_lcell_comb \ac_2x~0 (
	.dataa(!period_sel_addr_7),
	.datab(!\ac_h_2r~q ),
	.datac(!\ac_l_2r~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x~0 .extended_lut = "off";
defparam \ac_2x~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \ac_2x~0 .shared_arith = "off";

dffeas ac_1t(
	.clk(clk_3),
	.d(\ac_2x~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

arriaii_lcell_comb \ac_2x_r~0 (
	.dataa(!seq_ac_add_1t_ac_lat_internal),
	.datab(!\ac_2x~0_combout ),
	.datac(!\ac_1t~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x_r~0 .extended_lut = "off";
defparam \ac_2x_r~0 .lut_mask = 64'h2727272727272727;
defparam \ac_2x_r~0 .shared_arith = "off";

dffeas ac_h_r(
	.clk(phy_clk_1x),
	.d(\ac_h~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_r~q ),
	.prn(vcc));
defparam ac_h_r.is_wysiwyg = "true";
defparam ac_h_r.power_up = "low";

dffeas ac_l_r(
	.clk(phy_clk_1x),
	.d(\ac_h~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_r~q ),
	.prn(vcc));
defparam ac_l_r.is_wysiwyg = "true";
defparam ac_l_r.power_up = "low";

dffeas ac_h(
	.clk(phy_clk_1x),
	.d(\ac_h~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h~q ),
	.prn(vcc));
defparam ac_h.is_wysiwyg = "true";
defparam ac_h.power_up = "low";

arriaii_lcell_comb \ac_h~0 (
	.dataa(!seq_ac_sel),
	.datab(!seq_ac_rst_n_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_h~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_h~0 .extended_lut = "off";
defparam \ac_h~0 .lut_mask = 64'h7777777777777777;
defparam \ac_h~0 .shared_arith = "off";

endmodule

module ddr3_int_altddio_out_21 (
	outclock,
	dataout,
	aclr,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
inout 	[0:0] dataout;
input 	aclr;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_ddio_out_pgd_4 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.aclr(aclr),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module ddr3_int_ddio_out_pgd_4 (
	outclock,
	dataout,
	aclr,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
output 	[0:0] dataout;
input 	aclr;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



arriaii_ddio_out \ddio_outa[0] (
	.datainlo(datain_l[0]),
	.datainhi(datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(!aclr),
	.sreset(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "clear";
defparam \ddio_outa[0] .power_up = "low";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_ac_21 (
	phy_clk_1x,
	clk_3,
	dataout_0,
	seq_ac_add_1t_ac_lat_internal,
	period_sel_addr_7)/* synthesis synthesis_greybox=0 */;
input 	phy_clk_1x;
input 	clk_3;
output 	dataout_0;
input 	seq_ac_add_1t_ac_lat_internal;
input 	period_sel_addr_7;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ac_2x_r~q ;
wire \ac_2x_2r~q ;
wire \ac_h_2r~q ;
wire \ac_l_2r~q ;
wire \ac_2x~0_combout ;
wire \ac_1t~q ;
wire \ac_2x_r~0_combout ;
wire \ac_h_r~q ;
wire \ac_l_r~q ;
wire \ac_h_r~0_combout ;
wire \ac_l_r~0_combout ;


ddr3_int_altddio_out_22 \half_rate.addr_pin (
	.outclock(clk_3),
	.dataout({dataout_0}),
	.datain_l({\ac_2x_r~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_2x_r(
	.clk(clk_3),
	.d(\ac_2x_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_r~q ),
	.prn(vcc));
defparam ac_2x_r.is_wysiwyg = "true";
defparam ac_2x_r.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_3),
	.d(\ac_2x_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

dffeas ac_h_2r(
	.clk(clk_3),
	.d(\ac_h_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_2r~q ),
	.prn(vcc));
defparam ac_h_2r.is_wysiwyg = "true";
defparam ac_h_2r.power_up = "low";

dffeas ac_l_2r(
	.clk(clk_3),
	.d(\ac_l_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_2r~q ),
	.prn(vcc));
defparam ac_l_2r.is_wysiwyg = "true";
defparam ac_l_2r.power_up = "low";

arriaii_lcell_comb \ac_2x~0 (
	.dataa(!period_sel_addr_7),
	.datab(!\ac_h_2r~q ),
	.datac(!\ac_l_2r~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x~0 .extended_lut = "off";
defparam \ac_2x~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \ac_2x~0 .shared_arith = "off";

dffeas ac_1t(
	.clk(clk_3),
	.d(\ac_2x~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

arriaii_lcell_comb \ac_2x_r~0 (
	.dataa(!seq_ac_add_1t_ac_lat_internal),
	.datab(!\ac_2x~0_combout ),
	.datac(!\ac_1t~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x_r~0 .extended_lut = "off";
defparam \ac_2x_r~0 .lut_mask = 64'h2727272727272727;
defparam \ac_2x_r~0 .shared_arith = "off";

dffeas ac_h_r(
	.clk(phy_clk_1x),
	.d(\ac_h_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_r~q ),
	.prn(vcc));
defparam ac_h_r.is_wysiwyg = "true";
defparam ac_h_r.power_up = "low";

dffeas ac_l_r(
	.clk(phy_clk_1x),
	.d(\ac_l_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_r~q ),
	.prn(vcc));
defparam ac_l_r.is_wysiwyg = "true";
defparam ac_l_r.power_up = "low";

arriaii_lcell_comb \ac_h_r~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_h_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_h_r~0 .extended_lut = "off";
defparam \ac_h_r~0 .lut_mask = 64'h0000000000000000;
defparam \ac_h_r~0 .shared_arith = "off";

arriaii_lcell_comb \ac_l_r~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_l_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_l_r~0 .extended_lut = "off";
defparam \ac_l_r~0 .lut_mask = 64'h0000000000000000;
defparam \ac_l_r~0 .shared_arith = "off";

endmodule

module ddr3_int_altddio_out_22 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
inout 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_ddio_out_pgd_5 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module ddr3_int_ddio_out_pgd_5 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



arriaii_ddio_out \ddio_outa[0] (
	.datainlo(datain_l[0]),
	.datainhi(datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "clear";
defparam \ddio_outa[0] .power_up = "low";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_ac_22 (
	phy_clk_1x,
	clk_3,
	dataout_0,
	seq_ac_add_1t_ac_lat_internal,
	period_sel_addr_7,
	seq_ac_sel,
	afi_ras_n_0,
	seq_ac_ras_n_0,
	seq_ac_ras_n_1)/* synthesis synthesis_greybox=0 */;
input 	phy_clk_1x;
input 	clk_3;
output 	dataout_0;
input 	seq_ac_add_1t_ac_lat_internal;
input 	period_sel_addr_7;
input 	seq_ac_sel;
input 	afi_ras_n_0;
input 	seq_ac_ras_n_0;
input 	seq_ac_ras_n_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ac_h~q ;
wire \ac_l~q ;
wire \ac_2x_r~q ;
wire \ac_2x_2r~q ;
wire \ac_h_2r~q ;
wire \ac_l_2r~q ;
wire \ac_2x~0_combout ;
wire \ac_1t~q ;
wire \ac_2x_r~0_combout ;
wire \ac_h_r~q ;
wire \ac_l_r~q ;
wire \ac_h_r~0_combout ;
wire \ac_l_r~0_combout ;


ddr3_int_altddio_out_23 \half_rate.addr_pin (
	.outclock(clk_3),
	.dataout({dataout_0}),
	.datain_l({\ac_2x_r~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_h(
	.clk(phy_clk_1x),
	.d(seq_ac_ras_n_0),
	.asdata(afi_ras_n_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_h~q ),
	.prn(vcc));
defparam ac_h.is_wysiwyg = "true";
defparam ac_h.power_up = "low";

dffeas ac_l(
	.clk(phy_clk_1x),
	.d(seq_ac_ras_n_1),
	.asdata(afi_ras_n_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_l~q ),
	.prn(vcc));
defparam ac_l.is_wysiwyg = "true";
defparam ac_l.power_up = "low";

dffeas ac_2x_r(
	.clk(clk_3),
	.d(\ac_2x_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_r~q ),
	.prn(vcc));
defparam ac_2x_r.is_wysiwyg = "true";
defparam ac_2x_r.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_3),
	.d(\ac_2x_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

dffeas ac_h_2r(
	.clk(clk_3),
	.d(\ac_h_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_2r~q ),
	.prn(vcc));
defparam ac_h_2r.is_wysiwyg = "true";
defparam ac_h_2r.power_up = "low";

dffeas ac_l_2r(
	.clk(clk_3),
	.d(\ac_l_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_2r~q ),
	.prn(vcc));
defparam ac_l_2r.is_wysiwyg = "true";
defparam ac_l_2r.power_up = "low";

arriaii_lcell_comb \ac_2x~0 (
	.dataa(!period_sel_addr_7),
	.datab(!\ac_h_2r~q ),
	.datac(!\ac_l_2r~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x~0 .extended_lut = "off";
defparam \ac_2x~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \ac_2x~0 .shared_arith = "off";

dffeas ac_1t(
	.clk(clk_3),
	.d(\ac_2x~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

arriaii_lcell_comb \ac_2x_r~0 (
	.dataa(!seq_ac_add_1t_ac_lat_internal),
	.datab(!\ac_2x~0_combout ),
	.datac(!\ac_1t~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x_r~0 .extended_lut = "off";
defparam \ac_2x_r~0 .lut_mask = 64'h2727272727272727;
defparam \ac_2x_r~0 .shared_arith = "off";

dffeas ac_h_r(
	.clk(phy_clk_1x),
	.d(\ac_h_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_r~q ),
	.prn(vcc));
defparam ac_h_r.is_wysiwyg = "true";
defparam ac_h_r.power_up = "low";

dffeas ac_l_r(
	.clk(phy_clk_1x),
	.d(\ac_l_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_r~q ),
	.prn(vcc));
defparam ac_l_r.is_wysiwyg = "true";
defparam ac_l_r.power_up = "low";

arriaii_lcell_comb \ac_h_r~0 (
	.dataa(!\ac_h~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_h_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_h_r~0 .extended_lut = "off";
defparam \ac_h_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_h_r~0 .shared_arith = "off";

arriaii_lcell_comb \ac_l_r~0 (
	.dataa(!\ac_l~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_l_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_l_r~0 .extended_lut = "off";
defparam \ac_l_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_l_r~0 .shared_arith = "off";

endmodule

module ddr3_int_altddio_out_23 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
inout 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_ddio_out_6ed_16 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module ddr3_int_ddio_out_6ed_16 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



arriaii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_ac_23 (
	phy_clk_1x,
	clk_3,
	dataout_0,
	seq_ac_add_1t_ac_lat_internal,
	period_sel_addr_7,
	seq_ac_sel,
	afi_we_n_0,
	seq_ac_we_n_0,
	seq_ac_we_n_1)/* synthesis synthesis_greybox=0 */;
input 	phy_clk_1x;
input 	clk_3;
output 	dataout_0;
input 	seq_ac_add_1t_ac_lat_internal;
input 	period_sel_addr_7;
input 	seq_ac_sel;
input 	afi_we_n_0;
input 	seq_ac_we_n_0;
input 	seq_ac_we_n_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ac_h~q ;
wire \ac_l~q ;
wire \ac_2x_r~q ;
wire \ac_2x_2r~q ;
wire \ac_h_2r~q ;
wire \ac_l_2r~q ;
wire \ac_2x~0_combout ;
wire \ac_1t~q ;
wire \ac_2x_r~0_combout ;
wire \ac_h_r~q ;
wire \ac_l_r~q ;
wire \ac_h_r~0_combout ;
wire \ac_l_r~0_combout ;


ddr3_int_altddio_out_24 \half_rate.addr_pin (
	.outclock(clk_3),
	.dataout({dataout_0}),
	.datain_l({\ac_2x_r~q }),
	.datain_h({\ac_2x_2r~q }));

dffeas ac_h(
	.clk(phy_clk_1x),
	.d(seq_ac_we_n_0),
	.asdata(afi_we_n_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_h~q ),
	.prn(vcc));
defparam ac_h.is_wysiwyg = "true";
defparam ac_h.power_up = "low";

dffeas ac_l(
	.clk(phy_clk_1x),
	.d(seq_ac_we_n_1),
	.asdata(afi_we_n_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_ac_sel),
	.ena(vcc),
	.q(\ac_l~q ),
	.prn(vcc));
defparam ac_l.is_wysiwyg = "true";
defparam ac_l.power_up = "low";

dffeas ac_2x_r(
	.clk(clk_3),
	.d(\ac_2x_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_r~q ),
	.prn(vcc));
defparam ac_2x_r.is_wysiwyg = "true";
defparam ac_2x_r.power_up = "low";

dffeas ac_2x_2r(
	.clk(clk_3),
	.d(\ac_2x_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_2x_2r~q ),
	.prn(vcc));
defparam ac_2x_2r.is_wysiwyg = "true";
defparam ac_2x_2r.power_up = "low";

dffeas ac_h_2r(
	.clk(clk_3),
	.d(\ac_h_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_2r~q ),
	.prn(vcc));
defparam ac_h_2r.is_wysiwyg = "true";
defparam ac_h_2r.power_up = "low";

dffeas ac_l_2r(
	.clk(clk_3),
	.d(\ac_l_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_2r~q ),
	.prn(vcc));
defparam ac_l_2r.is_wysiwyg = "true";
defparam ac_l_2r.power_up = "low";

arriaii_lcell_comb \ac_2x~0 (
	.dataa(!period_sel_addr_7),
	.datab(!\ac_h_2r~q ),
	.datac(!\ac_l_2r~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x~0 .extended_lut = "off";
defparam \ac_2x~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \ac_2x~0 .shared_arith = "off";

dffeas ac_1t(
	.clk(clk_3),
	.d(\ac_2x~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_1t~q ),
	.prn(vcc));
defparam ac_1t.is_wysiwyg = "true";
defparam ac_1t.power_up = "low";

arriaii_lcell_comb \ac_2x_r~0 (
	.dataa(!seq_ac_add_1t_ac_lat_internal),
	.datab(!\ac_2x~0_combout ),
	.datac(!\ac_1t~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_2x_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_2x_r~0 .extended_lut = "off";
defparam \ac_2x_r~0 .lut_mask = 64'h2727272727272727;
defparam \ac_2x_r~0 .shared_arith = "off";

dffeas ac_h_r(
	.clk(phy_clk_1x),
	.d(\ac_h_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_h_r~q ),
	.prn(vcc));
defparam ac_h_r.is_wysiwyg = "true";
defparam ac_h_r.power_up = "low";

dffeas ac_l_r(
	.clk(phy_clk_1x),
	.d(\ac_l_r~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_l_r~q ),
	.prn(vcc));
defparam ac_l_r.is_wysiwyg = "true";
defparam ac_l_r.power_up = "low";

arriaii_lcell_comb \ac_h_r~0 (
	.dataa(!\ac_h~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_h_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_h_r~0 .extended_lut = "off";
defparam \ac_h_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_h_r~0 .shared_arith = "off";

arriaii_lcell_comb \ac_l_r~0 (
	.dataa(!\ac_l~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_l_r~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_l_r~0 .extended_lut = "off";
defparam \ac_l_r~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ac_l_r~0 .shared_arith = "off";

endmodule

module ddr3_int_altddio_out_24 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
inout 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_ddio_out_6ed_17 auto_generated(
	.outclock(outclock),
	.dataout({dataout[0]}),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}));

endmodule

module ddr3_int_ddio_out_6ed_17 (
	outclock,
	dataout,
	datain_l,
	datain_h)/* synthesis synthesis_greybox=0 */;
input 	outclock;
output 	[0:0] dataout;
input 	[0:0] datain_l;
input 	[0:0] datain_h;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



arriaii_ddio_out \ddio_outa[0] (
	.datainlo(!datain_l[0]),
	.datainhi(!datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "preset";
defparam \ddio_outa[0] .power_up = "high";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_clk_reset (
	clk_0,
	clk_1,
	clk_3,
	clk_4,
	clk_5,
	dqs_delay_ctrl,
	mem_clk_buf_in_0,
	mem_clk_n_buf_in_0,
	mimic_data_2x,
	fb_clk,
	reset_request_n,
	reset_phy_clk_1x_n1,
	ams_pipe_1,
	ams_pipe_11,
	ams_pipe_12,
	seq_rdp_reset_req_n,
	seq_pll_inc_dec_n,
	seq_pll_start_reconfig,
	ams_pipe_3,
	seq_pll_select,
	seq_mem_clk_disable,
	ams_pipe_31,
	ams_pipe_13,
	phs_shft_busy_siii1,
	global_reset_n,
	pll_ref_clk,
	soft_reset_n)/* synthesis synthesis_greybox=0 */;
output 	clk_0;
output 	clk_1;
output 	clk_3;
output 	clk_4;
output 	clk_5;
output 	[5:0] dqs_delay_ctrl;
output 	mem_clk_buf_in_0;
output 	mem_clk_n_buf_in_0;
output 	mimic_data_2x;
input 	fb_clk;
output 	reset_request_n;
output 	reset_phy_clk_1x_n1;
output 	ams_pipe_1;
output 	ams_pipe_11;
output 	ams_pipe_12;
input 	seq_rdp_reset_req_n;
input 	seq_pll_inc_dec_n;
input 	seq_pll_start_reconfig;
output 	ams_pipe_3;
input 	[2:0] seq_pll_select;
input 	seq_mem_clk_disable;
output 	ams_pipe_31;
output 	ams_pipe_13;
output 	phs_shft_busy_siii1;
input 	global_reset_n;
input 	pll_ref_clk;
input 	soft_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \half_rate.pll|altpll_component|auto_generated|phasedone ;
wire \half_rate.pll|altpll_component|auto_generated|pll1~LOCKED ;
wire \dll~UPNDNOUT ;
wire \half_rate.pll|altpll_component|auto_generated|pll_lock_sync~q ;
wire \pll_new_dir~q ;
wire \comb~0_combout ;
wire \seq_pll_inc_dec_ccd~q ;
wire \pll_reprogram_request_pulse_2r~q ;
wire \pll_new_phase[2]~q ;
wire \pll_new_phase[1]~q ;
wire \pll_new_phase[0]~q ;
wire \poa_clk_pipe|ams_pipe[0]~q ;
wire \always3~0_combout ;
wire \seq_pll_select_ccd[2]~q ;
wire \seq_pll_select_ccd[1]~q ;
wire \seq_pll_select_ccd[0]~q ;
wire \mem_clk_pdiff_in[0] ;
wire \phy_internal_reset_n~combout ;
wire \reset_master_ams~q ;
wire \global_pre_clear~q ;
wire \divider[1]~2_combout ;
wire \pll_reconfig_reset_n~0_combout ;
wire \clk_div_reset_ams_n~q ;
wire \clk_div_reset_ams_n_r~q ;
wire \divider[1]~q ;
wire \divider[2]~1_combout ;
wire \divider[2]~q ;
wire \divider~0_combout ;
wire \divider[0]~q ;
wire \scan_clk~0_combout ;
wire \scan_clk~q ;
wire \seq_pll_start_reconfig_ccd_pipe[0]~q ;
wire \seq_pll_start_reconfig_ccd_pipe[1]~q ;
wire \seq_pll_start_reconfig_ccd_pipe[2]~q ;
wire \pll_reconfig_reset_ams_n~q ;
wire \pll_reconfig_reset_ams_n_r~q ;
wire \seq_pll_start_reconfig_ams~q ;
wire \seq_pll_start_reconfig_r~q ;
wire \seq_pll_start_reconfig_2r~q ;
wire \seq_pll_start_reconfig_3r~q ;
wire \pll_phase_auto_calibrate_pulse~combout ;
wire \pll_reprogram_request_pulse~q ;
wire \pll_reprogram_request_pulse_r~q ;
wire \pll_reprogram_request_long_pulse~combout ;
wire \pll_reprogram_request~q ;
wire \phs_shft_busy_siii~0_combout ;

wire [5:0] dll_DELAYCTRLOUT_bus;

assign dqs_delay_ctrl[0] = dll_DELAYCTRLOUT_bus[0];
assign dqs_delay_ctrl[1] = dll_DELAYCTRLOUT_bus[1];
assign dqs_delay_ctrl[2] = dll_DELAYCTRLOUT_bus[2];
assign dqs_delay_ctrl[3] = dll_DELAYCTRLOUT_bus[3];
assign dqs_delay_ctrl[4] = dll_DELAYCTRLOUT_bus[4];
assign dqs_delay_ctrl[5] = dll_DELAYCTRLOUT_bus[5];

ddr3_int_ddr3_int_phy_alt_mem_phy_pll \half_rate.pll (
	.phasedone(\half_rate.pll|altpll_component|auto_generated|phasedone ),
	.pll1(\half_rate.pll|altpll_component|auto_generated|pll1~LOCKED ),
	.clk_0(clk_0),
	.clk_1(clk_1),
	.clk_3(clk_3),
	.clk_4(clk_4),
	.clk_5(clk_5),
	.pll_lock_sync(\half_rate.pll|altpll_component|auto_generated|pll_lock_sync~q ),
	.locked(reset_request_n),
	.pll_new_dir(\pll_new_dir~q ),
	.pll_reprogram_request(\pll_reprogram_request~q ),
	.scan_clk(\scan_clk~q ),
	.pll_new_phase_2(\pll_new_phase[2]~q ),
	.pll_new_phase_1(\pll_new_phase[1]~q ),
	.pll_new_phase_0(\pll_new_phase[0]~q ),
	.global_reset_n(global_reset_n),
	.pll_ref_clk(pll_ref_clk));

ddr3_int_ddr3_int_phy_alt_mem_phy_reset_pipe_6 reset_rdp_phy_clk_pipe(
	.clock(clk_0),
	.ams_pipe_1(ams_pipe_1),
	.pre_clear(\comb~0_combout ));

ddr3_int_ddr3_int_phy_alt_mem_phy_reset_pipe_3 mem_clk_pipe(
	.clock(clk_1),
	.pre_clear(\global_pre_clear~q ),
	.ams_pipe_3(ams_pipe_31));

ddr3_int_ddr3_int_phy_alt_mem_phy_reset_pipe_5 poa_clk_pipe(
	.clock(clk_4),
	.pre_clear(\comb~0_combout ),
	.ams_pipe_0(\poa_clk_pipe|ams_pipe[0]~q ));

ddr3_int_ddr3_int_phy_alt_mem_phy_reset_pipe_8 write_clk_pipe(
	.clock(clk_3),
	.ams_pipe_1(ams_pipe_11),
	.pre_clear(\global_pre_clear~q ),
	.ams_pipe_3(ams_pipe_3));

ddr3_int_ddr3_int_phy_alt_mem_phy_reset_pipe ac_clk_pipe_2x(
	.clock(clk_3),
	.ams_pipe_1(ams_pipe_11),
	.pre_clear(\global_pre_clear~q ));

ddr3_int_ddr3_int_phy_alt_mem_phy_reset_pipe_2 measure_clk_pipe(
	.clock(clk_5),
	.pre_clear(\global_pre_clear~q ),
	.ams_pipe_1(ams_pipe_13));

ddr3_int_ddr3_int_phy_alt_mem_phy_reset_pipe_7 resync_clk_2x_pipe(
	.clock(clk_4),
	.ams_pipe_1(ams_pipe_12),
	.pre_clear(\comb~0_combout ),
	.ams_pipe_0(\poa_clk_pipe|ams_pipe[0]~q ));

dffeas pll_new_dir(
	.clk(\scan_clk~q ),
	.d(\seq_pll_inc_dec_ccd~q ),
	.asdata(vcc),
	.clrn(\pll_reconfig_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pll_phase_auto_calibrate_pulse~combout ),
	.q(\pll_new_dir~q ),
	.prn(vcc));
defparam pll_new_dir.is_wysiwyg = "true";
defparam pll_new_dir.power_up = "low";

arriaii_lcell_comb \comb~0 (
	.dataa(!\global_pre_clear~q ),
	.datab(!seq_rdp_reset_req_n),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\comb~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~0 .extended_lut = "off";
defparam \comb~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \comb~0 .shared_arith = "off";

dffeas seq_pll_inc_dec_ccd(
	.clk(clk_0),
	.d(seq_pll_inc_dec_n),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\seq_pll_inc_dec_ccd~q ),
	.prn(vcc));
defparam seq_pll_inc_dec_ccd.is_wysiwyg = "true";
defparam seq_pll_inc_dec_ccd.power_up = "low";

dffeas pll_reprogram_request_pulse_2r(
	.clk(\scan_clk~q ),
	.d(\pll_reprogram_request_pulse_r~q ),
	.asdata(vcc),
	.clrn(\pll_reconfig_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pll_reprogram_request_pulse_2r~q ),
	.prn(vcc));
defparam pll_reprogram_request_pulse_2r.is_wysiwyg = "true";
defparam pll_reprogram_request_pulse_2r.power_up = "low";

dffeas \pll_new_phase[2] (
	.clk(\scan_clk~q ),
	.d(\seq_pll_select_ccd[2]~q ),
	.asdata(vcc),
	.clrn(\pll_reconfig_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pll_phase_auto_calibrate_pulse~combout ),
	.q(\pll_new_phase[2]~q ),
	.prn(vcc));
defparam \pll_new_phase[2] .is_wysiwyg = "true";
defparam \pll_new_phase[2] .power_up = "low";

dffeas \pll_new_phase[1] (
	.clk(\scan_clk~q ),
	.d(\seq_pll_select_ccd[1]~q ),
	.asdata(vcc),
	.clrn(\pll_reconfig_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pll_phase_auto_calibrate_pulse~combout ),
	.q(\pll_new_phase[1]~q ),
	.prn(vcc));
defparam \pll_new_phase[1] .is_wysiwyg = "true";
defparam \pll_new_phase[1] .power_up = "low";

dffeas \pll_new_phase[0] (
	.clk(\scan_clk~q ),
	.d(\seq_pll_select_ccd[0]~q ),
	.asdata(vcc),
	.clrn(\pll_reconfig_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pll_phase_auto_calibrate_pulse~combout ),
	.q(\pll_new_phase[0]~q ),
	.prn(vcc));
defparam \pll_new_phase[0] .is_wysiwyg = "true";
defparam \pll_new_phase[0] .power_up = "low";

arriaii_lcell_comb \always3~0 (
	.dataa(!seq_pll_start_reconfig),
	.datab(!\seq_pll_start_reconfig_ccd_pipe[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always3~0 .extended_lut = "off";
defparam \always3~0 .lut_mask = 64'h4444444444444444;
defparam \always3~0 .shared_arith = "off";

dffeas \seq_pll_select_ccd[2] (
	.clk(clk_0),
	.d(seq_pll_select[0]),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\seq_pll_select_ccd[2]~q ),
	.prn(vcc));
defparam \seq_pll_select_ccd[2] .is_wysiwyg = "true";
defparam \seq_pll_select_ccd[2] .power_up = "low";

dffeas \seq_pll_select_ccd[1] (
	.clk(clk_0),
	.d(seq_pll_select[1]),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\seq_pll_select_ccd[1]~q ),
	.prn(vcc));
defparam \seq_pll_select_ccd[1] .is_wysiwyg = "true";
defparam \seq_pll_select_ccd[1] .power_up = "low";

dffeas \seq_pll_select_ccd[0] (
	.clk(clk_0),
	.d(seq_pll_select[0]),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always3~0_combout ),
	.q(\seq_pll_select_ccd[0]~q ),
	.prn(vcc));
defparam \seq_pll_select_ccd[0] .is_wysiwyg = "true";
defparam \seq_pll_select_ccd[0] .power_up = "low";

arriaii_dll dll(
	.clk(clk_1),
	.aload(reset_request_n),
	.upndnin(vcc),
	.upndninclkena(vcc),
	.dqsupdate(),
	.upndnout(\dll~UPNDNOUT ),
	.offsetdelayctrlclkout(),
	.offsetdelayctrlout(),
	.delayctrlout(dll_DELAYCTRLOUT_bus));
defparam dll.delay_buffer_mode = "high";
defparam dll.delay_chain_length = 10;
defparam dll.delayctrlout_mode = "normal";
defparam dll.dual_phase_comparators = "true";
defparam dll.input_frequency = "3333ps";
defparam dll.jitter_reduction = "true";
defparam dll.sim_buffer_delay_increment = 10;
defparam dll.sim_high_buffer_intrinsic_delay = 175;
defparam dll.sim_low_buffer_intrinsic_delay = 350;
defparam dll.sim_valid_lock = 1280;
defparam dll.sim_valid_lockcount = 0;
defparam dll.static_delay_ctrl = 0;
defparam dll.use_upndnin = "false";
defparam dll.use_upndninclkena = "false";

arriaii_pseudo_diff_out \DDR_CLK_OUT[0].mem_clk_pdiff (
	.i(\mem_clk_pdiff_in[0] ),
	.o(mem_clk_buf_in_0),
	.obar(mem_clk_n_buf_in_0));

arriaii_ddio_in ddio_mimic(
	.datain(fb_clk),
	.clk(clk_5),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(),
	.regouthi(mimic_data_2x),
	.dfflo());
defparam ddio_mimic.async_mode = "none";
defparam ddio_mimic.power_up = "low";
defparam ddio_mimic.sync_mode = "none";
defparam ddio_mimic.use_clkn = "false";

dffeas reset_phy_clk_1x_n(
	.clk(clk_0),
	.d(vcc),
	.asdata(vcc),
	.clrn(\global_pre_clear~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(reset_phy_clk_1x_n1),
	.prn(vcc));
defparam reset_phy_clk_1x_n.is_wysiwyg = "true";
defparam reset_phy_clk_1x_n.power_up = "low";

dffeas phs_shft_busy_siii(
	.clk(\scan_clk~q ),
	.d(\phs_shft_busy_siii~0_combout ),
	.asdata(vcc),
	.clrn(\pll_reconfig_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(phs_shft_busy_siii1),
	.prn(vcc));
defparam phs_shft_busy_siii.is_wysiwyg = "true";
defparam phs_shft_busy_siii.power_up = "low";

arriaii_ddio_out \DDR_CLK_OUT[0].mem_clk_ddio (
	.datainlo(gnd),
	.datainhi(vcc),
	.clkhi(clk_1),
	.clklo(clk_1),
	.muxsel(clk_1),
	.ena(vcc),
	.areset(gnd),
	.sreset(!seq_mem_clk_disable),
	.clk(gnd),
	.dataout(\mem_clk_pdiff_in[0] ),
	.dfflo(),
	.dffhi());
defparam \DDR_CLK_OUT[0].mem_clk_ddio .async_mode = "none";
defparam \DDR_CLK_OUT[0].mem_clk_ddio .power_up = "low";
defparam \DDR_CLK_OUT[0].mem_clk_ddio .sync_mode = "clear";
defparam \DDR_CLK_OUT[0].mem_clk_ddio .use_new_clocking_model = "true";

arriaii_lcell_comb phy_internal_reset_n(
	.dataa(!\half_rate.pll|altpll_component|auto_generated|pll1~LOCKED ),
	.datab(!\half_rate.pll|altpll_component|auto_generated|pll_lock_sync~q ),
	.datac(!global_reset_n),
	.datad(!soft_reset_n),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\phy_internal_reset_n~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam phy_internal_reset_n.extended_lut = "off";
defparam phy_internal_reset_n.lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam phy_internal_reset_n.shared_arith = "off";

dffeas reset_master_ams(
	.clk(clk_0),
	.d(vcc),
	.asdata(vcc),
	.clrn(!\phy_internal_reset_n~combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\reset_master_ams~q ),
	.prn(vcc));
defparam reset_master_ams.is_wysiwyg = "true";
defparam reset_master_ams.power_up = "low";

dffeas global_pre_clear(
	.clk(clk_0),
	.d(\reset_master_ams~q ),
	.asdata(vcc),
	.clrn(!\phy_internal_reset_n~combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\global_pre_clear~q ),
	.prn(vcc));
defparam global_pre_clear.is_wysiwyg = "true";
defparam global_pre_clear.power_up = "low";

arriaii_lcell_comb \divider[1]~2 (
	.dataa(!\divider[0]~q ),
	.datab(!\divider[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\divider[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \divider[1]~2 .extended_lut = "off";
defparam \divider[1]~2 .lut_mask = 64'h6666666666666666;
defparam \divider[1]~2 .shared_arith = "off";

arriaii_lcell_comb \pll_reconfig_reset_n~0 (
	.dataa(!\half_rate.pll|altpll_component|auto_generated|pll1~LOCKED ),
	.datab(!\half_rate.pll|altpll_component|auto_generated|pll_lock_sync~q ),
	.datac(!global_reset_n),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pll_reconfig_reset_n~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pll_reconfig_reset_n~0 .extended_lut = "off";
defparam \pll_reconfig_reset_n~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \pll_reconfig_reset_n~0 .shared_arith = "off";

dffeas clk_div_reset_ams_n(
	.clk(clk_0),
	.d(vcc),
	.asdata(vcc),
	.clrn(!\pll_reconfig_reset_n~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\clk_div_reset_ams_n~q ),
	.prn(vcc));
defparam clk_div_reset_ams_n.is_wysiwyg = "true";
defparam clk_div_reset_ams_n.power_up = "low";

dffeas clk_div_reset_ams_n_r(
	.clk(clk_0),
	.d(\clk_div_reset_ams_n~q ),
	.asdata(vcc),
	.clrn(!\pll_reconfig_reset_n~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\clk_div_reset_ams_n_r~q ),
	.prn(vcc));
defparam clk_div_reset_ams_n_r.is_wysiwyg = "true";
defparam clk_div_reset_ams_n_r.power_up = "low";

dffeas \divider[1] (
	.clk(clk_0),
	.d(\divider[1]~2_combout ),
	.asdata(vcc),
	.clrn(\clk_div_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\divider[1]~q ),
	.prn(vcc));
defparam \divider[1] .is_wysiwyg = "true";
defparam \divider[1] .power_up = "low";

arriaii_lcell_comb \divider[2]~1 (
	.dataa(!\divider[0]~q ),
	.datab(!\divider[2]~q ),
	.datac(!\divider[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\divider[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \divider[2]~1 .extended_lut = "off";
defparam \divider[2]~1 .lut_mask = 64'h3636363636363636;
defparam \divider[2]~1 .shared_arith = "off";

dffeas \divider[2] (
	.clk(clk_0),
	.d(\divider[2]~1_combout ),
	.asdata(vcc),
	.clrn(\clk_div_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\divider[2]~q ),
	.prn(vcc));
defparam \divider[2] .is_wysiwyg = "true";
defparam \divider[2] .power_up = "low";

arriaii_lcell_comb \divider~0 (
	.dataa(!\divider[0]~q ),
	.datab(!\divider[2]~q ),
	.datac(!\divider[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\divider~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \divider~0 .extended_lut = "off";
defparam \divider~0 .lut_mask = 64'h2A2A2A2A2A2A2A2A;
defparam \divider~0 .shared_arith = "off";

dffeas \divider[0] (
	.clk(clk_0),
	.d(\divider~0_combout ),
	.asdata(vcc),
	.clrn(\clk_div_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\divider[0]~q ),
	.prn(vcc));
defparam \divider[0] .is_wysiwyg = "true";
defparam \divider[0] .power_up = "low";

arriaii_lcell_comb \scan_clk~0 (
	.dataa(!\scan_clk~q ),
	.datab(!\divider[0]~q ),
	.datac(!\divider[2]~q ),
	.datad(!\divider[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\scan_clk~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \scan_clk~0 .extended_lut = "off";
defparam \scan_clk~0 .lut_mask = 64'h9555955595559555;
defparam \scan_clk~0 .shared_arith = "off";

dffeas scan_clk(
	.clk(clk_0),
	.d(\scan_clk~0_combout ),
	.asdata(vcc),
	.clrn(\clk_div_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\scan_clk~q ),
	.prn(vcc));
defparam scan_clk.is_wysiwyg = "true";
defparam scan_clk.power_up = "low";

dffeas \seq_pll_start_reconfig_ccd_pipe[0] (
	.clk(clk_0),
	.d(seq_pll_start_reconfig),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_pll_start_reconfig_ccd_pipe[0]~q ),
	.prn(vcc));
defparam \seq_pll_start_reconfig_ccd_pipe[0] .is_wysiwyg = "true";
defparam \seq_pll_start_reconfig_ccd_pipe[0] .power_up = "low";

dffeas \seq_pll_start_reconfig_ccd_pipe[1] (
	.clk(clk_0),
	.d(\seq_pll_start_reconfig_ccd_pipe[0]~q ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_pll_start_reconfig_ccd_pipe[1]~q ),
	.prn(vcc));
defparam \seq_pll_start_reconfig_ccd_pipe[1] .is_wysiwyg = "true";
defparam \seq_pll_start_reconfig_ccd_pipe[1] .power_up = "low";

dffeas \seq_pll_start_reconfig_ccd_pipe[2] (
	.clk(clk_0),
	.d(\seq_pll_start_reconfig_ccd_pipe[1]~q ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_pll_start_reconfig_ccd_pipe[2]~q ),
	.prn(vcc));
defparam \seq_pll_start_reconfig_ccd_pipe[2] .is_wysiwyg = "true";
defparam \seq_pll_start_reconfig_ccd_pipe[2] .power_up = "low";

dffeas pll_reconfig_reset_ams_n(
	.clk(\scan_clk~q ),
	.d(vcc),
	.asdata(vcc),
	.clrn(!\pll_reconfig_reset_n~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pll_reconfig_reset_ams_n~q ),
	.prn(vcc));
defparam pll_reconfig_reset_ams_n.is_wysiwyg = "true";
defparam pll_reconfig_reset_ams_n.power_up = "low";

dffeas pll_reconfig_reset_ams_n_r(
	.clk(\scan_clk~q ),
	.d(\pll_reconfig_reset_ams_n~q ),
	.asdata(vcc),
	.clrn(!\pll_reconfig_reset_n~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pll_reconfig_reset_ams_n_r~q ),
	.prn(vcc));
defparam pll_reconfig_reset_ams_n_r.is_wysiwyg = "true";
defparam pll_reconfig_reset_ams_n_r.power_up = "low";

dffeas seq_pll_start_reconfig_ams(
	.clk(\scan_clk~q ),
	.d(\seq_pll_start_reconfig_ccd_pipe[2]~q ),
	.asdata(vcc),
	.clrn(\pll_reconfig_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_pll_start_reconfig_ams~q ),
	.prn(vcc));
defparam seq_pll_start_reconfig_ams.is_wysiwyg = "true";
defparam seq_pll_start_reconfig_ams.power_up = "low";

dffeas seq_pll_start_reconfig_r(
	.clk(\scan_clk~q ),
	.d(\seq_pll_start_reconfig_ams~q ),
	.asdata(vcc),
	.clrn(\pll_reconfig_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_pll_start_reconfig_r~q ),
	.prn(vcc));
defparam seq_pll_start_reconfig_r.is_wysiwyg = "true";
defparam seq_pll_start_reconfig_r.power_up = "low";

dffeas seq_pll_start_reconfig_2r(
	.clk(\scan_clk~q ),
	.d(\seq_pll_start_reconfig_r~q ),
	.asdata(vcc),
	.clrn(\pll_reconfig_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_pll_start_reconfig_2r~q ),
	.prn(vcc));
defparam seq_pll_start_reconfig_2r.is_wysiwyg = "true";
defparam seq_pll_start_reconfig_2r.power_up = "low";

dffeas seq_pll_start_reconfig_3r(
	.clk(\scan_clk~q ),
	.d(\seq_pll_start_reconfig_2r~q ),
	.asdata(vcc),
	.clrn(\pll_reconfig_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_pll_start_reconfig_3r~q ),
	.prn(vcc));
defparam seq_pll_start_reconfig_3r.is_wysiwyg = "true";
defparam seq_pll_start_reconfig_3r.power_up = "low";

arriaii_lcell_comb pll_phase_auto_calibrate_pulse(
	.dataa(!\seq_pll_start_reconfig_2r~q ),
	.datab(!\seq_pll_start_reconfig_3r~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pll_phase_auto_calibrate_pulse~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam pll_phase_auto_calibrate_pulse.extended_lut = "off";
defparam pll_phase_auto_calibrate_pulse.lut_mask = 64'h4444444444444444;
defparam pll_phase_auto_calibrate_pulse.shared_arith = "off";

dffeas pll_reprogram_request_pulse(
	.clk(\scan_clk~q ),
	.d(\pll_phase_auto_calibrate_pulse~combout ),
	.asdata(vcc),
	.clrn(\pll_reconfig_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pll_reprogram_request_pulse~q ),
	.prn(vcc));
defparam pll_reprogram_request_pulse.is_wysiwyg = "true";
defparam pll_reprogram_request_pulse.power_up = "low";

dffeas pll_reprogram_request_pulse_r(
	.clk(\scan_clk~q ),
	.d(\pll_reprogram_request_pulse~q ),
	.asdata(vcc),
	.clrn(\pll_reconfig_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pll_reprogram_request_pulse_r~q ),
	.prn(vcc));
defparam pll_reprogram_request_pulse_r.is_wysiwyg = "true";
defparam pll_reprogram_request_pulse_r.power_up = "low";

arriaii_lcell_comb pll_reprogram_request_long_pulse(
	.dataa(!\pll_reprogram_request_pulse_2r~q ),
	.datab(!\pll_reprogram_request_pulse~q ),
	.datac(!\pll_reprogram_request_pulse_r~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pll_reprogram_request_long_pulse~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam pll_reprogram_request_long_pulse.extended_lut = "off";
defparam pll_reprogram_request_long_pulse.lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam pll_reprogram_request_long_pulse.shared_arith = "off";

dffeas pll_reprogram_request(
	.clk(\scan_clk~q ),
	.d(\pll_reprogram_request_long_pulse~combout ),
	.asdata(vcc),
	.clrn(\pll_reconfig_reset_ams_n_r~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pll_reprogram_request~q ),
	.prn(vcc));
defparam pll_reprogram_request.is_wysiwyg = "true";
defparam pll_reprogram_request.power_up = "low";

arriaii_lcell_comb \phs_shft_busy_siii~0 (
	.dataa(!\half_rate.pll|altpll_component|auto_generated|phasedone ),
	.datab(!\pll_reprogram_request~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\phs_shft_busy_siii~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \phs_shft_busy_siii~0 .extended_lut = "off";
defparam \phs_shft_busy_siii~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \phs_shft_busy_siii~0 .shared_arith = "off";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_pll (
	phasedone,
	pll1,
	clk_0,
	clk_1,
	clk_3,
	clk_4,
	clk_5,
	pll_lock_sync,
	locked,
	pll_new_dir,
	pll_reprogram_request,
	scan_clk,
	pll_new_phase_2,
	pll_new_phase_1,
	pll_new_phase_0,
	global_reset_n,
	pll_ref_clk)/* synthesis synthesis_greybox=0 */;
output 	phasedone;
output 	pll1;
output 	clk_0;
output 	clk_1;
output 	clk_3;
output 	clk_4;
output 	clk_5;
output 	pll_lock_sync;
output 	locked;
input 	pll_new_dir;
input 	pll_reprogram_request;
input 	scan_clk;
input 	pll_new_phase_2;
input 	pll_new_phase_1;
input 	pll_new_phase_0;
input 	global_reset_n;
input 	pll_ref_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_altpll_1 altpll_component(
	.phasedone(phasedone),
	.pll1(pll1),
	.clk_0(clk_0),
	.clk_1(clk_1),
	.clk_3(clk_3),
	.clk_4(clk_4),
	.clk_5(clk_5),
	.pll_lock_sync(pll_lock_sync),
	.locked(locked),
	.phaseupdown(pll_new_dir),
	.phasestep(pll_reprogram_request),
	.scanclk(scan_clk),
	.pll_new_phase_2(pll_new_phase_2),
	.pll_new_phase_1(pll_new_phase_1),
	.pll_new_phase_0(pll_new_phase_0),
	.areset(global_reset_n),
	.inclk({gnd,pll_ref_clk}));

endmodule

module ddr3_int_altpll_1 (
	phasedone,
	pll1,
	clk_0,
	clk_1,
	clk_3,
	clk_4,
	clk_5,
	pll_lock_sync,
	locked,
	phaseupdown,
	phasestep,
	scanclk,
	pll_new_phase_2,
	pll_new_phase_1,
	pll_new_phase_0,
	areset,
	inclk)/* synthesis synthesis_greybox=0 */;
output 	phasedone;
output 	pll1;
output 	clk_0;
output 	clk_1;
output 	clk_3;
output 	clk_4;
output 	clk_5;
output 	pll_lock_sync;
output 	locked;
input 	phaseupdown;
input 	phasestep;
input 	scanclk;
input 	pll_new_phase_2;
input 	pll_new_phase_1;
input 	pll_new_phase_0;
input 	areset;
input 	[1:0] inclk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_altpll_f5p3 auto_generated(
	.phasedone(phasedone),
	.pll11(pll1),
	.clk({clk_unconnected_wire_6,clk_5,clk_4,clk_3,clk_unconnected_wire_2,clk_1,clk_0}),
	.pll_lock_sync1(pll_lock_sync),
	.locked1(locked),
	.phaseupdown(phaseupdown),
	.phasestep(phasestep),
	.scanclk(scanclk),
	.pll_new_phase_2(pll_new_phase_2),
	.pll_new_phase_1(pll_new_phase_1),
	.pll_new_phase_0(pll_new_phase_0),
	.areset(areset),
	.inclk({gnd,inclk[0]}));

endmodule

module ddr3_int_altpll_f5p3 (
	phasedone,
	pll11,
	clk,
	pll_lock_sync1,
	locked1,
	phaseupdown,
	phasestep,
	scanclk,
	pll_new_phase_2,
	pll_new_phase_1,
	pll_new_phase_0,
	areset,
	inclk)/* synthesis synthesis_greybox=0 */;
output 	phasedone;
output 	pll11;
output 	[6:0] clk;
output 	pll_lock_sync1;
output 	locked1;
input 	phaseupdown;
input 	phasestep;
input 	scanclk;
input 	pll_new_phase_2;
input 	pll_new_phase_1;
input 	pll_new_phase_0;
input 	areset;
input 	[1:0] inclk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \clk[2] ;
wire \clk[6] ;
wire \pll1~CLK7 ;
wire \pll1~CLK8 ;
wire \pll1~CLK9 ;
wire \altpll_dyn_phase_le2|combout ;
wire \altpll_dyn_phase_le4|combout ;
wire \altpll_dyn_phase_le5|combout ;
wire \altpll_dyn_phase_le6|combout ;
wire \remap_decoy_le3a[0]~combout ;
wire \remap_decoy_le3a[1]~combout ;
wire \remap_decoy_le3a[2]~combout ;
wire \remap_decoy_le3a[3]~combout ;
wire \pll1~FBOUT ;

wire [9:0] pll1_CLK_bus;

assign clk[0] = pll1_CLK_bus[0];
assign clk[1] = pll1_CLK_bus[1];
assign \clk[2]  = pll1_CLK_bus[2];
assign clk[3] = pll1_CLK_bus[3];
assign clk[4] = pll1_CLK_bus[4];
assign clk[5] = pll1_CLK_bus[5];
assign \clk[6]  = pll1_CLK_bus[6];
assign \pll1~CLK7  = pll1_CLK_bus[7];
assign \pll1~CLK8  = pll1_CLK_bus[8];
assign \pll1~CLK9  = pll1_CLK_bus[9];

ddr3_int_altpll_dyn_phase_le_jdo altpll_dyn_phase_le2(
	.combout(\altpll_dyn_phase_le2|combout ),
	.remap_decoy_le3a_0(\remap_decoy_le3a[0]~combout ),
	.remap_decoy_le3a_1(\remap_decoy_le3a[1]~combout ),
	.remap_decoy_le3a_2(\remap_decoy_le3a[2]~combout ),
	.remap_decoy_le3a_3(\remap_decoy_le3a[3]~combout ));

ddr3_int_altpll_dyn_phase_le_kdo altpll_dyn_phase_le4(
	.combout(\altpll_dyn_phase_le4|combout ),
	.remap_decoy_le3a_0(\remap_decoy_le3a[0]~combout ),
	.remap_decoy_le3a_1(\remap_decoy_le3a[1]~combout ),
	.remap_decoy_le3a_2(\remap_decoy_le3a[2]~combout ),
	.remap_decoy_le3a_3(\remap_decoy_le3a[3]~combout ));

ddr3_int_altpll_dyn_phase_le_ldo altpll_dyn_phase_le5(
	.combout(\altpll_dyn_phase_le5|combout ),
	.remap_decoy_le3a_0(\remap_decoy_le3a[0]~combout ),
	.remap_decoy_le3a_1(\remap_decoy_le3a[1]~combout ),
	.remap_decoy_le3a_2(\remap_decoy_le3a[2]~combout ),
	.remap_decoy_le3a_3(\remap_decoy_le3a[3]~combout ));

ddr3_int_altpll_dyn_phase_le_mdo altpll_dyn_phase_le6(
	.combout(\altpll_dyn_phase_le6|combout ),
	.remap_decoy_le3a_0(\remap_decoy_le3a[0]~combout ),
	.remap_decoy_le3a_1(\remap_decoy_le3a[1]~combout ),
	.remap_decoy_le3a_2(\remap_decoy_le3a[2]~combout ),
	.remap_decoy_le3a_3(\remap_decoy_le3a[3]~combout ));

arriaii_lcell_comb \remap_decoy_le3a[0] (
	.dataa(!pll_new_phase_2),
	.datab(!pll_new_phase_1),
	.datac(!pll_new_phase_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\remap_decoy_le3a[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \remap_decoy_le3a[0] .extended_lut = "off";
defparam \remap_decoy_le3a[0] .lut_mask = 64'h6B6B6B6B6B6B6B6B;
defparam \remap_decoy_le3a[0] .shared_arith = "off";

arriaii_lcell_comb \remap_decoy_le3a[1] (
	.dataa(!pll_new_phase_2),
	.datab(!pll_new_phase_1),
	.datac(!pll_new_phase_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\remap_decoy_le3a[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \remap_decoy_le3a[1] .extended_lut = "off";
defparam \remap_decoy_le3a[1] .lut_mask = 64'hEDEDEDEDEDEDEDED;
defparam \remap_decoy_le3a[1] .shared_arith = "off";

arriaii_lcell_comb \remap_decoy_le3a[2] (
	.dataa(!pll_new_phase_2),
	.datab(!pll_new_phase_1),
	.datac(!pll_new_phase_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\remap_decoy_le3a[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \remap_decoy_le3a[2] .extended_lut = "off";
defparam \remap_decoy_le3a[2] .lut_mask = 64'h6767676767676767;
defparam \remap_decoy_le3a[2] .shared_arith = "off";

arriaii_lcell_comb \remap_decoy_le3a[3] (
	.dataa(!pll_new_phase_2),
	.datab(!pll_new_phase_1),
	.datac(!pll_new_phase_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\remap_decoy_le3a[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \remap_decoy_le3a[3] .extended_lut = "off";
defparam \remap_decoy_le3a[3] .lut_mask = 64'h7070707070707070;
defparam \remap_decoy_le3a[3] .shared_arith = "off";

arriaii_pll pll1(
	.areset(!areset),
	.pfdena(vcc),
	.fbin(\pll1~FBOUT ),
	.phaseupdown(phaseupdown),
	.phasestep(phasestep),
	.scandata(gnd),
	.scanclk(scanclk),
	.scanclkena(vcc),
	.configupdate(gnd),
	.clkswitch(gnd),
	.inclk({gnd,inclk[0]}),
	.phasecounterselect({\altpll_dyn_phase_le6|combout ,\altpll_dyn_phase_le5|combout ,\altpll_dyn_phase_le4|combout ,\altpll_dyn_phase_le2|combout }),
	.phasedone(phasedone),
	.scandataout(),
	.scandone(),
	.activeclock(),
	.locked(pll11),
	.vcooverrange(),
	.vcounderrange(),
	.fbout(\pll1~FBOUT ),
	.clk(pll1_CLK_bus),
	.clkbad());
defparam pll1.auto_settings = "false";
defparam pll1.bandwidth_type = "medium";
defparam pll1.c0_high = 4;
defparam pll1.c0_initial = 2;
defparam pll1.c0_low = 4;
defparam pll1.c0_mode = "even";
defparam pll1.c0_ph = 5;
defparam pll1.c1_high = 2;
defparam pll1.c1_initial = 2;
defparam pll1.c1_low = 2;
defparam pll1.c1_mode = "even";
defparam pll1.c1_ph = 0;
defparam pll1.c1_use_casc_in = "off";
defparam pll1.c2_high = 2;
defparam pll1.c2_initial = 1;
defparam pll1.c2_low = 2;
defparam pll1.c2_mode = "even";
defparam pll1.c2_ph = 0;
defparam pll1.c2_use_casc_in = "off";
defparam pll1.c3_high = 2;
defparam pll1.c3_initial = 2;
defparam pll1.c3_low = 2;
defparam pll1.c3_mode = "even";
defparam pll1.c3_ph = 0;
defparam pll1.c3_use_casc_in = "off";
defparam pll1.c4_high = 2;
defparam pll1.c4_initial = 2;
defparam pll1.c4_low = 2;
defparam pll1.c4_mode = "even";
defparam pll1.c4_ph = 0;
defparam pll1.c4_use_casc_in = "off";
defparam pll1.c5_high = 0;
defparam pll1.c5_initial = 0;
defparam pll1.c5_low = 0;
defparam pll1.c5_mode = "bypass";
defparam pll1.c5_ph = 0;
defparam pll1.c5_use_casc_in = "off";
defparam pll1.c6_high = 0;
defparam pll1.c6_initial = 0;
defparam pll1.c6_low = 0;
defparam pll1.c6_mode = "bypass";
defparam pll1.c6_ph = 0;
defparam pll1.c6_use_casc_in = "off";
defparam pll1.c7_high = 0;
defparam pll1.c7_initial = 0;
defparam pll1.c7_low = 0;
defparam pll1.c7_mode = "bypass";
defparam pll1.c7_ph = 0;
defparam pll1.c7_use_casc_in = "off";
defparam pll1.c8_high = 0;
defparam pll1.c8_initial = 0;
defparam pll1.c8_low = 0;
defparam pll1.c8_mode = "bypass";
defparam pll1.c8_ph = 0;
defparam pll1.c8_use_casc_in = "off";
defparam pll1.c9_high = 0;
defparam pll1.c9_initial = 0;
defparam pll1.c9_low = 0;
defparam pll1.c9_mode = "bypass";
defparam pll1.c9_ph = 0;
defparam pll1.c9_use_casc_in = "off";
defparam pll1.charge_pump_current_bits = 1;
defparam pll1.clk0_counter = "c0";
defparam pll1.clk0_divide_by = 1;
defparam pll1.clk0_duty_cycle = 50;
defparam pll1.clk0_multiply_by = 6;
defparam pll1.clk0_phase_shift = "521";
defparam pll1.clk1_counter = "c1";
defparam pll1.clk1_divide_by = 1;
defparam pll1.clk1_duty_cycle = 50;
defparam pll1.clk1_multiply_by = 12;
defparam pll1.clk1_phase_shift = "0";
defparam pll1.clk2_counter = "unused";
defparam pll1.clk2_divide_by = 0;
defparam pll1.clk2_duty_cycle = 50;
defparam pll1.clk2_multiply_by = 0;
defparam pll1.clk2_phase_shift = "0";
defparam pll1.clk3_counter = "c2";
defparam pll1.clk3_divide_by = 1;
defparam pll1.clk3_duty_cycle = 50;
defparam pll1.clk3_multiply_by = 12;
defparam pll1.clk3_phase_shift = "-833";
defparam pll1.clk4_counter = "c3";
defparam pll1.clk4_divide_by = 1;
defparam pll1.clk4_duty_cycle = 50;
defparam pll1.clk4_multiply_by = 12;
defparam pll1.clk4_phase_shift = "0";
defparam pll1.clk5_counter = "c4";
defparam pll1.clk5_divide_by = 1;
defparam pll1.clk5_duty_cycle = 50;
defparam pll1.clk5_multiply_by = 12;
defparam pll1.clk5_phase_shift = "0";
defparam pll1.clk6_counter = "unused";
defparam pll1.clk6_divide_by = 0;
defparam pll1.clk6_duty_cycle = 50;
defparam pll1.clk6_multiply_by = 0;
defparam pll1.clk6_phase_shift = "0";
defparam pll1.clk7_counter = "unused";
defparam pll1.clk7_divide_by = 0;
defparam pll1.clk7_duty_cycle = 50;
defparam pll1.clk7_multiply_by = 0;
defparam pll1.clk7_phase_shift = "0";
defparam pll1.clk8_counter = "unused";
defparam pll1.clk8_divide_by = 0;
defparam pll1.clk8_duty_cycle = 50;
defparam pll1.clk8_multiply_by = 0;
defparam pll1.clk8_phase_shift = "0";
defparam pll1.clk9_counter = "unused";
defparam pll1.clk9_divide_by = 0;
defparam pll1.clk9_duty_cycle = 50;
defparam pll1.clk9_multiply_by = 0;
defparam pll1.clk9_phase_shift = "0";
defparam pll1.dpa_divide_by = 0;
defparam pll1.dpa_divider = 1;
defparam pll1.dpa_multiply_by = 0;
defparam pll1.inclk0_input_frequency = 40000;
defparam pll1.inclk1_input_frequency = 0;
defparam pll1.loop_filter_c_bits = 0;
defparam pll1.loop_filter_r_bits = 24;
defparam pll1.m = 48;
defparam pll1.m_initial = 2;
defparam pll1.m_ph = 0;
defparam pll1.n = 1;
defparam pll1.operation_mode = "no compensation";
defparam pll1.pfd_max = 200000;
defparam pll1.pfd_min = 3076;
defparam pll1.pll_type = "fast";
defparam pll1.self_reset_on_loss_lock = "off";
defparam pll1.simulation_type = "timing";
defparam pll1.switch_over_type = "auto";
defparam pll1.vco_center = 769;
defparam pll1.vco_divide_by = 0;
defparam pll1.vco_frequency_control = "auto";
defparam pll1.vco_max = 1666;
defparam pll1.vco_min = 769;
defparam pll1.vco_multiply_by = 0;
defparam pll1.vco_phase_shift_step = 104;
defparam pll1.vco_post_scale = 1;

dffeas pll_lock_sync(
	.clk(pll11),
	.d(vcc),
	.asdata(vcc),
	.clrn(areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(pll_lock_sync1),
	.prn(vcc));
defparam pll_lock_sync.is_wysiwyg = "true";
defparam pll_lock_sync.power_up = "low";

arriaii_lcell_comb locked(
	.dataa(!pll11),
	.datab(!pll_lock_sync1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(locked1),
	.sumout(),
	.cout(),
	.shareout());
defparam locked.extended_lut = "off";
defparam locked.lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam locked.shared_arith = "off";

endmodule

module ddr3_int_altpll_dyn_phase_le_jdo (
	combout,
	remap_decoy_le3a_0,
	remap_decoy_le3a_1,
	remap_decoy_le3a_2,
	remap_decoy_le3a_3)/* synthesis synthesis_greybox=0 */;
output 	combout;
input 	remap_decoy_le3a_0;
input 	remap_decoy_le3a_1;
input 	remap_decoy_le3a_2;
input 	remap_decoy_le3a_3;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



arriaii_lcell_comb le_comb7(
	.dataa(!remap_decoy_le3a_0),
	.datab(!remap_decoy_le3a_1),
	.datac(!remap_decoy_le3a_2),
	.datad(!remap_decoy_le3a_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(combout),
	.sumout(),
	.cout(),
	.shareout());
defparam le_comb7.extended_lut = "off";
defparam le_comb7.lut_mask = 64'h5555555555555555;
defparam le_comb7.shared_arith = "off";

endmodule

module ddr3_int_altpll_dyn_phase_le_kdo (
	combout,
	remap_decoy_le3a_0,
	remap_decoy_le3a_1,
	remap_decoy_le3a_2,
	remap_decoy_le3a_3)/* synthesis synthesis_greybox=0 */;
output 	combout;
input 	remap_decoy_le3a_0;
input 	remap_decoy_le3a_1;
input 	remap_decoy_le3a_2;
input 	remap_decoy_le3a_3;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



arriaii_lcell_comb le_comb8(
	.dataa(!remap_decoy_le3a_0),
	.datab(!remap_decoy_le3a_1),
	.datac(!remap_decoy_le3a_2),
	.datad(!remap_decoy_le3a_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(combout),
	.sumout(),
	.cout(),
	.shareout());
defparam le_comb8.extended_lut = "off";
defparam le_comb8.lut_mask = 64'h3333333333333333;
defparam le_comb8.shared_arith = "off";

endmodule

module ddr3_int_altpll_dyn_phase_le_ldo (
	combout,
	remap_decoy_le3a_0,
	remap_decoy_le3a_1,
	remap_decoy_le3a_2,
	remap_decoy_le3a_3)/* synthesis synthesis_greybox=0 */;
output 	combout;
input 	remap_decoy_le3a_0;
input 	remap_decoy_le3a_1;
input 	remap_decoy_le3a_2;
input 	remap_decoy_le3a_3;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



arriaii_lcell_comb le_comb9(
	.dataa(!remap_decoy_le3a_0),
	.datab(!remap_decoy_le3a_1),
	.datac(!remap_decoy_le3a_2),
	.datad(!remap_decoy_le3a_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(combout),
	.sumout(),
	.cout(),
	.shareout());
defparam le_comb9.extended_lut = "off";
defparam le_comb9.lut_mask = 64'h0F0F0F0F0F0F0F0F;
defparam le_comb9.shared_arith = "off";

endmodule

module ddr3_int_altpll_dyn_phase_le_mdo (
	combout,
	remap_decoy_le3a_0,
	remap_decoy_le3a_1,
	remap_decoy_le3a_2,
	remap_decoy_le3a_3)/* synthesis synthesis_greybox=0 */;
output 	combout;
input 	remap_decoy_le3a_0;
input 	remap_decoy_le3a_1;
input 	remap_decoy_le3a_2;
input 	remap_decoy_le3a_3;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



arriaii_lcell_comb le_comb10(
	.dataa(!remap_decoy_le3a_0),
	.datab(!remap_decoy_le3a_1),
	.datac(!remap_decoy_le3a_2),
	.datad(!remap_decoy_le3a_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(combout),
	.sumout(),
	.cout(),
	.shareout());
defparam le_comb10.extended_lut = "off";
defparam le_comb10.lut_mask = 64'h00FF00FF00FF00FF;
defparam le_comb10.shared_arith = "off";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_reset_pipe (
	clock,
	ams_pipe_1,
	pre_clear)/* synthesis synthesis_greybox=0 */;
input 	clock;
output 	ams_pipe_1;
input 	pre_clear;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ams_pipe[0]~q ;


dffeas \ams_pipe[1] (
	.clk(clock),
	.d(\ams_pipe[0]~q ),
	.asdata(vcc),
	.clrn(pre_clear),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ams_pipe_1),
	.prn(vcc));
defparam \ams_pipe[1] .is_wysiwyg = "true";
defparam \ams_pipe[1] .power_up = "low";

dffeas \ams_pipe[0] (
	.clk(clock),
	.d(vcc),
	.asdata(vcc),
	.clrn(pre_clear),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ams_pipe[0]~q ),
	.prn(vcc));
defparam \ams_pipe[0] .is_wysiwyg = "true";
defparam \ams_pipe[0] .power_up = "low";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_reset_pipe_2 (
	clock,
	pre_clear,
	ams_pipe_1)/* synthesis synthesis_greybox=0 */;
input 	clock;
input 	pre_clear;
output 	ams_pipe_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ams_pipe[0]~q ;


dffeas \ams_pipe[1] (
	.clk(clock),
	.d(\ams_pipe[0]~q ),
	.asdata(vcc),
	.clrn(pre_clear),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ams_pipe_1),
	.prn(vcc));
defparam \ams_pipe[1] .is_wysiwyg = "true";
defparam \ams_pipe[1] .power_up = "low";

dffeas \ams_pipe[0] (
	.clk(clock),
	.d(vcc),
	.asdata(vcc),
	.clrn(pre_clear),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ams_pipe[0]~q ),
	.prn(vcc));
defparam \ams_pipe[0] .is_wysiwyg = "true";
defparam \ams_pipe[0] .power_up = "low";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_reset_pipe_3 (
	clock,
	pre_clear,
	ams_pipe_3)/* synthesis synthesis_greybox=0 */;
input 	clock;
input 	pre_clear;
output 	ams_pipe_3;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ams_pipe[0]~q ;
wire \ams_pipe[1]~q ;
wire \ams_pipe[2]~q ;


dffeas \ams_pipe[3] (
	.clk(clock),
	.d(\ams_pipe[2]~q ),
	.asdata(vcc),
	.clrn(pre_clear),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ams_pipe_3),
	.prn(vcc));
defparam \ams_pipe[3] .is_wysiwyg = "true";
defparam \ams_pipe[3] .power_up = "low";

dffeas \ams_pipe[0] (
	.clk(clock),
	.d(vcc),
	.asdata(vcc),
	.clrn(pre_clear),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ams_pipe[0]~q ),
	.prn(vcc));
defparam \ams_pipe[0] .is_wysiwyg = "true";
defparam \ams_pipe[0] .power_up = "low";

dffeas \ams_pipe[1] (
	.clk(clock),
	.d(\ams_pipe[0]~q ),
	.asdata(vcc),
	.clrn(pre_clear),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ams_pipe[1]~q ),
	.prn(vcc));
defparam \ams_pipe[1] .is_wysiwyg = "true";
defparam \ams_pipe[1] .power_up = "low";

dffeas \ams_pipe[2] (
	.clk(clock),
	.d(\ams_pipe[1]~q ),
	.asdata(vcc),
	.clrn(pre_clear),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ams_pipe[2]~q ),
	.prn(vcc));
defparam \ams_pipe[2] .is_wysiwyg = "true";
defparam \ams_pipe[2] .power_up = "low";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_reset_pipe_5 (
	clock,
	pre_clear,
	ams_pipe_0)/* synthesis synthesis_greybox=0 */;
input 	clock;
input 	pre_clear;
output 	ams_pipe_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \ams_pipe[0] (
	.clk(clock),
	.d(vcc),
	.asdata(vcc),
	.clrn(!pre_clear),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ams_pipe_0),
	.prn(vcc));
defparam \ams_pipe[0] .is_wysiwyg = "true";
defparam \ams_pipe[0] .power_up = "low";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_reset_pipe_6 (
	clock,
	ams_pipe_1,
	pre_clear)/* synthesis synthesis_greybox=0 */;
input 	clock;
output 	ams_pipe_1;
input 	pre_clear;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ams_pipe[0]~q ;


dffeas \ams_pipe[1] (
	.clk(clock),
	.d(\ams_pipe[0]~q ),
	.asdata(vcc),
	.clrn(!pre_clear),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ams_pipe_1),
	.prn(vcc));
defparam \ams_pipe[1] .is_wysiwyg = "true";
defparam \ams_pipe[1] .power_up = "low";

dffeas \ams_pipe[0] (
	.clk(clock),
	.d(vcc),
	.asdata(vcc),
	.clrn(!pre_clear),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ams_pipe[0]~q ),
	.prn(vcc));
defparam \ams_pipe[0] .is_wysiwyg = "true";
defparam \ams_pipe[0] .power_up = "low";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_reset_pipe_7 (
	clock,
	ams_pipe_1,
	pre_clear,
	ams_pipe_0)/* synthesis synthesis_greybox=0 */;
input 	clock;
output 	ams_pipe_1;
input 	pre_clear;
input 	ams_pipe_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \ams_pipe[1] (
	.clk(clock),
	.d(ams_pipe_0),
	.asdata(vcc),
	.clrn(!pre_clear),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ams_pipe_1),
	.prn(vcc));
defparam \ams_pipe[1] .is_wysiwyg = "true";
defparam \ams_pipe[1] .power_up = "low";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_reset_pipe_8 (
	clock,
	ams_pipe_1,
	pre_clear,
	ams_pipe_3)/* synthesis synthesis_greybox=0 */;
input 	clock;
input 	ams_pipe_1;
input 	pre_clear;
output 	ams_pipe_3;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ams_pipe[2]~q ;


dffeas \ams_pipe[3] (
	.clk(clock),
	.d(\ams_pipe[2]~q ),
	.asdata(vcc),
	.clrn(pre_clear),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ams_pipe_3),
	.prn(vcc));
defparam \ams_pipe[3] .is_wysiwyg = "true";
defparam \ams_pipe[3] .power_up = "low";

dffeas \ams_pipe[2] (
	.clk(clock),
	.d(ams_pipe_1),
	.asdata(vcc),
	.clrn(pre_clear),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ams_pipe[2]~q ),
	.prn(vcc));
defparam \ams_pipe[2] .is_wysiwyg = "true";
defparam \ams_pipe[2] .power_up = "low";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_dp_io (
	clk_1,
	clk_3,
	resync_clk_2x,
	dqs_delay_ctrl_0,
	dqs_delay_ctrl_1,
	dqs_delay_ctrl_2,
	dqs_delay_ctrl_3,
	dqs_delay_ctrl_4,
	dqs_delay_ctrl_5,
	wire_output_dq_0_output_ddio_out_inst_dataout,
	wire_output_dq_0_output_ddio_out_inst_dataout1,
	wire_output_dq_0_output_ddio_out_inst_dataout2,
	wire_output_dq_0_output_ddio_out_inst_dataout3,
	wdp_dm_l_2x_0,
	wdp_dm_h_2x_0,
	wdp_dm_l_2x_1,
	wdp_dm_h_2x_1,
	wdp_dm_l_2x_2,
	wdp_dm_h_2x_2,
	wdp_dm_l_2x_3,
	wdp_dm_h_2x_3,
	wire_bidir_dq_0_output_ddio_out_inst_dataout,
	wire_bidir_dq_1_output_ddio_out_inst_dataout,
	wire_bidir_dq_2_output_ddio_out_inst_dataout,
	wire_bidir_dq_3_output_ddio_out_inst_dataout,
	wire_bidir_dq_4_output_ddio_out_inst_dataout,
	wire_bidir_dq_5_output_ddio_out_inst_dataout,
	wire_bidir_dq_6_output_ddio_out_inst_dataout,
	wire_bidir_dq_7_output_ddio_out_inst_dataout,
	wire_bidir_dq_0_output_ddio_out_inst_dataout1,
	wire_bidir_dq_1_output_ddio_out_inst_dataout1,
	wire_bidir_dq_2_output_ddio_out_inst_dataout1,
	wire_bidir_dq_3_output_ddio_out_inst_dataout1,
	wire_bidir_dq_4_output_ddio_out_inst_dataout1,
	wire_bidir_dq_5_output_ddio_out_inst_dataout1,
	wire_bidir_dq_6_output_ddio_out_inst_dataout1,
	wire_bidir_dq_7_output_ddio_out_inst_dataout1,
	wire_bidir_dq_0_output_ddio_out_inst_dataout2,
	wire_bidir_dq_1_output_ddio_out_inst_dataout2,
	wire_bidir_dq_2_output_ddio_out_inst_dataout2,
	wire_bidir_dq_3_output_ddio_out_inst_dataout2,
	wire_bidir_dq_4_output_ddio_out_inst_dataout2,
	wire_bidir_dq_5_output_ddio_out_inst_dataout2,
	wire_bidir_dq_6_output_ddio_out_inst_dataout2,
	wire_bidir_dq_7_output_ddio_out_inst_dataout2,
	wire_bidir_dq_0_output_ddio_out_inst_dataout3,
	wire_bidir_dq_1_output_ddio_out_inst_dataout3,
	wire_bidir_dq_2_output_ddio_out_inst_dataout3,
	wire_bidir_dq_3_output_ddio_out_inst_dataout3,
	wire_bidir_dq_4_output_ddio_out_inst_dataout3,
	wire_bidir_dq_5_output_ddio_out_inst_dataout3,
	wire_bidir_dq_6_output_ddio_out_inst_dataout3,
	wire_bidir_dq_7_output_ddio_out_inst_dataout3,
	dqs_pseudo_diff_out_0,
	dqsn_pseudo_diff_out_0,
	dqs_pseudo_diff_out_1,
	dqsn_pseudo_diff_out_1,
	dqs_pseudo_diff_out_2,
	dqsn_pseudo_diff_out_2,
	dqs_pseudo_diff_out_3,
	dqsn_pseudo_diff_out_3,
	wdp_wdata_l_2x_0,
	wdp_wdata_h_2x_0,
	dq_oe_2x_0,
	wdp_wdata_l_2x_1,
	wdp_wdata_h_2x_1,
	wdp_wdata_l_2x_2,
	wdp_wdata_h_2x_2,
	wdp_wdata_l_2x_3,
	wdp_wdata_h_2x_3,
	wdp_wdata_l_2x_4,
	wdp_wdata_h_2x_4,
	dq_oe_2x_1,
	wdp_wdata_l_2x_5,
	wdp_wdata_h_2x_5,
	wdp_wdata_l_2x_6,
	wdp_wdata_h_2x_6,
	wdp_wdata_l_2x_7,
	wdp_wdata_h_2x_7,
	wdp_wdata_l_2x_8,
	wdp_wdata_h_2x_8,
	dq_oe_2x_2,
	wdp_wdata_l_2x_9,
	wdp_wdata_h_2x_9,
	wdp_wdata_l_2x_10,
	wdp_wdata_h_2x_10,
	wdp_wdata_l_2x_11,
	wdp_wdata_h_2x_11,
	wdp_wdata_l_2x_12,
	wdp_wdata_h_2x_12,
	dq_oe_2x_3,
	wdp_wdata_l_2x_13,
	wdp_wdata_h_2x_13,
	wdp_wdata_l_2x_14,
	wdp_wdata_h_2x_14,
	wdp_wdata_l_2x_15,
	wdp_wdata_h_2x_15,
	wdp_wdata_l_2x_16,
	wdp_wdata_h_2x_16,
	dq_oe_2x_4,
	wdp_wdata_l_2x_17,
	wdp_wdata_h_2x_17,
	wdp_wdata_l_2x_18,
	wdp_wdata_h_2x_18,
	wdp_wdata_l_2x_19,
	wdp_wdata_h_2x_19,
	wdp_wdata_l_2x_20,
	wdp_wdata_h_2x_20,
	dq_oe_2x_5,
	wdp_wdata_l_2x_21,
	wdp_wdata_h_2x_21,
	wdp_wdata_l_2x_22,
	wdp_wdata_h_2x_22,
	wdp_wdata_l_2x_23,
	wdp_wdata_h_2x_23,
	wdp_wdata_l_2x_24,
	wdp_wdata_h_2x_24,
	dq_oe_2x_6,
	wdp_wdata_l_2x_25,
	wdp_wdata_h_2x_25,
	wdp_wdata_l_2x_26,
	wdp_wdata_h_2x_26,
	wdp_wdata_l_2x_27,
	wdp_wdata_h_2x_27,
	wdp_wdata_l_2x_28,
	wdp_wdata_h_2x_28,
	dq_oe_2x_7,
	wdp_wdata_l_2x_29,
	wdp_wdata_h_2x_29,
	wdp_wdata_l_2x_30,
	wdp_wdata_h_2x_30,
	wdp_wdata_l_2x_31,
	wdp_wdata_h_2x_31,
	dq_datain_0,
	dq_datain_1,
	dq_datain_2,
	dq_datain_3,
	dq_datain_4,
	dq_datain_5,
	dq_datain_6,
	dq_datain_7,
	dq_datain_8,
	dq_datain_9,
	dq_datain_10,
	dq_datain_11,
	dq_datain_12,
	dq_datain_13,
	dq_datain_14,
	dq_datain_15,
	dq_datain_16,
	dq_datain_17,
	dq_datain_18,
	dq_datain_19,
	dq_datain_20,
	dq_datain_21,
	dq_datain_22,
	dq_datain_23,
	dq_datain_24,
	dq_datain_25,
	dq_datain_26,
	dq_datain_27,
	dq_datain_28,
	dq_datain_29,
	dq_datain_30,
	dq_datain_31,
	dqs_buffered_0,
	dqs_buffered_1,
	dqs_buffered_2,
	dqs_buffered_3,
	dio_rdata_h_2x_0,
	dio_rdata_h_2x_1,
	dio_rdata_h_2x_2,
	dio_rdata_h_2x_3,
	dio_rdata_h_2x_4,
	dio_rdata_h_2x_5,
	dio_rdata_h_2x_6,
	dio_rdata_h_2x_7,
	dio_rdata_h_2x_8,
	dio_rdata_h_2x_9,
	dio_rdata_h_2x_10,
	dio_rdata_h_2x_11,
	dio_rdata_h_2x_12,
	dio_rdata_h_2x_13,
	dio_rdata_h_2x_14,
	dio_rdata_h_2x_15,
	dio_rdata_h_2x_16,
	dio_rdata_h_2x_17,
	dio_rdata_h_2x_18,
	dio_rdata_h_2x_19,
	dio_rdata_h_2x_20,
	dio_rdata_h_2x_21,
	dio_rdata_h_2x_22,
	dio_rdata_h_2x_23,
	dio_rdata_h_2x_24,
	dio_rdata_h_2x_25,
	dio_rdata_h_2x_26,
	dio_rdata_h_2x_27,
	dio_rdata_h_2x_28,
	dio_rdata_h_2x_29,
	dio_rdata_h_2x_30,
	dio_rdata_h_2x_31,
	dio_rdata_l_2x_0,
	dio_rdata_l_2x_1,
	dio_rdata_l_2x_2,
	dio_rdata_l_2x_3,
	dio_rdata_l_2x_4,
	dio_rdata_l_2x_5,
	dio_rdata_l_2x_6,
	dio_rdata_l_2x_7,
	dio_rdata_l_2x_8,
	dio_rdata_l_2x_9,
	dio_rdata_l_2x_10,
	dio_rdata_l_2x_11,
	dio_rdata_l_2x_12,
	dio_rdata_l_2x_13,
	dio_rdata_l_2x_14,
	dio_rdata_l_2x_15,
	dio_rdata_l_2x_16,
	dio_rdata_l_2x_17,
	dio_rdata_l_2x_18,
	dio_rdata_l_2x_19,
	dio_rdata_l_2x_20,
	dio_rdata_l_2x_21,
	dio_rdata_l_2x_22,
	dio_rdata_l_2x_23,
	dio_rdata_l_2x_24,
	dio_rdata_l_2x_25,
	dio_rdata_l_2x_26,
	dio_rdata_l_2x_27,
	dio_rdata_l_2x_28,
	dio_rdata_l_2x_29,
	dio_rdata_l_2x_30,
	dio_rdata_l_2x_31,
	bidir_dq_0_oe_ff_inst,
	bidir_dq_1_oe_ff_inst,
	bidir_dq_2_oe_ff_inst,
	bidir_dq_3_oe_ff_inst,
	bidir_dq_4_oe_ff_inst,
	bidir_dq_5_oe_ff_inst,
	bidir_dq_6_oe_ff_inst,
	bidir_dq_7_oe_ff_inst,
	bidir_dq_0_oe_ff_inst1,
	bidir_dq_1_oe_ff_inst1,
	bidir_dq_2_oe_ff_inst1,
	bidir_dq_3_oe_ff_inst1,
	bidir_dq_4_oe_ff_inst1,
	bidir_dq_5_oe_ff_inst1,
	bidir_dq_6_oe_ff_inst1,
	bidir_dq_7_oe_ff_inst1,
	bidir_dq_0_oe_ff_inst2,
	bidir_dq_1_oe_ff_inst2,
	bidir_dq_2_oe_ff_inst2,
	bidir_dq_3_oe_ff_inst2,
	bidir_dq_4_oe_ff_inst2,
	bidir_dq_5_oe_ff_inst2,
	bidir_dq_6_oe_ff_inst2,
	bidir_dq_7_oe_ff_inst2,
	bidir_dq_0_oe_ff_inst3,
	bidir_dq_1_oe_ff_inst3,
	bidir_dq_2_oe_ff_inst3,
	bidir_dq_3_oe_ff_inst3,
	bidir_dq_4_oe_ff_inst3,
	bidir_dq_5_oe_ff_inst3,
	bidir_dq_6_oe_ff_inst3,
	bidir_dq_7_oe_ff_inst3,
	dqs_0_oe_ff_inst,
	dqs_0_oe_ff_inst1,
	dqs_0_oe_ff_inst2,
	dqs_0_oe_ff_inst3,
	dqsn_0_oe_ff_inst,
	dqsn_0_oe_ff_inst1,
	dqsn_0_oe_ff_inst2,
	dqsn_0_oe_ff_inst3,
	ams_pipe_3,
	dqs_burst_2x_r3_0,
	dqs_burst_2x_r3_1,
	dqs_burst_2x_r3_2,
	dqs_burst_2x_r3_3,
	postamble_en_pos_2x_0,
	postamble_en_pos_2x_1,
	postamble_en_pos_2x_2,
	postamble_en_pos_2x_3)/* synthesis synthesis_greybox=0 */;
input 	clk_1;
input 	clk_3;
input 	resync_clk_2x;
input 	dqs_delay_ctrl_0;
input 	dqs_delay_ctrl_1;
input 	dqs_delay_ctrl_2;
input 	dqs_delay_ctrl_3;
input 	dqs_delay_ctrl_4;
input 	dqs_delay_ctrl_5;
output 	wire_output_dq_0_output_ddio_out_inst_dataout;
output 	wire_output_dq_0_output_ddio_out_inst_dataout1;
output 	wire_output_dq_0_output_ddio_out_inst_dataout2;
output 	wire_output_dq_0_output_ddio_out_inst_dataout3;
input 	wdp_dm_l_2x_0;
input 	wdp_dm_h_2x_0;
input 	wdp_dm_l_2x_1;
input 	wdp_dm_h_2x_1;
input 	wdp_dm_l_2x_2;
input 	wdp_dm_h_2x_2;
input 	wdp_dm_l_2x_3;
input 	wdp_dm_h_2x_3;
output 	wire_bidir_dq_0_output_ddio_out_inst_dataout;
output 	wire_bidir_dq_1_output_ddio_out_inst_dataout;
output 	wire_bidir_dq_2_output_ddio_out_inst_dataout;
output 	wire_bidir_dq_3_output_ddio_out_inst_dataout;
output 	wire_bidir_dq_4_output_ddio_out_inst_dataout;
output 	wire_bidir_dq_5_output_ddio_out_inst_dataout;
output 	wire_bidir_dq_6_output_ddio_out_inst_dataout;
output 	wire_bidir_dq_7_output_ddio_out_inst_dataout;
output 	wire_bidir_dq_0_output_ddio_out_inst_dataout1;
output 	wire_bidir_dq_1_output_ddio_out_inst_dataout1;
output 	wire_bidir_dq_2_output_ddio_out_inst_dataout1;
output 	wire_bidir_dq_3_output_ddio_out_inst_dataout1;
output 	wire_bidir_dq_4_output_ddio_out_inst_dataout1;
output 	wire_bidir_dq_5_output_ddio_out_inst_dataout1;
output 	wire_bidir_dq_6_output_ddio_out_inst_dataout1;
output 	wire_bidir_dq_7_output_ddio_out_inst_dataout1;
output 	wire_bidir_dq_0_output_ddio_out_inst_dataout2;
output 	wire_bidir_dq_1_output_ddio_out_inst_dataout2;
output 	wire_bidir_dq_2_output_ddio_out_inst_dataout2;
output 	wire_bidir_dq_3_output_ddio_out_inst_dataout2;
output 	wire_bidir_dq_4_output_ddio_out_inst_dataout2;
output 	wire_bidir_dq_5_output_ddio_out_inst_dataout2;
output 	wire_bidir_dq_6_output_ddio_out_inst_dataout2;
output 	wire_bidir_dq_7_output_ddio_out_inst_dataout2;
output 	wire_bidir_dq_0_output_ddio_out_inst_dataout3;
output 	wire_bidir_dq_1_output_ddio_out_inst_dataout3;
output 	wire_bidir_dq_2_output_ddio_out_inst_dataout3;
output 	wire_bidir_dq_3_output_ddio_out_inst_dataout3;
output 	wire_bidir_dq_4_output_ddio_out_inst_dataout3;
output 	wire_bidir_dq_5_output_ddio_out_inst_dataout3;
output 	wire_bidir_dq_6_output_ddio_out_inst_dataout3;
output 	wire_bidir_dq_7_output_ddio_out_inst_dataout3;
output 	dqs_pseudo_diff_out_0;
output 	dqsn_pseudo_diff_out_0;
output 	dqs_pseudo_diff_out_1;
output 	dqsn_pseudo_diff_out_1;
output 	dqs_pseudo_diff_out_2;
output 	dqsn_pseudo_diff_out_2;
output 	dqs_pseudo_diff_out_3;
output 	dqsn_pseudo_diff_out_3;
input 	wdp_wdata_l_2x_0;
input 	wdp_wdata_h_2x_0;
input 	dq_oe_2x_0;
input 	wdp_wdata_l_2x_1;
input 	wdp_wdata_h_2x_1;
input 	wdp_wdata_l_2x_2;
input 	wdp_wdata_h_2x_2;
input 	wdp_wdata_l_2x_3;
input 	wdp_wdata_h_2x_3;
input 	wdp_wdata_l_2x_4;
input 	wdp_wdata_h_2x_4;
input 	dq_oe_2x_1;
input 	wdp_wdata_l_2x_5;
input 	wdp_wdata_h_2x_5;
input 	wdp_wdata_l_2x_6;
input 	wdp_wdata_h_2x_6;
input 	wdp_wdata_l_2x_7;
input 	wdp_wdata_h_2x_7;
input 	wdp_wdata_l_2x_8;
input 	wdp_wdata_h_2x_8;
input 	dq_oe_2x_2;
input 	wdp_wdata_l_2x_9;
input 	wdp_wdata_h_2x_9;
input 	wdp_wdata_l_2x_10;
input 	wdp_wdata_h_2x_10;
input 	wdp_wdata_l_2x_11;
input 	wdp_wdata_h_2x_11;
input 	wdp_wdata_l_2x_12;
input 	wdp_wdata_h_2x_12;
input 	dq_oe_2x_3;
input 	wdp_wdata_l_2x_13;
input 	wdp_wdata_h_2x_13;
input 	wdp_wdata_l_2x_14;
input 	wdp_wdata_h_2x_14;
input 	wdp_wdata_l_2x_15;
input 	wdp_wdata_h_2x_15;
input 	wdp_wdata_l_2x_16;
input 	wdp_wdata_h_2x_16;
input 	dq_oe_2x_4;
input 	wdp_wdata_l_2x_17;
input 	wdp_wdata_h_2x_17;
input 	wdp_wdata_l_2x_18;
input 	wdp_wdata_h_2x_18;
input 	wdp_wdata_l_2x_19;
input 	wdp_wdata_h_2x_19;
input 	wdp_wdata_l_2x_20;
input 	wdp_wdata_h_2x_20;
input 	dq_oe_2x_5;
input 	wdp_wdata_l_2x_21;
input 	wdp_wdata_h_2x_21;
input 	wdp_wdata_l_2x_22;
input 	wdp_wdata_h_2x_22;
input 	wdp_wdata_l_2x_23;
input 	wdp_wdata_h_2x_23;
input 	wdp_wdata_l_2x_24;
input 	wdp_wdata_h_2x_24;
input 	dq_oe_2x_6;
input 	wdp_wdata_l_2x_25;
input 	wdp_wdata_h_2x_25;
input 	wdp_wdata_l_2x_26;
input 	wdp_wdata_h_2x_26;
input 	wdp_wdata_l_2x_27;
input 	wdp_wdata_h_2x_27;
input 	wdp_wdata_l_2x_28;
input 	wdp_wdata_h_2x_28;
input 	dq_oe_2x_7;
input 	wdp_wdata_l_2x_29;
input 	wdp_wdata_h_2x_29;
input 	wdp_wdata_l_2x_30;
input 	wdp_wdata_h_2x_30;
input 	wdp_wdata_l_2x_31;
input 	wdp_wdata_h_2x_31;
input 	dq_datain_0;
input 	dq_datain_1;
input 	dq_datain_2;
input 	dq_datain_3;
input 	dq_datain_4;
input 	dq_datain_5;
input 	dq_datain_6;
input 	dq_datain_7;
input 	dq_datain_8;
input 	dq_datain_9;
input 	dq_datain_10;
input 	dq_datain_11;
input 	dq_datain_12;
input 	dq_datain_13;
input 	dq_datain_14;
input 	dq_datain_15;
input 	dq_datain_16;
input 	dq_datain_17;
input 	dq_datain_18;
input 	dq_datain_19;
input 	dq_datain_20;
input 	dq_datain_21;
input 	dq_datain_22;
input 	dq_datain_23;
input 	dq_datain_24;
input 	dq_datain_25;
input 	dq_datain_26;
input 	dq_datain_27;
input 	dq_datain_28;
input 	dq_datain_29;
input 	dq_datain_30;
input 	dq_datain_31;
input 	dqs_buffered_0;
input 	dqs_buffered_1;
input 	dqs_buffered_2;
input 	dqs_buffered_3;
output 	dio_rdata_h_2x_0;
output 	dio_rdata_h_2x_1;
output 	dio_rdata_h_2x_2;
output 	dio_rdata_h_2x_3;
output 	dio_rdata_h_2x_4;
output 	dio_rdata_h_2x_5;
output 	dio_rdata_h_2x_6;
output 	dio_rdata_h_2x_7;
output 	dio_rdata_h_2x_8;
output 	dio_rdata_h_2x_9;
output 	dio_rdata_h_2x_10;
output 	dio_rdata_h_2x_11;
output 	dio_rdata_h_2x_12;
output 	dio_rdata_h_2x_13;
output 	dio_rdata_h_2x_14;
output 	dio_rdata_h_2x_15;
output 	dio_rdata_h_2x_16;
output 	dio_rdata_h_2x_17;
output 	dio_rdata_h_2x_18;
output 	dio_rdata_h_2x_19;
output 	dio_rdata_h_2x_20;
output 	dio_rdata_h_2x_21;
output 	dio_rdata_h_2x_22;
output 	dio_rdata_h_2x_23;
output 	dio_rdata_h_2x_24;
output 	dio_rdata_h_2x_25;
output 	dio_rdata_h_2x_26;
output 	dio_rdata_h_2x_27;
output 	dio_rdata_h_2x_28;
output 	dio_rdata_h_2x_29;
output 	dio_rdata_h_2x_30;
output 	dio_rdata_h_2x_31;
output 	dio_rdata_l_2x_0;
output 	dio_rdata_l_2x_1;
output 	dio_rdata_l_2x_2;
output 	dio_rdata_l_2x_3;
output 	dio_rdata_l_2x_4;
output 	dio_rdata_l_2x_5;
output 	dio_rdata_l_2x_6;
output 	dio_rdata_l_2x_7;
output 	dio_rdata_l_2x_8;
output 	dio_rdata_l_2x_9;
output 	dio_rdata_l_2x_10;
output 	dio_rdata_l_2x_11;
output 	dio_rdata_l_2x_12;
output 	dio_rdata_l_2x_13;
output 	dio_rdata_l_2x_14;
output 	dio_rdata_l_2x_15;
output 	dio_rdata_l_2x_16;
output 	dio_rdata_l_2x_17;
output 	dio_rdata_l_2x_18;
output 	dio_rdata_l_2x_19;
output 	dio_rdata_l_2x_20;
output 	dio_rdata_l_2x_21;
output 	dio_rdata_l_2x_22;
output 	dio_rdata_l_2x_23;
output 	dio_rdata_l_2x_24;
output 	dio_rdata_l_2x_25;
output 	dio_rdata_l_2x_26;
output 	dio_rdata_l_2x_27;
output 	dio_rdata_l_2x_28;
output 	dio_rdata_l_2x_29;
output 	dio_rdata_l_2x_30;
output 	dio_rdata_l_2x_31;
output 	bidir_dq_0_oe_ff_inst;
output 	bidir_dq_1_oe_ff_inst;
output 	bidir_dq_2_oe_ff_inst;
output 	bidir_dq_3_oe_ff_inst;
output 	bidir_dq_4_oe_ff_inst;
output 	bidir_dq_5_oe_ff_inst;
output 	bidir_dq_6_oe_ff_inst;
output 	bidir_dq_7_oe_ff_inst;
output 	bidir_dq_0_oe_ff_inst1;
output 	bidir_dq_1_oe_ff_inst1;
output 	bidir_dq_2_oe_ff_inst1;
output 	bidir_dq_3_oe_ff_inst1;
output 	bidir_dq_4_oe_ff_inst1;
output 	bidir_dq_5_oe_ff_inst1;
output 	bidir_dq_6_oe_ff_inst1;
output 	bidir_dq_7_oe_ff_inst1;
output 	bidir_dq_0_oe_ff_inst2;
output 	bidir_dq_1_oe_ff_inst2;
output 	bidir_dq_2_oe_ff_inst2;
output 	bidir_dq_3_oe_ff_inst2;
output 	bidir_dq_4_oe_ff_inst2;
output 	bidir_dq_5_oe_ff_inst2;
output 	bidir_dq_6_oe_ff_inst2;
output 	bidir_dq_7_oe_ff_inst2;
output 	bidir_dq_0_oe_ff_inst3;
output 	bidir_dq_1_oe_ff_inst3;
output 	bidir_dq_2_oe_ff_inst3;
output 	bidir_dq_3_oe_ff_inst3;
output 	bidir_dq_4_oe_ff_inst3;
output 	bidir_dq_5_oe_ff_inst3;
output 	bidir_dq_6_oe_ff_inst3;
output 	bidir_dq_7_oe_ff_inst3;
output 	dqs_0_oe_ff_inst;
output 	dqs_0_oe_ff_inst1;
output 	dqs_0_oe_ff_inst2;
output 	dqs_0_oe_ff_inst3;
output 	dqsn_0_oe_ff_inst;
output 	dqsn_0_oe_ff_inst1;
output 	dqsn_0_oe_ff_inst2;
output 	dqsn_0_oe_ff_inst3;
input 	ams_pipe_3;
input 	dqs_burst_2x_r3_0;
input 	dqs_burst_2x_r3_1;
input 	dqs_burst_2x_r3_2;
input 	dqs_burst_2x_r3_3;
input 	postamble_en_pos_2x_0;
input 	postamble_en_pos_2x_1;
input 	postamble_en_pos_2x_2;
input 	postamble_en_pos_2x_3;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \dqs_group[0].dq_dqs|wire_bidir_dq_0_ddio_in_inst_regoutlo ;
wire \dqs_group[0].dq_dqs|wire_bidir_dq_0_ddio_in_inst_regouthi ;
wire \dqs_group[0].dq_dqs|wire_bidir_dq_1_ddio_in_inst_regoutlo ;
wire \dqs_group[0].dq_dqs|wire_bidir_dq_1_ddio_in_inst_regouthi ;
wire \dqs_group[0].dq_dqs|wire_bidir_dq_2_ddio_in_inst_regoutlo ;
wire \dqs_group[0].dq_dqs|wire_bidir_dq_2_ddio_in_inst_regouthi ;
wire \dqs_group[0].dq_dqs|wire_bidir_dq_3_ddio_in_inst_regoutlo ;
wire \dqs_group[0].dq_dqs|wire_bidir_dq_3_ddio_in_inst_regouthi ;
wire \dqs_group[0].dq_dqs|wire_bidir_dq_4_ddio_in_inst_regoutlo ;
wire \dqs_group[0].dq_dqs|wire_bidir_dq_4_ddio_in_inst_regouthi ;
wire \dqs_group[0].dq_dqs|wire_bidir_dq_5_ddio_in_inst_regoutlo ;
wire \dqs_group[0].dq_dqs|wire_bidir_dq_5_ddio_in_inst_regouthi ;
wire \dqs_group[0].dq_dqs|wire_bidir_dq_6_ddio_in_inst_regoutlo ;
wire \dqs_group[0].dq_dqs|wire_bidir_dq_6_ddio_in_inst_regouthi ;
wire \dqs_group[0].dq_dqs|wire_bidir_dq_7_ddio_in_inst_regoutlo ;
wire \dqs_group[0].dq_dqs|wire_bidir_dq_7_ddio_in_inst_regouthi ;
wire \dqs_group[1].dq_dqs|wire_bidir_dq_0_ddio_in_inst_regoutlo ;
wire \dqs_group[1].dq_dqs|wire_bidir_dq_0_ddio_in_inst_regouthi ;
wire \dqs_group[1].dq_dqs|wire_bidir_dq_1_ddio_in_inst_regoutlo ;
wire \dqs_group[1].dq_dqs|wire_bidir_dq_1_ddio_in_inst_regouthi ;
wire \dqs_group[1].dq_dqs|wire_bidir_dq_2_ddio_in_inst_regoutlo ;
wire \dqs_group[1].dq_dqs|wire_bidir_dq_2_ddio_in_inst_regouthi ;
wire \dqs_group[1].dq_dqs|wire_bidir_dq_3_ddio_in_inst_regoutlo ;
wire \dqs_group[1].dq_dqs|wire_bidir_dq_3_ddio_in_inst_regouthi ;
wire \dqs_group[1].dq_dqs|wire_bidir_dq_4_ddio_in_inst_regoutlo ;
wire \dqs_group[1].dq_dqs|wire_bidir_dq_4_ddio_in_inst_regouthi ;
wire \dqs_group[1].dq_dqs|wire_bidir_dq_5_ddio_in_inst_regoutlo ;
wire \dqs_group[1].dq_dqs|wire_bidir_dq_5_ddio_in_inst_regouthi ;
wire \dqs_group[1].dq_dqs|wire_bidir_dq_6_ddio_in_inst_regoutlo ;
wire \dqs_group[1].dq_dqs|wire_bidir_dq_6_ddio_in_inst_regouthi ;
wire \dqs_group[1].dq_dqs|wire_bidir_dq_7_ddio_in_inst_regoutlo ;
wire \dqs_group[1].dq_dqs|wire_bidir_dq_7_ddio_in_inst_regouthi ;
wire \dqs_group[2].dq_dqs|wire_bidir_dq_0_ddio_in_inst_regoutlo ;
wire \dqs_group[2].dq_dqs|wire_bidir_dq_0_ddio_in_inst_regouthi ;
wire \dqs_group[2].dq_dqs|wire_bidir_dq_1_ddio_in_inst_regoutlo ;
wire \dqs_group[2].dq_dqs|wire_bidir_dq_1_ddio_in_inst_regouthi ;
wire \dqs_group[2].dq_dqs|wire_bidir_dq_2_ddio_in_inst_regoutlo ;
wire \dqs_group[2].dq_dqs|wire_bidir_dq_2_ddio_in_inst_regouthi ;
wire \dqs_group[2].dq_dqs|wire_bidir_dq_3_ddio_in_inst_regoutlo ;
wire \dqs_group[2].dq_dqs|wire_bidir_dq_3_ddio_in_inst_regouthi ;
wire \dqs_group[2].dq_dqs|wire_bidir_dq_4_ddio_in_inst_regoutlo ;
wire \dqs_group[2].dq_dqs|wire_bidir_dq_4_ddio_in_inst_regouthi ;
wire \dqs_group[2].dq_dqs|wire_bidir_dq_5_ddio_in_inst_regoutlo ;
wire \dqs_group[2].dq_dqs|wire_bidir_dq_5_ddio_in_inst_regouthi ;
wire \dqs_group[2].dq_dqs|wire_bidir_dq_6_ddio_in_inst_regoutlo ;
wire \dqs_group[2].dq_dqs|wire_bidir_dq_6_ddio_in_inst_regouthi ;
wire \dqs_group[2].dq_dqs|wire_bidir_dq_7_ddio_in_inst_regoutlo ;
wire \dqs_group[2].dq_dqs|wire_bidir_dq_7_ddio_in_inst_regouthi ;
wire \dqs_group[3].dq_dqs|wire_bidir_dq_0_ddio_in_inst_regoutlo ;
wire \dqs_group[3].dq_dqs|wire_bidir_dq_0_ddio_in_inst_regouthi ;
wire \dqs_group[3].dq_dqs|wire_bidir_dq_1_ddio_in_inst_regoutlo ;
wire \dqs_group[3].dq_dqs|wire_bidir_dq_1_ddio_in_inst_regouthi ;
wire \dqs_group[3].dq_dqs|wire_bidir_dq_2_ddio_in_inst_regoutlo ;
wire \dqs_group[3].dq_dqs|wire_bidir_dq_2_ddio_in_inst_regouthi ;
wire \dqs_group[3].dq_dqs|wire_bidir_dq_3_ddio_in_inst_regoutlo ;
wire \dqs_group[3].dq_dqs|wire_bidir_dq_3_ddio_in_inst_regouthi ;
wire \dqs_group[3].dq_dqs|wire_bidir_dq_4_ddio_in_inst_regoutlo ;
wire \dqs_group[3].dq_dqs|wire_bidir_dq_4_ddio_in_inst_regouthi ;
wire \dqs_group[3].dq_dqs|wire_bidir_dq_5_ddio_in_inst_regoutlo ;
wire \dqs_group[3].dq_dqs|wire_bidir_dq_5_ddio_in_inst_regouthi ;
wire \dqs_group[3].dq_dqs|wire_bidir_dq_6_ddio_in_inst_regoutlo ;
wire \dqs_group[3].dq_dqs|wire_bidir_dq_6_ddio_in_inst_regouthi ;
wire \dqs_group[3].dq_dqs|wire_bidir_dq_7_ddio_in_inst_regoutlo ;
wire \dqs_group[3].dq_dqs|wire_bidir_dq_7_ddio_in_inst_regouthi ;
wire \dqs_group[0].dq_dqs|wire_dqs_0_output_ddio_out_inst_dataout ;
wire \dqs_group[1].dq_dqs|wire_dqs_0_output_ddio_out_inst_dataout ;
wire \dqs_group[2].dq_dqs|wire_dqs_0_output_ddio_out_inst_dataout ;
wire \dqs_group[3].dq_dqs|wire_dqs_0_output_ddio_out_inst_dataout ;
wire \rdata_p_ams[0]~0_combout ;
wire \rdata_p_ams[0]~q ;
wire \dio_rdata_h_2x[0]~0_combout ;
wire \rdata_p_ams[1]~1_combout ;
wire \rdata_p_ams[1]~q ;
wire \dio_rdata_h_2x[1]~1_combout ;
wire \rdata_p_ams[2]~2_combout ;
wire \rdata_p_ams[2]~q ;
wire \dio_rdata_h_2x[2]~2_combout ;
wire \rdata_p_ams[3]~3_combout ;
wire \rdata_p_ams[3]~q ;
wire \dio_rdata_h_2x[3]~3_combout ;
wire \rdata_p_ams[4]~4_combout ;
wire \rdata_p_ams[4]~q ;
wire \dio_rdata_h_2x[4]~4_combout ;
wire \rdata_p_ams[5]~5_combout ;
wire \rdata_p_ams[5]~q ;
wire \dio_rdata_h_2x[5]~5_combout ;
wire \rdata_p_ams[6]~6_combout ;
wire \rdata_p_ams[6]~q ;
wire \dio_rdata_h_2x[6]~6_combout ;
wire \rdata_p_ams[7]~7_combout ;
wire \rdata_p_ams[7]~q ;
wire \dio_rdata_h_2x[7]~7_combout ;
wire \rdata_p_ams[8]~8_combout ;
wire \rdata_p_ams[8]~q ;
wire \dio_rdata_h_2x[8]~8_combout ;
wire \rdata_p_ams[9]~9_combout ;
wire \rdata_p_ams[9]~q ;
wire \dio_rdata_h_2x[9]~9_combout ;
wire \rdata_p_ams[10]~10_combout ;
wire \rdata_p_ams[10]~q ;
wire \dio_rdata_h_2x[10]~10_combout ;
wire \rdata_p_ams[11]~11_combout ;
wire \rdata_p_ams[11]~q ;
wire \dio_rdata_h_2x[11]~11_combout ;
wire \rdata_p_ams[12]~12_combout ;
wire \rdata_p_ams[12]~q ;
wire \dio_rdata_h_2x[12]~12_combout ;
wire \rdata_p_ams[13]~13_combout ;
wire \rdata_p_ams[13]~q ;
wire \dio_rdata_h_2x[13]~13_combout ;
wire \rdata_p_ams[14]~14_combout ;
wire \rdata_p_ams[14]~q ;
wire \dio_rdata_h_2x[14]~14_combout ;
wire \rdata_p_ams[15]~15_combout ;
wire \rdata_p_ams[15]~q ;
wire \dio_rdata_h_2x[15]~15_combout ;
wire \rdata_p_ams[16]~16_combout ;
wire \rdata_p_ams[16]~q ;
wire \dio_rdata_h_2x[16]~16_combout ;
wire \rdata_p_ams[17]~17_combout ;
wire \rdata_p_ams[17]~q ;
wire \dio_rdata_h_2x[17]~17_combout ;
wire \rdata_p_ams[18]~18_combout ;
wire \rdata_p_ams[18]~q ;
wire \dio_rdata_h_2x[18]~18_combout ;
wire \rdata_p_ams[19]~19_combout ;
wire \rdata_p_ams[19]~q ;
wire \dio_rdata_h_2x[19]~19_combout ;
wire \rdata_p_ams[20]~20_combout ;
wire \rdata_p_ams[20]~q ;
wire \dio_rdata_h_2x[20]~20_combout ;
wire \rdata_p_ams[21]~21_combout ;
wire \rdata_p_ams[21]~q ;
wire \dio_rdata_h_2x[21]~21_combout ;
wire \rdata_p_ams[22]~22_combout ;
wire \rdata_p_ams[22]~q ;
wire \dio_rdata_h_2x[22]~22_combout ;
wire \rdata_p_ams[23]~23_combout ;
wire \rdata_p_ams[23]~q ;
wire \dio_rdata_h_2x[23]~23_combout ;
wire \rdata_p_ams[24]~24_combout ;
wire \rdata_p_ams[24]~q ;
wire \dio_rdata_h_2x[24]~24_combout ;
wire \rdata_p_ams[25]~25_combout ;
wire \rdata_p_ams[25]~q ;
wire \dio_rdata_h_2x[25]~25_combout ;
wire \rdata_p_ams[26]~26_combout ;
wire \rdata_p_ams[26]~q ;
wire \dio_rdata_h_2x[26]~26_combout ;
wire \rdata_p_ams[27]~27_combout ;
wire \rdata_p_ams[27]~q ;
wire \dio_rdata_h_2x[27]~27_combout ;
wire \rdata_p_ams[28]~28_combout ;
wire \rdata_p_ams[28]~q ;
wire \dio_rdata_h_2x[28]~28_combout ;
wire \rdata_p_ams[29]~29_combout ;
wire \rdata_p_ams[29]~q ;
wire \dio_rdata_h_2x[29]~29_combout ;
wire \rdata_p_ams[30]~30_combout ;
wire \rdata_p_ams[30]~q ;
wire \dio_rdata_h_2x[30]~30_combout ;
wire \rdata_p_ams[31]~31_combout ;
wire \rdata_p_ams[31]~q ;
wire \dio_rdata_h_2x[31]~31_combout ;
wire \rdata_n_ams[0]~0_combout ;
wire \rdata_n_ams[0]~q ;
wire \dio_rdata_l_2x[0]~0_combout ;
wire \rdata_n_ams[1]~1_combout ;
wire \rdata_n_ams[1]~q ;
wire \dio_rdata_l_2x[1]~1_combout ;
wire \rdata_n_ams[2]~2_combout ;
wire \rdata_n_ams[2]~q ;
wire \dio_rdata_l_2x[2]~2_combout ;
wire \rdata_n_ams[3]~3_combout ;
wire \rdata_n_ams[3]~q ;
wire \dio_rdata_l_2x[3]~3_combout ;
wire \rdata_n_ams[4]~4_combout ;
wire \rdata_n_ams[4]~q ;
wire \dio_rdata_l_2x[4]~4_combout ;
wire \rdata_n_ams[5]~5_combout ;
wire \rdata_n_ams[5]~q ;
wire \dio_rdata_l_2x[5]~5_combout ;
wire \rdata_n_ams[6]~6_combout ;
wire \rdata_n_ams[6]~q ;
wire \dio_rdata_l_2x[6]~6_combout ;
wire \rdata_n_ams[7]~7_combout ;
wire \rdata_n_ams[7]~q ;
wire \dio_rdata_l_2x[7]~7_combout ;
wire \rdata_n_ams[8]~8_combout ;
wire \rdata_n_ams[8]~q ;
wire \dio_rdata_l_2x[8]~8_combout ;
wire \rdata_n_ams[9]~9_combout ;
wire \rdata_n_ams[9]~q ;
wire \dio_rdata_l_2x[9]~9_combout ;
wire \rdata_n_ams[10]~10_combout ;
wire \rdata_n_ams[10]~q ;
wire \dio_rdata_l_2x[10]~10_combout ;
wire \rdata_n_ams[11]~11_combout ;
wire \rdata_n_ams[11]~q ;
wire \dio_rdata_l_2x[11]~11_combout ;
wire \rdata_n_ams[12]~12_combout ;
wire \rdata_n_ams[12]~q ;
wire \dio_rdata_l_2x[12]~12_combout ;
wire \rdata_n_ams[13]~13_combout ;
wire \rdata_n_ams[13]~q ;
wire \dio_rdata_l_2x[13]~13_combout ;
wire \rdata_n_ams[14]~14_combout ;
wire \rdata_n_ams[14]~q ;
wire \dio_rdata_l_2x[14]~14_combout ;
wire \rdata_n_ams[15]~15_combout ;
wire \rdata_n_ams[15]~q ;
wire \dio_rdata_l_2x[15]~15_combout ;
wire \rdata_n_ams[16]~16_combout ;
wire \rdata_n_ams[16]~q ;
wire \dio_rdata_l_2x[16]~16_combout ;
wire \rdata_n_ams[17]~17_combout ;
wire \rdata_n_ams[17]~q ;
wire \dio_rdata_l_2x[17]~17_combout ;
wire \rdata_n_ams[18]~18_combout ;
wire \rdata_n_ams[18]~q ;
wire \dio_rdata_l_2x[18]~18_combout ;
wire \rdata_n_ams[19]~19_combout ;
wire \rdata_n_ams[19]~q ;
wire \dio_rdata_l_2x[19]~19_combout ;
wire \rdata_n_ams[20]~20_combout ;
wire \rdata_n_ams[20]~q ;
wire \dio_rdata_l_2x[20]~20_combout ;
wire \rdata_n_ams[21]~21_combout ;
wire \rdata_n_ams[21]~q ;
wire \dio_rdata_l_2x[21]~21_combout ;
wire \rdata_n_ams[22]~22_combout ;
wire \rdata_n_ams[22]~q ;
wire \dio_rdata_l_2x[22]~22_combout ;
wire \rdata_n_ams[23]~23_combout ;
wire \rdata_n_ams[23]~q ;
wire \dio_rdata_l_2x[23]~23_combout ;
wire \rdata_n_ams[24]~24_combout ;
wire \rdata_n_ams[24]~q ;
wire \dio_rdata_l_2x[24]~24_combout ;
wire \rdata_n_ams[25]~25_combout ;
wire \rdata_n_ams[25]~q ;
wire \dio_rdata_l_2x[25]~25_combout ;
wire \rdata_n_ams[26]~26_combout ;
wire \rdata_n_ams[26]~q ;
wire \dio_rdata_l_2x[26]~26_combout ;
wire \rdata_n_ams[27]~27_combout ;
wire \rdata_n_ams[27]~q ;
wire \dio_rdata_l_2x[27]~27_combout ;
wire \rdata_n_ams[28]~28_combout ;
wire \rdata_n_ams[28]~q ;
wire \dio_rdata_l_2x[28]~28_combout ;
wire \rdata_n_ams[29]~29_combout ;
wire \rdata_n_ams[29]~q ;
wire \dio_rdata_l_2x[29]~29_combout ;
wire \rdata_n_ams[30]~30_combout ;
wire \rdata_n_ams[30]~q ;
wire \dio_rdata_l_2x[30]~30_combout ;
wire \rdata_n_ams[31]~31_combout ;
wire \rdata_n_ams[31]~q ;
wire \dio_rdata_l_2x[31]~31_combout ;


ddr3_int_ddr3_int_phy_alt_mem_phy_dq_dqs \dqs_group[0].dq_dqs (
	.dqs_output_reg_clk(clk_1),
	.dq_output_reg_clk(clk_3),
	.dqs_enable_ctrl_clk(resync_clk_2x),
	.dll_delayctrlin({dqs_delay_ctrl_5,dqs_delay_ctrl_4,dqs_delay_ctrl_3,dqs_delay_ctrl_2,dqs_delay_ctrl_1,dqs_delay_ctrl_0}),
	.output_dq_output_data_out({wire_output_dq_0_output_ddio_out_inst_dataout}),
	.output_dq_output_data_in_low({wdp_dm_l_2x_0}),
	.output_dq_output_data_in_high({wdp_dm_h_2x_0}),
	.bidir_dq_output_data_out({wire_bidir_dq_7_output_ddio_out_inst_dataout,wire_bidir_dq_6_output_ddio_out_inst_dataout,wire_bidir_dq_5_output_ddio_out_inst_dataout,wire_bidir_dq_4_output_ddio_out_inst_dataout,wire_bidir_dq_3_output_ddio_out_inst_dataout,
wire_bidir_dq_2_output_ddio_out_inst_dataout,wire_bidir_dq_1_output_ddio_out_inst_dataout,wire_bidir_dq_0_output_ddio_out_inst_dataout}),
	.bidir_dq_input_data_out_low({\dqs_group[0].dq_dqs|wire_bidir_dq_7_ddio_in_inst_regoutlo ,\dqs_group[0].dq_dqs|wire_bidir_dq_6_ddio_in_inst_regoutlo ,\dqs_group[0].dq_dqs|wire_bidir_dq_5_ddio_in_inst_regoutlo ,\dqs_group[0].dq_dqs|wire_bidir_dq_4_ddio_in_inst_regoutlo ,
\dqs_group[0].dq_dqs|wire_bidir_dq_3_ddio_in_inst_regoutlo ,\dqs_group[0].dq_dqs|wire_bidir_dq_2_ddio_in_inst_regoutlo ,\dqs_group[0].dq_dqs|wire_bidir_dq_1_ddio_in_inst_regoutlo ,\dqs_group[0].dq_dqs|wire_bidir_dq_0_ddio_in_inst_regoutlo }),
	.bidir_dq_input_data_out_high({\dqs_group[0].dq_dqs|wire_bidir_dq_7_ddio_in_inst_regouthi ,\dqs_group[0].dq_dqs|wire_bidir_dq_6_ddio_in_inst_regouthi ,\dqs_group[0].dq_dqs|wire_bidir_dq_5_ddio_in_inst_regouthi ,\dqs_group[0].dq_dqs|wire_bidir_dq_4_ddio_in_inst_regouthi ,
\dqs_group[0].dq_dqs|wire_bidir_dq_3_ddio_in_inst_regouthi ,\dqs_group[0].dq_dqs|wire_bidir_dq_2_ddio_in_inst_regouthi ,\dqs_group[0].dq_dqs|wire_bidir_dq_1_ddio_in_inst_regouthi ,\dqs_group[0].dq_dqs|wire_bidir_dq_0_ddio_in_inst_regouthi }),
	.bidir_dq_output_data_in_low({wdp_wdata_l_2x_7,wdp_wdata_l_2x_6,wdp_wdata_l_2x_5,wdp_wdata_l_2x_4,wdp_wdata_l_2x_3,wdp_wdata_l_2x_2,wdp_wdata_l_2x_1,wdp_wdata_l_2x_0}),
	.bidir_dq_output_data_in_high({wdp_wdata_h_2x_7,wdp_wdata_h_2x_6,wdp_wdata_h_2x_5,wdp_wdata_h_2x_4,wdp_wdata_h_2x_3,wdp_wdata_h_2x_2,wdp_wdata_h_2x_1,wdp_wdata_h_2x_0}),
	.dq_oe_2x_0(dq_oe_2x_0),
	.dq_oe_2x_1(dq_oe_2x_1),
	.dqs_output_data_out({\dqs_group[0].dq_dqs|wire_dqs_0_output_ddio_out_inst_dataout }),
	.bidir_dq_input_data_in({dq_datain_7,dq_datain_6,dq_datain_5,dq_datain_4,dq_datain_3,dq_datain_2,dq_datain_1,dq_datain_0}),
	.dqs_input_data_in({dqs_buffered_0}),
	.bidir_dq_0_oe_ff_inst1(bidir_dq_0_oe_ff_inst),
	.bidir_dq_1_oe_ff_inst1(bidir_dq_1_oe_ff_inst),
	.bidir_dq_2_oe_ff_inst1(bidir_dq_2_oe_ff_inst),
	.bidir_dq_3_oe_ff_inst1(bidir_dq_3_oe_ff_inst),
	.bidir_dq_4_oe_ff_inst1(bidir_dq_4_oe_ff_inst),
	.bidir_dq_5_oe_ff_inst1(bidir_dq_5_oe_ff_inst),
	.bidir_dq_6_oe_ff_inst1(bidir_dq_6_oe_ff_inst),
	.bidir_dq_7_oe_ff_inst1(bidir_dq_7_oe_ff_inst),
	.dqs_0_oe_ff_inst1(dqs_0_oe_ff_inst),
	.dqsn_0_oe_ff_inst1(dqsn_0_oe_ff_inst),
	.bidir_dq_areset({ams_pipe_3,ams_pipe_3,ams_pipe_3,ams_pipe_3,ams_pipe_3,ams_pipe_3,ams_pipe_3,ams_pipe_3}),
	.dqs_output_data_in_high({dqs_burst_2x_r3_0}),
	.dqs_enable_ctrl_in(postamble_en_pos_2x_0));

ddr3_int_ddr3_int_phy_alt_mem_phy_dq_dqs_1 \dqs_group[1].dq_dqs (
	.dqs_output_reg_clk(clk_1),
	.dq_output_reg_clk(clk_3),
	.dqs_enable_ctrl_clk(resync_clk_2x),
	.dll_delayctrlin({dqs_delay_ctrl_5,dqs_delay_ctrl_4,dqs_delay_ctrl_3,dqs_delay_ctrl_2,dqs_delay_ctrl_1,dqs_delay_ctrl_0}),
	.output_dq_output_data_out({wire_output_dq_0_output_ddio_out_inst_dataout1}),
	.output_dq_output_data_in_low({wdp_dm_l_2x_1}),
	.output_dq_output_data_in_high({wdp_dm_h_2x_1}),
	.bidir_dq_output_data_out({wire_bidir_dq_7_output_ddio_out_inst_dataout1,wire_bidir_dq_6_output_ddio_out_inst_dataout1,wire_bidir_dq_5_output_ddio_out_inst_dataout1,wire_bidir_dq_4_output_ddio_out_inst_dataout1,wire_bidir_dq_3_output_ddio_out_inst_dataout1,
wire_bidir_dq_2_output_ddio_out_inst_dataout1,wire_bidir_dq_1_output_ddio_out_inst_dataout1,wire_bidir_dq_0_output_ddio_out_inst_dataout1}),
	.bidir_dq_input_data_out_low({\dqs_group[1].dq_dqs|wire_bidir_dq_7_ddio_in_inst_regoutlo ,\dqs_group[1].dq_dqs|wire_bidir_dq_6_ddio_in_inst_regoutlo ,\dqs_group[1].dq_dqs|wire_bidir_dq_5_ddio_in_inst_regoutlo ,\dqs_group[1].dq_dqs|wire_bidir_dq_4_ddio_in_inst_regoutlo ,
\dqs_group[1].dq_dqs|wire_bidir_dq_3_ddio_in_inst_regoutlo ,\dqs_group[1].dq_dqs|wire_bidir_dq_2_ddio_in_inst_regoutlo ,\dqs_group[1].dq_dqs|wire_bidir_dq_1_ddio_in_inst_regoutlo ,\dqs_group[1].dq_dqs|wire_bidir_dq_0_ddio_in_inst_regoutlo }),
	.bidir_dq_input_data_out_high({\dqs_group[1].dq_dqs|wire_bidir_dq_7_ddio_in_inst_regouthi ,\dqs_group[1].dq_dqs|wire_bidir_dq_6_ddio_in_inst_regouthi ,\dqs_group[1].dq_dqs|wire_bidir_dq_5_ddio_in_inst_regouthi ,\dqs_group[1].dq_dqs|wire_bidir_dq_4_ddio_in_inst_regouthi ,
\dqs_group[1].dq_dqs|wire_bidir_dq_3_ddio_in_inst_regouthi ,\dqs_group[1].dq_dqs|wire_bidir_dq_2_ddio_in_inst_regouthi ,\dqs_group[1].dq_dqs|wire_bidir_dq_1_ddio_in_inst_regouthi ,\dqs_group[1].dq_dqs|wire_bidir_dq_0_ddio_in_inst_regouthi }),
	.bidir_dq_output_data_in_low({wdp_wdata_l_2x_15,wdp_wdata_l_2x_14,wdp_wdata_l_2x_13,wdp_wdata_l_2x_12,wdp_wdata_l_2x_11,wdp_wdata_l_2x_10,wdp_wdata_l_2x_9,wdp_wdata_l_2x_8}),
	.bidir_dq_output_data_in_high({wdp_wdata_h_2x_15,wdp_wdata_h_2x_14,wdp_wdata_h_2x_13,wdp_wdata_h_2x_12,wdp_wdata_h_2x_11,wdp_wdata_h_2x_10,wdp_wdata_h_2x_9,wdp_wdata_h_2x_8}),
	.dq_oe_2x_2(dq_oe_2x_2),
	.dq_oe_2x_3(dq_oe_2x_3),
	.dqs_output_data_out({\dqs_group[1].dq_dqs|wire_dqs_0_output_ddio_out_inst_dataout }),
	.bidir_dq_input_data_in({dq_datain_15,dq_datain_14,dq_datain_13,dq_datain_12,dq_datain_11,dq_datain_10,dq_datain_9,dq_datain_8}),
	.dqs_input_data_in({dqs_buffered_1}),
	.bidir_dq_0_oe_ff_inst1(bidir_dq_0_oe_ff_inst1),
	.bidir_dq_1_oe_ff_inst1(bidir_dq_1_oe_ff_inst1),
	.bidir_dq_2_oe_ff_inst1(bidir_dq_2_oe_ff_inst1),
	.bidir_dq_3_oe_ff_inst1(bidir_dq_3_oe_ff_inst1),
	.bidir_dq_4_oe_ff_inst1(bidir_dq_4_oe_ff_inst1),
	.bidir_dq_5_oe_ff_inst1(bidir_dq_5_oe_ff_inst1),
	.bidir_dq_6_oe_ff_inst1(bidir_dq_6_oe_ff_inst1),
	.bidir_dq_7_oe_ff_inst1(bidir_dq_7_oe_ff_inst1),
	.dqs_0_oe_ff_inst1(dqs_0_oe_ff_inst1),
	.dqsn_0_oe_ff_inst1(dqsn_0_oe_ff_inst1),
	.bidir_dq_areset({ams_pipe_3,ams_pipe_3,ams_pipe_3,ams_pipe_3,ams_pipe_3,ams_pipe_3,ams_pipe_3,ams_pipe_3}),
	.dqs_output_data_in_high({dqs_burst_2x_r3_1}),
	.dqs_enable_ctrl_in(postamble_en_pos_2x_1));

ddr3_int_ddr3_int_phy_alt_mem_phy_dq_dqs_2 \dqs_group[2].dq_dqs (
	.dqs_output_reg_clk(clk_1),
	.dq_output_reg_clk(clk_3),
	.dqs_enable_ctrl_clk(resync_clk_2x),
	.dll_delayctrlin({dqs_delay_ctrl_5,dqs_delay_ctrl_4,dqs_delay_ctrl_3,dqs_delay_ctrl_2,dqs_delay_ctrl_1,dqs_delay_ctrl_0}),
	.output_dq_output_data_out({wire_output_dq_0_output_ddio_out_inst_dataout2}),
	.output_dq_output_data_in_low({wdp_dm_l_2x_2}),
	.output_dq_output_data_in_high({wdp_dm_h_2x_2}),
	.bidir_dq_output_data_out({wire_bidir_dq_7_output_ddio_out_inst_dataout2,wire_bidir_dq_6_output_ddio_out_inst_dataout2,wire_bidir_dq_5_output_ddio_out_inst_dataout2,wire_bidir_dq_4_output_ddio_out_inst_dataout2,wire_bidir_dq_3_output_ddio_out_inst_dataout2,
wire_bidir_dq_2_output_ddio_out_inst_dataout2,wire_bidir_dq_1_output_ddio_out_inst_dataout2,wire_bidir_dq_0_output_ddio_out_inst_dataout2}),
	.bidir_dq_input_data_out_low({\dqs_group[2].dq_dqs|wire_bidir_dq_7_ddio_in_inst_regoutlo ,\dqs_group[2].dq_dqs|wire_bidir_dq_6_ddio_in_inst_regoutlo ,\dqs_group[2].dq_dqs|wire_bidir_dq_5_ddio_in_inst_regoutlo ,\dqs_group[2].dq_dqs|wire_bidir_dq_4_ddio_in_inst_regoutlo ,
\dqs_group[2].dq_dqs|wire_bidir_dq_3_ddio_in_inst_regoutlo ,\dqs_group[2].dq_dqs|wire_bidir_dq_2_ddio_in_inst_regoutlo ,\dqs_group[2].dq_dqs|wire_bidir_dq_1_ddio_in_inst_regoutlo ,\dqs_group[2].dq_dqs|wire_bidir_dq_0_ddio_in_inst_regoutlo }),
	.bidir_dq_input_data_out_high({\dqs_group[2].dq_dqs|wire_bidir_dq_7_ddio_in_inst_regouthi ,\dqs_group[2].dq_dqs|wire_bidir_dq_6_ddio_in_inst_regouthi ,\dqs_group[2].dq_dqs|wire_bidir_dq_5_ddio_in_inst_regouthi ,\dqs_group[2].dq_dqs|wire_bidir_dq_4_ddio_in_inst_regouthi ,
\dqs_group[2].dq_dqs|wire_bidir_dq_3_ddio_in_inst_regouthi ,\dqs_group[2].dq_dqs|wire_bidir_dq_2_ddio_in_inst_regouthi ,\dqs_group[2].dq_dqs|wire_bidir_dq_1_ddio_in_inst_regouthi ,\dqs_group[2].dq_dqs|wire_bidir_dq_0_ddio_in_inst_regouthi }),
	.bidir_dq_output_data_in_low({wdp_wdata_l_2x_23,wdp_wdata_l_2x_22,wdp_wdata_l_2x_21,wdp_wdata_l_2x_20,wdp_wdata_l_2x_19,wdp_wdata_l_2x_18,wdp_wdata_l_2x_17,wdp_wdata_l_2x_16}),
	.bidir_dq_output_data_in_high({wdp_wdata_h_2x_23,wdp_wdata_h_2x_22,wdp_wdata_h_2x_21,wdp_wdata_h_2x_20,wdp_wdata_h_2x_19,wdp_wdata_h_2x_18,wdp_wdata_h_2x_17,wdp_wdata_h_2x_16}),
	.dq_oe_2x_4(dq_oe_2x_4),
	.dq_oe_2x_5(dq_oe_2x_5),
	.dqs_output_data_out({\dqs_group[2].dq_dqs|wire_dqs_0_output_ddio_out_inst_dataout }),
	.bidir_dq_input_data_in({dq_datain_23,dq_datain_22,dq_datain_21,dq_datain_20,dq_datain_19,dq_datain_18,dq_datain_17,dq_datain_16}),
	.dqs_input_data_in({dqs_buffered_2}),
	.bidir_dq_0_oe_ff_inst1(bidir_dq_0_oe_ff_inst2),
	.bidir_dq_1_oe_ff_inst1(bidir_dq_1_oe_ff_inst2),
	.bidir_dq_2_oe_ff_inst1(bidir_dq_2_oe_ff_inst2),
	.bidir_dq_3_oe_ff_inst1(bidir_dq_3_oe_ff_inst2),
	.bidir_dq_4_oe_ff_inst1(bidir_dq_4_oe_ff_inst2),
	.bidir_dq_5_oe_ff_inst1(bidir_dq_5_oe_ff_inst2),
	.bidir_dq_6_oe_ff_inst1(bidir_dq_6_oe_ff_inst2),
	.bidir_dq_7_oe_ff_inst1(bidir_dq_7_oe_ff_inst2),
	.dqs_0_oe_ff_inst1(dqs_0_oe_ff_inst2),
	.dqsn_0_oe_ff_inst1(dqsn_0_oe_ff_inst2),
	.bidir_dq_areset({ams_pipe_3,ams_pipe_3,ams_pipe_3,ams_pipe_3,ams_pipe_3,ams_pipe_3,ams_pipe_3,ams_pipe_3}),
	.dqs_output_data_in_high({dqs_burst_2x_r3_2}),
	.dqs_enable_ctrl_in(postamble_en_pos_2x_2));

ddr3_int_ddr3_int_phy_alt_mem_phy_dq_dqs_3 \dqs_group[3].dq_dqs (
	.dqs_output_reg_clk(clk_1),
	.dq_output_reg_clk(clk_3),
	.dqs_enable_ctrl_clk(resync_clk_2x),
	.dll_delayctrlin({dqs_delay_ctrl_5,dqs_delay_ctrl_4,dqs_delay_ctrl_3,dqs_delay_ctrl_2,dqs_delay_ctrl_1,dqs_delay_ctrl_0}),
	.output_dq_output_data_out({wire_output_dq_0_output_ddio_out_inst_dataout3}),
	.output_dq_output_data_in_low({wdp_dm_l_2x_3}),
	.output_dq_output_data_in_high({wdp_dm_h_2x_3}),
	.bidir_dq_output_data_out({wire_bidir_dq_7_output_ddio_out_inst_dataout3,wire_bidir_dq_6_output_ddio_out_inst_dataout3,wire_bidir_dq_5_output_ddio_out_inst_dataout3,wire_bidir_dq_4_output_ddio_out_inst_dataout3,wire_bidir_dq_3_output_ddio_out_inst_dataout3,
wire_bidir_dq_2_output_ddio_out_inst_dataout3,wire_bidir_dq_1_output_ddio_out_inst_dataout3,wire_bidir_dq_0_output_ddio_out_inst_dataout3}),
	.bidir_dq_input_data_out_low({\dqs_group[3].dq_dqs|wire_bidir_dq_7_ddio_in_inst_regoutlo ,\dqs_group[3].dq_dqs|wire_bidir_dq_6_ddio_in_inst_regoutlo ,\dqs_group[3].dq_dqs|wire_bidir_dq_5_ddio_in_inst_regoutlo ,\dqs_group[3].dq_dqs|wire_bidir_dq_4_ddio_in_inst_regoutlo ,
\dqs_group[3].dq_dqs|wire_bidir_dq_3_ddio_in_inst_regoutlo ,\dqs_group[3].dq_dqs|wire_bidir_dq_2_ddio_in_inst_regoutlo ,\dqs_group[3].dq_dqs|wire_bidir_dq_1_ddio_in_inst_regoutlo ,\dqs_group[3].dq_dqs|wire_bidir_dq_0_ddio_in_inst_regoutlo }),
	.bidir_dq_input_data_out_high({\dqs_group[3].dq_dqs|wire_bidir_dq_7_ddio_in_inst_regouthi ,\dqs_group[3].dq_dqs|wire_bidir_dq_6_ddio_in_inst_regouthi ,\dqs_group[3].dq_dqs|wire_bidir_dq_5_ddio_in_inst_regouthi ,\dqs_group[3].dq_dqs|wire_bidir_dq_4_ddio_in_inst_regouthi ,
\dqs_group[3].dq_dqs|wire_bidir_dq_3_ddio_in_inst_regouthi ,\dqs_group[3].dq_dqs|wire_bidir_dq_2_ddio_in_inst_regouthi ,\dqs_group[3].dq_dqs|wire_bidir_dq_1_ddio_in_inst_regouthi ,\dqs_group[3].dq_dqs|wire_bidir_dq_0_ddio_in_inst_regouthi }),
	.bidir_dq_output_data_in_low({wdp_wdata_l_2x_31,wdp_wdata_l_2x_30,wdp_wdata_l_2x_29,wdp_wdata_l_2x_28,wdp_wdata_l_2x_27,wdp_wdata_l_2x_26,wdp_wdata_l_2x_25,wdp_wdata_l_2x_24}),
	.bidir_dq_output_data_in_high({wdp_wdata_h_2x_31,wdp_wdata_h_2x_30,wdp_wdata_h_2x_29,wdp_wdata_h_2x_28,wdp_wdata_h_2x_27,wdp_wdata_h_2x_26,wdp_wdata_h_2x_25,wdp_wdata_h_2x_24}),
	.dq_oe_2x_6(dq_oe_2x_6),
	.dq_oe_2x_7(dq_oe_2x_7),
	.dqs_output_data_out({\dqs_group[3].dq_dqs|wire_dqs_0_output_ddio_out_inst_dataout }),
	.bidir_dq_input_data_in({dq_datain_31,dq_datain_30,dq_datain_29,dq_datain_28,dq_datain_27,dq_datain_26,dq_datain_25,dq_datain_24}),
	.dqs_input_data_in({dqs_buffered_3}),
	.bidir_dq_0_oe_ff_inst1(bidir_dq_0_oe_ff_inst3),
	.bidir_dq_1_oe_ff_inst1(bidir_dq_1_oe_ff_inst3),
	.bidir_dq_2_oe_ff_inst1(bidir_dq_2_oe_ff_inst3),
	.bidir_dq_3_oe_ff_inst1(bidir_dq_3_oe_ff_inst3),
	.bidir_dq_4_oe_ff_inst1(bidir_dq_4_oe_ff_inst3),
	.bidir_dq_5_oe_ff_inst1(bidir_dq_5_oe_ff_inst3),
	.bidir_dq_6_oe_ff_inst1(bidir_dq_6_oe_ff_inst3),
	.bidir_dq_7_oe_ff_inst1(bidir_dq_7_oe_ff_inst3),
	.dqs_0_oe_ff_inst1(dqs_0_oe_ff_inst3),
	.dqsn_0_oe_ff_inst1(dqsn_0_oe_ff_inst3),
	.bidir_dq_areset({ams_pipe_3,ams_pipe_3,ams_pipe_3,ams_pipe_3,ams_pipe_3,ams_pipe_3,ams_pipe_3,ams_pipe_3}),
	.dqs_output_data_in_high({dqs_burst_2x_r3_3}),
	.dqs_enable_ctrl_in(postamble_en_pos_2x_3));

arriaii_pseudo_diff_out \dqs_group[0].ddr2_with_dqsn_buf_gen.dqs_pdiff_out (
	.i(\dqs_group[0].dq_dqs|wire_dqs_0_output_ddio_out_inst_dataout ),
	.o(dqs_pseudo_diff_out_0),
	.obar(dqsn_pseudo_diff_out_0));

arriaii_pseudo_diff_out \dqs_group[1].ddr2_with_dqsn_buf_gen.dqs_pdiff_out (
	.i(\dqs_group[1].dq_dqs|wire_dqs_0_output_ddio_out_inst_dataout ),
	.o(dqs_pseudo_diff_out_1),
	.obar(dqsn_pseudo_diff_out_1));

arriaii_pseudo_diff_out \dqs_group[2].ddr2_with_dqsn_buf_gen.dqs_pdiff_out (
	.i(\dqs_group[2].dq_dqs|wire_dqs_0_output_ddio_out_inst_dataout ),
	.o(dqs_pseudo_diff_out_2),
	.obar(dqsn_pseudo_diff_out_2));

arriaii_pseudo_diff_out \dqs_group[3].ddr2_with_dqsn_buf_gen.dqs_pdiff_out (
	.i(\dqs_group[3].dq_dqs|wire_dqs_0_output_ddio_out_inst_dataout ),
	.o(dqs_pseudo_diff_out_3),
	.obar(dqsn_pseudo_diff_out_3));

dffeas \dio_rdata_h_2x[0] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_h_2x[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_0),
	.prn(vcc));
defparam \dio_rdata_h_2x[0] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[0] .power_up = "low";

dffeas \dio_rdata_h_2x[1] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_h_2x[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_1),
	.prn(vcc));
defparam \dio_rdata_h_2x[1] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[1] .power_up = "low";

dffeas \dio_rdata_h_2x[2] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_h_2x[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_2),
	.prn(vcc));
defparam \dio_rdata_h_2x[2] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[2] .power_up = "low";

dffeas \dio_rdata_h_2x[3] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_h_2x[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_3),
	.prn(vcc));
defparam \dio_rdata_h_2x[3] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[3] .power_up = "low";

dffeas \dio_rdata_h_2x[4] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_h_2x[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_4),
	.prn(vcc));
defparam \dio_rdata_h_2x[4] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[4] .power_up = "low";

dffeas \dio_rdata_h_2x[5] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_h_2x[5]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_5),
	.prn(vcc));
defparam \dio_rdata_h_2x[5] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[5] .power_up = "low";

dffeas \dio_rdata_h_2x[6] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_h_2x[6]~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_6),
	.prn(vcc));
defparam \dio_rdata_h_2x[6] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[6] .power_up = "low";

dffeas \dio_rdata_h_2x[7] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_h_2x[7]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_7),
	.prn(vcc));
defparam \dio_rdata_h_2x[7] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[7] .power_up = "low";

dffeas \dio_rdata_h_2x[8] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_h_2x[8]~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_8),
	.prn(vcc));
defparam \dio_rdata_h_2x[8] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[8] .power_up = "low";

dffeas \dio_rdata_h_2x[9] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_h_2x[9]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_9),
	.prn(vcc));
defparam \dio_rdata_h_2x[9] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[9] .power_up = "low";

dffeas \dio_rdata_h_2x[10] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_h_2x[10]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_10),
	.prn(vcc));
defparam \dio_rdata_h_2x[10] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[10] .power_up = "low";

dffeas \dio_rdata_h_2x[11] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_h_2x[11]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_11),
	.prn(vcc));
defparam \dio_rdata_h_2x[11] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[11] .power_up = "low";

dffeas \dio_rdata_h_2x[12] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_h_2x[12]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_12),
	.prn(vcc));
defparam \dio_rdata_h_2x[12] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[12] .power_up = "low";

dffeas \dio_rdata_h_2x[13] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_h_2x[13]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_13),
	.prn(vcc));
defparam \dio_rdata_h_2x[13] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[13] .power_up = "low";

dffeas \dio_rdata_h_2x[14] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_h_2x[14]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_14),
	.prn(vcc));
defparam \dio_rdata_h_2x[14] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[14] .power_up = "low";

dffeas \dio_rdata_h_2x[15] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_h_2x[15]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_15),
	.prn(vcc));
defparam \dio_rdata_h_2x[15] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[15] .power_up = "low";

dffeas \dio_rdata_h_2x[16] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_h_2x[16]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_16),
	.prn(vcc));
defparam \dio_rdata_h_2x[16] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[16] .power_up = "low";

dffeas \dio_rdata_h_2x[17] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_h_2x[17]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_17),
	.prn(vcc));
defparam \dio_rdata_h_2x[17] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[17] .power_up = "low";

dffeas \dio_rdata_h_2x[18] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_h_2x[18]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_18),
	.prn(vcc));
defparam \dio_rdata_h_2x[18] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[18] .power_up = "low";

dffeas \dio_rdata_h_2x[19] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_h_2x[19]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_19),
	.prn(vcc));
defparam \dio_rdata_h_2x[19] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[19] .power_up = "low";

dffeas \dio_rdata_h_2x[20] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_h_2x[20]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_20),
	.prn(vcc));
defparam \dio_rdata_h_2x[20] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[20] .power_up = "low";

dffeas \dio_rdata_h_2x[21] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_h_2x[21]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_21),
	.prn(vcc));
defparam \dio_rdata_h_2x[21] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[21] .power_up = "low";

dffeas \dio_rdata_h_2x[22] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_h_2x[22]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_22),
	.prn(vcc));
defparam \dio_rdata_h_2x[22] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[22] .power_up = "low";

dffeas \dio_rdata_h_2x[23] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_h_2x[23]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_23),
	.prn(vcc));
defparam \dio_rdata_h_2x[23] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[23] .power_up = "low";

dffeas \dio_rdata_h_2x[24] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_h_2x[24]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_24),
	.prn(vcc));
defparam \dio_rdata_h_2x[24] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[24] .power_up = "low";

dffeas \dio_rdata_h_2x[25] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_h_2x[25]~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_25),
	.prn(vcc));
defparam \dio_rdata_h_2x[25] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[25] .power_up = "low";

dffeas \dio_rdata_h_2x[26] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_h_2x[26]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_26),
	.prn(vcc));
defparam \dio_rdata_h_2x[26] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[26] .power_up = "low";

dffeas \dio_rdata_h_2x[27] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_h_2x[27]~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_27),
	.prn(vcc));
defparam \dio_rdata_h_2x[27] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[27] .power_up = "low";

dffeas \dio_rdata_h_2x[28] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_h_2x[28]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_28),
	.prn(vcc));
defparam \dio_rdata_h_2x[28] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[28] .power_up = "low";

dffeas \dio_rdata_h_2x[29] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_h_2x[29]~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_29),
	.prn(vcc));
defparam \dio_rdata_h_2x[29] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[29] .power_up = "low";

dffeas \dio_rdata_h_2x[30] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_h_2x[30]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_30),
	.prn(vcc));
defparam \dio_rdata_h_2x[30] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[30] .power_up = "low";

dffeas \dio_rdata_h_2x[31] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_h_2x[31]~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_h_2x_31),
	.prn(vcc));
defparam \dio_rdata_h_2x[31] .is_wysiwyg = "true";
defparam \dio_rdata_h_2x[31] .power_up = "low";

dffeas \dio_rdata_l_2x[0] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_l_2x[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_0),
	.prn(vcc));
defparam \dio_rdata_l_2x[0] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[0] .power_up = "low";

dffeas \dio_rdata_l_2x[1] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_l_2x[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_1),
	.prn(vcc));
defparam \dio_rdata_l_2x[1] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[1] .power_up = "low";

dffeas \dio_rdata_l_2x[2] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_l_2x[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_2),
	.prn(vcc));
defparam \dio_rdata_l_2x[2] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[2] .power_up = "low";

dffeas \dio_rdata_l_2x[3] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_l_2x[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_3),
	.prn(vcc));
defparam \dio_rdata_l_2x[3] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[3] .power_up = "low";

dffeas \dio_rdata_l_2x[4] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_l_2x[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_4),
	.prn(vcc));
defparam \dio_rdata_l_2x[4] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[4] .power_up = "low";

dffeas \dio_rdata_l_2x[5] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_l_2x[5]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_5),
	.prn(vcc));
defparam \dio_rdata_l_2x[5] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[5] .power_up = "low";

dffeas \dio_rdata_l_2x[6] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_l_2x[6]~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_6),
	.prn(vcc));
defparam \dio_rdata_l_2x[6] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[6] .power_up = "low";

dffeas \dio_rdata_l_2x[7] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_l_2x[7]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_7),
	.prn(vcc));
defparam \dio_rdata_l_2x[7] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[7] .power_up = "low";

dffeas \dio_rdata_l_2x[8] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_l_2x[8]~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_8),
	.prn(vcc));
defparam \dio_rdata_l_2x[8] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[8] .power_up = "low";

dffeas \dio_rdata_l_2x[9] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_l_2x[9]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_9),
	.prn(vcc));
defparam \dio_rdata_l_2x[9] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[9] .power_up = "low";

dffeas \dio_rdata_l_2x[10] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_l_2x[10]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_10),
	.prn(vcc));
defparam \dio_rdata_l_2x[10] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[10] .power_up = "low";

dffeas \dio_rdata_l_2x[11] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_l_2x[11]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_11),
	.prn(vcc));
defparam \dio_rdata_l_2x[11] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[11] .power_up = "low";

dffeas \dio_rdata_l_2x[12] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_l_2x[12]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_12),
	.prn(vcc));
defparam \dio_rdata_l_2x[12] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[12] .power_up = "low";

dffeas \dio_rdata_l_2x[13] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_l_2x[13]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_13),
	.prn(vcc));
defparam \dio_rdata_l_2x[13] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[13] .power_up = "low";

dffeas \dio_rdata_l_2x[14] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_l_2x[14]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_14),
	.prn(vcc));
defparam \dio_rdata_l_2x[14] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[14] .power_up = "low";

dffeas \dio_rdata_l_2x[15] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_l_2x[15]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_15),
	.prn(vcc));
defparam \dio_rdata_l_2x[15] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[15] .power_up = "low";

dffeas \dio_rdata_l_2x[16] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_l_2x[16]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_16),
	.prn(vcc));
defparam \dio_rdata_l_2x[16] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[16] .power_up = "low";

dffeas \dio_rdata_l_2x[17] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_l_2x[17]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_17),
	.prn(vcc));
defparam \dio_rdata_l_2x[17] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[17] .power_up = "low";

dffeas \dio_rdata_l_2x[18] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_l_2x[18]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_18),
	.prn(vcc));
defparam \dio_rdata_l_2x[18] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[18] .power_up = "low";

dffeas \dio_rdata_l_2x[19] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_l_2x[19]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_19),
	.prn(vcc));
defparam \dio_rdata_l_2x[19] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[19] .power_up = "low";

dffeas \dio_rdata_l_2x[20] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_l_2x[20]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_20),
	.prn(vcc));
defparam \dio_rdata_l_2x[20] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[20] .power_up = "low";

dffeas \dio_rdata_l_2x[21] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_l_2x[21]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_21),
	.prn(vcc));
defparam \dio_rdata_l_2x[21] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[21] .power_up = "low";

dffeas \dio_rdata_l_2x[22] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_l_2x[22]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_22),
	.prn(vcc));
defparam \dio_rdata_l_2x[22] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[22] .power_up = "low";

dffeas \dio_rdata_l_2x[23] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_l_2x[23]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_23),
	.prn(vcc));
defparam \dio_rdata_l_2x[23] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[23] .power_up = "low";

dffeas \dio_rdata_l_2x[24] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_l_2x[24]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_24),
	.prn(vcc));
defparam \dio_rdata_l_2x[24] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[24] .power_up = "low";

dffeas \dio_rdata_l_2x[25] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_l_2x[25]~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_25),
	.prn(vcc));
defparam \dio_rdata_l_2x[25] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[25] .power_up = "low";

dffeas \dio_rdata_l_2x[26] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_l_2x[26]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_26),
	.prn(vcc));
defparam \dio_rdata_l_2x[26] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[26] .power_up = "low";

dffeas \dio_rdata_l_2x[27] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_l_2x[27]~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_27),
	.prn(vcc));
defparam \dio_rdata_l_2x[27] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[27] .power_up = "low";

dffeas \dio_rdata_l_2x[28] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_l_2x[28]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_28),
	.prn(vcc));
defparam \dio_rdata_l_2x[28] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[28] .power_up = "low";

dffeas \dio_rdata_l_2x[29] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_l_2x[29]~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_29),
	.prn(vcc));
defparam \dio_rdata_l_2x[29] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[29] .power_up = "low";

dffeas \dio_rdata_l_2x[30] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_l_2x[30]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_30),
	.prn(vcc));
defparam \dio_rdata_l_2x[30] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[30] .power_up = "low";

dffeas \dio_rdata_l_2x[31] (
	.clk(resync_clk_2x),
	.d(\dio_rdata_l_2x[31]~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dio_rdata_l_2x_31),
	.prn(vcc));
defparam \dio_rdata_l_2x[31] .is_wysiwyg = "true";
defparam \dio_rdata_l_2x[31] .power_up = "low";

arriaii_lcell_comb \rdata_p_ams[0]~0 (
	.dataa(!\dqs_group[0].dq_dqs|wire_bidir_dq_0_ddio_in_inst_regoutlo ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_p_ams[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_p_ams[0]~0 .extended_lut = "off";
defparam \rdata_p_ams[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_p_ams[0]~0 .shared_arith = "off";

dffeas \rdata_p_ams[0] (
	.clk(resync_clk_2x),
	.d(\rdata_p_ams[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[0]~q ),
	.prn(vcc));
defparam \rdata_p_ams[0] .is_wysiwyg = "true";
defparam \rdata_p_ams[0] .power_up = "low";

arriaii_lcell_comb \dio_rdata_h_2x[0]~0 (
	.dataa(!\rdata_p_ams[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_h_2x[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_h_2x[0]~0 .extended_lut = "off";
defparam \dio_rdata_h_2x[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_h_2x[0]~0 .shared_arith = "off";

arriaii_lcell_comb \rdata_p_ams[1]~1 (
	.dataa(!\dqs_group[0].dq_dqs|wire_bidir_dq_1_ddio_in_inst_regoutlo ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_p_ams[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_p_ams[1]~1 .extended_lut = "off";
defparam \rdata_p_ams[1]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_p_ams[1]~1 .shared_arith = "off";

dffeas \rdata_p_ams[1] (
	.clk(resync_clk_2x),
	.d(\rdata_p_ams[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[1]~q ),
	.prn(vcc));
defparam \rdata_p_ams[1] .is_wysiwyg = "true";
defparam \rdata_p_ams[1] .power_up = "low";

arriaii_lcell_comb \dio_rdata_h_2x[1]~1 (
	.dataa(!\rdata_p_ams[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_h_2x[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_h_2x[1]~1 .extended_lut = "off";
defparam \dio_rdata_h_2x[1]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_h_2x[1]~1 .shared_arith = "off";

arriaii_lcell_comb \rdata_p_ams[2]~2 (
	.dataa(!\dqs_group[0].dq_dqs|wire_bidir_dq_2_ddio_in_inst_regoutlo ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_p_ams[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_p_ams[2]~2 .extended_lut = "off";
defparam \rdata_p_ams[2]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_p_ams[2]~2 .shared_arith = "off";

dffeas \rdata_p_ams[2] (
	.clk(resync_clk_2x),
	.d(\rdata_p_ams[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[2]~q ),
	.prn(vcc));
defparam \rdata_p_ams[2] .is_wysiwyg = "true";
defparam \rdata_p_ams[2] .power_up = "low";

arriaii_lcell_comb \dio_rdata_h_2x[2]~2 (
	.dataa(!\rdata_p_ams[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_h_2x[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_h_2x[2]~2 .extended_lut = "off";
defparam \dio_rdata_h_2x[2]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_h_2x[2]~2 .shared_arith = "off";

arriaii_lcell_comb \rdata_p_ams[3]~3 (
	.dataa(!\dqs_group[0].dq_dqs|wire_bidir_dq_3_ddio_in_inst_regoutlo ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_p_ams[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_p_ams[3]~3 .extended_lut = "off";
defparam \rdata_p_ams[3]~3 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_p_ams[3]~3 .shared_arith = "off";

dffeas \rdata_p_ams[3] (
	.clk(resync_clk_2x),
	.d(\rdata_p_ams[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[3]~q ),
	.prn(vcc));
defparam \rdata_p_ams[3] .is_wysiwyg = "true";
defparam \rdata_p_ams[3] .power_up = "low";

arriaii_lcell_comb \dio_rdata_h_2x[3]~3 (
	.dataa(!\rdata_p_ams[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_h_2x[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_h_2x[3]~3 .extended_lut = "off";
defparam \dio_rdata_h_2x[3]~3 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_h_2x[3]~3 .shared_arith = "off";

arriaii_lcell_comb \rdata_p_ams[4]~4 (
	.dataa(!\dqs_group[0].dq_dqs|wire_bidir_dq_4_ddio_in_inst_regoutlo ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_p_ams[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_p_ams[4]~4 .extended_lut = "off";
defparam \rdata_p_ams[4]~4 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_p_ams[4]~4 .shared_arith = "off";

dffeas \rdata_p_ams[4] (
	.clk(resync_clk_2x),
	.d(\rdata_p_ams[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[4]~q ),
	.prn(vcc));
defparam \rdata_p_ams[4] .is_wysiwyg = "true";
defparam \rdata_p_ams[4] .power_up = "low";

arriaii_lcell_comb \dio_rdata_h_2x[4]~4 (
	.dataa(!\rdata_p_ams[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_h_2x[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_h_2x[4]~4 .extended_lut = "off";
defparam \dio_rdata_h_2x[4]~4 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_h_2x[4]~4 .shared_arith = "off";

arriaii_lcell_comb \rdata_p_ams[5]~5 (
	.dataa(!\dqs_group[0].dq_dqs|wire_bidir_dq_5_ddio_in_inst_regoutlo ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_p_ams[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_p_ams[5]~5 .extended_lut = "off";
defparam \rdata_p_ams[5]~5 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_p_ams[5]~5 .shared_arith = "off";

dffeas \rdata_p_ams[5] (
	.clk(resync_clk_2x),
	.d(\rdata_p_ams[5]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[5]~q ),
	.prn(vcc));
defparam \rdata_p_ams[5] .is_wysiwyg = "true";
defparam \rdata_p_ams[5] .power_up = "low";

arriaii_lcell_comb \dio_rdata_h_2x[5]~5 (
	.dataa(!\rdata_p_ams[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_h_2x[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_h_2x[5]~5 .extended_lut = "off";
defparam \dio_rdata_h_2x[5]~5 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_h_2x[5]~5 .shared_arith = "off";

arriaii_lcell_comb \rdata_p_ams[6]~6 (
	.dataa(!\dqs_group[0].dq_dqs|wire_bidir_dq_6_ddio_in_inst_regoutlo ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_p_ams[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_p_ams[6]~6 .extended_lut = "off";
defparam \rdata_p_ams[6]~6 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_p_ams[6]~6 .shared_arith = "off";

dffeas \rdata_p_ams[6] (
	.clk(resync_clk_2x),
	.d(\rdata_p_ams[6]~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[6]~q ),
	.prn(vcc));
defparam \rdata_p_ams[6] .is_wysiwyg = "true";
defparam \rdata_p_ams[6] .power_up = "low";

arriaii_lcell_comb \dio_rdata_h_2x[6]~6 (
	.dataa(!\rdata_p_ams[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_h_2x[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_h_2x[6]~6 .extended_lut = "off";
defparam \dio_rdata_h_2x[6]~6 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_h_2x[6]~6 .shared_arith = "off";

arriaii_lcell_comb \rdata_p_ams[7]~7 (
	.dataa(!\dqs_group[0].dq_dqs|wire_bidir_dq_7_ddio_in_inst_regoutlo ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_p_ams[7]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_p_ams[7]~7 .extended_lut = "off";
defparam \rdata_p_ams[7]~7 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_p_ams[7]~7 .shared_arith = "off";

dffeas \rdata_p_ams[7] (
	.clk(resync_clk_2x),
	.d(\rdata_p_ams[7]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[7]~q ),
	.prn(vcc));
defparam \rdata_p_ams[7] .is_wysiwyg = "true";
defparam \rdata_p_ams[7] .power_up = "low";

arriaii_lcell_comb \dio_rdata_h_2x[7]~7 (
	.dataa(!\rdata_p_ams[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_h_2x[7]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_h_2x[7]~7 .extended_lut = "off";
defparam \dio_rdata_h_2x[7]~7 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_h_2x[7]~7 .shared_arith = "off";

arriaii_lcell_comb \rdata_p_ams[8]~8 (
	.dataa(!\dqs_group[1].dq_dqs|wire_bidir_dq_0_ddio_in_inst_regoutlo ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_p_ams[8]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_p_ams[8]~8 .extended_lut = "off";
defparam \rdata_p_ams[8]~8 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_p_ams[8]~8 .shared_arith = "off";

dffeas \rdata_p_ams[8] (
	.clk(resync_clk_2x),
	.d(\rdata_p_ams[8]~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[8]~q ),
	.prn(vcc));
defparam \rdata_p_ams[8] .is_wysiwyg = "true";
defparam \rdata_p_ams[8] .power_up = "low";

arriaii_lcell_comb \dio_rdata_h_2x[8]~8 (
	.dataa(!\rdata_p_ams[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_h_2x[8]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_h_2x[8]~8 .extended_lut = "off";
defparam \dio_rdata_h_2x[8]~8 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_h_2x[8]~8 .shared_arith = "off";

arriaii_lcell_comb \rdata_p_ams[9]~9 (
	.dataa(!\dqs_group[1].dq_dqs|wire_bidir_dq_1_ddio_in_inst_regoutlo ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_p_ams[9]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_p_ams[9]~9 .extended_lut = "off";
defparam \rdata_p_ams[9]~9 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_p_ams[9]~9 .shared_arith = "off";

dffeas \rdata_p_ams[9] (
	.clk(resync_clk_2x),
	.d(\rdata_p_ams[9]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[9]~q ),
	.prn(vcc));
defparam \rdata_p_ams[9] .is_wysiwyg = "true";
defparam \rdata_p_ams[9] .power_up = "low";

arriaii_lcell_comb \dio_rdata_h_2x[9]~9 (
	.dataa(!\rdata_p_ams[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_h_2x[9]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_h_2x[9]~9 .extended_lut = "off";
defparam \dio_rdata_h_2x[9]~9 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_h_2x[9]~9 .shared_arith = "off";

arriaii_lcell_comb \rdata_p_ams[10]~10 (
	.dataa(!\dqs_group[1].dq_dqs|wire_bidir_dq_2_ddio_in_inst_regoutlo ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_p_ams[10]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_p_ams[10]~10 .extended_lut = "off";
defparam \rdata_p_ams[10]~10 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_p_ams[10]~10 .shared_arith = "off";

dffeas \rdata_p_ams[10] (
	.clk(resync_clk_2x),
	.d(\rdata_p_ams[10]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[10]~q ),
	.prn(vcc));
defparam \rdata_p_ams[10] .is_wysiwyg = "true";
defparam \rdata_p_ams[10] .power_up = "low";

arriaii_lcell_comb \dio_rdata_h_2x[10]~10 (
	.dataa(!\rdata_p_ams[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_h_2x[10]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_h_2x[10]~10 .extended_lut = "off";
defparam \dio_rdata_h_2x[10]~10 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_h_2x[10]~10 .shared_arith = "off";

arriaii_lcell_comb \rdata_p_ams[11]~11 (
	.dataa(!\dqs_group[1].dq_dqs|wire_bidir_dq_3_ddio_in_inst_regoutlo ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_p_ams[11]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_p_ams[11]~11 .extended_lut = "off";
defparam \rdata_p_ams[11]~11 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_p_ams[11]~11 .shared_arith = "off";

dffeas \rdata_p_ams[11] (
	.clk(resync_clk_2x),
	.d(\rdata_p_ams[11]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[11]~q ),
	.prn(vcc));
defparam \rdata_p_ams[11] .is_wysiwyg = "true";
defparam \rdata_p_ams[11] .power_up = "low";

arriaii_lcell_comb \dio_rdata_h_2x[11]~11 (
	.dataa(!\rdata_p_ams[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_h_2x[11]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_h_2x[11]~11 .extended_lut = "off";
defparam \dio_rdata_h_2x[11]~11 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_h_2x[11]~11 .shared_arith = "off";

arriaii_lcell_comb \rdata_p_ams[12]~12 (
	.dataa(!\dqs_group[1].dq_dqs|wire_bidir_dq_4_ddio_in_inst_regoutlo ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_p_ams[12]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_p_ams[12]~12 .extended_lut = "off";
defparam \rdata_p_ams[12]~12 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_p_ams[12]~12 .shared_arith = "off";

dffeas \rdata_p_ams[12] (
	.clk(resync_clk_2x),
	.d(\rdata_p_ams[12]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[12]~q ),
	.prn(vcc));
defparam \rdata_p_ams[12] .is_wysiwyg = "true";
defparam \rdata_p_ams[12] .power_up = "low";

arriaii_lcell_comb \dio_rdata_h_2x[12]~12 (
	.dataa(!\rdata_p_ams[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_h_2x[12]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_h_2x[12]~12 .extended_lut = "off";
defparam \dio_rdata_h_2x[12]~12 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_h_2x[12]~12 .shared_arith = "off";

arriaii_lcell_comb \rdata_p_ams[13]~13 (
	.dataa(!\dqs_group[1].dq_dqs|wire_bidir_dq_5_ddio_in_inst_regoutlo ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_p_ams[13]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_p_ams[13]~13 .extended_lut = "off";
defparam \rdata_p_ams[13]~13 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_p_ams[13]~13 .shared_arith = "off";

dffeas \rdata_p_ams[13] (
	.clk(resync_clk_2x),
	.d(\rdata_p_ams[13]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[13]~q ),
	.prn(vcc));
defparam \rdata_p_ams[13] .is_wysiwyg = "true";
defparam \rdata_p_ams[13] .power_up = "low";

arriaii_lcell_comb \dio_rdata_h_2x[13]~13 (
	.dataa(!\rdata_p_ams[13]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_h_2x[13]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_h_2x[13]~13 .extended_lut = "off";
defparam \dio_rdata_h_2x[13]~13 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_h_2x[13]~13 .shared_arith = "off";

arriaii_lcell_comb \rdata_p_ams[14]~14 (
	.dataa(!\dqs_group[1].dq_dqs|wire_bidir_dq_6_ddio_in_inst_regoutlo ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_p_ams[14]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_p_ams[14]~14 .extended_lut = "off";
defparam \rdata_p_ams[14]~14 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_p_ams[14]~14 .shared_arith = "off";

dffeas \rdata_p_ams[14] (
	.clk(resync_clk_2x),
	.d(\rdata_p_ams[14]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[14]~q ),
	.prn(vcc));
defparam \rdata_p_ams[14] .is_wysiwyg = "true";
defparam \rdata_p_ams[14] .power_up = "low";

arriaii_lcell_comb \dio_rdata_h_2x[14]~14 (
	.dataa(!\rdata_p_ams[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_h_2x[14]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_h_2x[14]~14 .extended_lut = "off";
defparam \dio_rdata_h_2x[14]~14 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_h_2x[14]~14 .shared_arith = "off";

arriaii_lcell_comb \rdata_p_ams[15]~15 (
	.dataa(!\dqs_group[1].dq_dqs|wire_bidir_dq_7_ddio_in_inst_regoutlo ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_p_ams[15]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_p_ams[15]~15 .extended_lut = "off";
defparam \rdata_p_ams[15]~15 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_p_ams[15]~15 .shared_arith = "off";

dffeas \rdata_p_ams[15] (
	.clk(resync_clk_2x),
	.d(\rdata_p_ams[15]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[15]~q ),
	.prn(vcc));
defparam \rdata_p_ams[15] .is_wysiwyg = "true";
defparam \rdata_p_ams[15] .power_up = "low";

arriaii_lcell_comb \dio_rdata_h_2x[15]~15 (
	.dataa(!\rdata_p_ams[15]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_h_2x[15]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_h_2x[15]~15 .extended_lut = "off";
defparam \dio_rdata_h_2x[15]~15 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_h_2x[15]~15 .shared_arith = "off";

arriaii_lcell_comb \rdata_p_ams[16]~16 (
	.dataa(!\dqs_group[2].dq_dqs|wire_bidir_dq_0_ddio_in_inst_regoutlo ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_p_ams[16]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_p_ams[16]~16 .extended_lut = "off";
defparam \rdata_p_ams[16]~16 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_p_ams[16]~16 .shared_arith = "off";

dffeas \rdata_p_ams[16] (
	.clk(resync_clk_2x),
	.d(\rdata_p_ams[16]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[16]~q ),
	.prn(vcc));
defparam \rdata_p_ams[16] .is_wysiwyg = "true";
defparam \rdata_p_ams[16] .power_up = "low";

arriaii_lcell_comb \dio_rdata_h_2x[16]~16 (
	.dataa(!\rdata_p_ams[16]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_h_2x[16]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_h_2x[16]~16 .extended_lut = "off";
defparam \dio_rdata_h_2x[16]~16 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_h_2x[16]~16 .shared_arith = "off";

arriaii_lcell_comb \rdata_p_ams[17]~17 (
	.dataa(!\dqs_group[2].dq_dqs|wire_bidir_dq_1_ddio_in_inst_regoutlo ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_p_ams[17]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_p_ams[17]~17 .extended_lut = "off";
defparam \rdata_p_ams[17]~17 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_p_ams[17]~17 .shared_arith = "off";

dffeas \rdata_p_ams[17] (
	.clk(resync_clk_2x),
	.d(\rdata_p_ams[17]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[17]~q ),
	.prn(vcc));
defparam \rdata_p_ams[17] .is_wysiwyg = "true";
defparam \rdata_p_ams[17] .power_up = "low";

arriaii_lcell_comb \dio_rdata_h_2x[17]~17 (
	.dataa(!\rdata_p_ams[17]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_h_2x[17]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_h_2x[17]~17 .extended_lut = "off";
defparam \dio_rdata_h_2x[17]~17 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_h_2x[17]~17 .shared_arith = "off";

arriaii_lcell_comb \rdata_p_ams[18]~18 (
	.dataa(!\dqs_group[2].dq_dqs|wire_bidir_dq_2_ddio_in_inst_regoutlo ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_p_ams[18]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_p_ams[18]~18 .extended_lut = "off";
defparam \rdata_p_ams[18]~18 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_p_ams[18]~18 .shared_arith = "off";

dffeas \rdata_p_ams[18] (
	.clk(resync_clk_2x),
	.d(\rdata_p_ams[18]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[18]~q ),
	.prn(vcc));
defparam \rdata_p_ams[18] .is_wysiwyg = "true";
defparam \rdata_p_ams[18] .power_up = "low";

arriaii_lcell_comb \dio_rdata_h_2x[18]~18 (
	.dataa(!\rdata_p_ams[18]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_h_2x[18]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_h_2x[18]~18 .extended_lut = "off";
defparam \dio_rdata_h_2x[18]~18 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_h_2x[18]~18 .shared_arith = "off";

arriaii_lcell_comb \rdata_p_ams[19]~19 (
	.dataa(!\dqs_group[2].dq_dqs|wire_bidir_dq_3_ddio_in_inst_regoutlo ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_p_ams[19]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_p_ams[19]~19 .extended_lut = "off";
defparam \rdata_p_ams[19]~19 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_p_ams[19]~19 .shared_arith = "off";

dffeas \rdata_p_ams[19] (
	.clk(resync_clk_2x),
	.d(\rdata_p_ams[19]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[19]~q ),
	.prn(vcc));
defparam \rdata_p_ams[19] .is_wysiwyg = "true";
defparam \rdata_p_ams[19] .power_up = "low";

arriaii_lcell_comb \dio_rdata_h_2x[19]~19 (
	.dataa(!\rdata_p_ams[19]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_h_2x[19]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_h_2x[19]~19 .extended_lut = "off";
defparam \dio_rdata_h_2x[19]~19 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_h_2x[19]~19 .shared_arith = "off";

arriaii_lcell_comb \rdata_p_ams[20]~20 (
	.dataa(!\dqs_group[2].dq_dqs|wire_bidir_dq_4_ddio_in_inst_regoutlo ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_p_ams[20]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_p_ams[20]~20 .extended_lut = "off";
defparam \rdata_p_ams[20]~20 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_p_ams[20]~20 .shared_arith = "off";

dffeas \rdata_p_ams[20] (
	.clk(resync_clk_2x),
	.d(\rdata_p_ams[20]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[20]~q ),
	.prn(vcc));
defparam \rdata_p_ams[20] .is_wysiwyg = "true";
defparam \rdata_p_ams[20] .power_up = "low";

arriaii_lcell_comb \dio_rdata_h_2x[20]~20 (
	.dataa(!\rdata_p_ams[20]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_h_2x[20]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_h_2x[20]~20 .extended_lut = "off";
defparam \dio_rdata_h_2x[20]~20 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_h_2x[20]~20 .shared_arith = "off";

arriaii_lcell_comb \rdata_p_ams[21]~21 (
	.dataa(!\dqs_group[2].dq_dqs|wire_bidir_dq_5_ddio_in_inst_regoutlo ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_p_ams[21]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_p_ams[21]~21 .extended_lut = "off";
defparam \rdata_p_ams[21]~21 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_p_ams[21]~21 .shared_arith = "off";

dffeas \rdata_p_ams[21] (
	.clk(resync_clk_2x),
	.d(\rdata_p_ams[21]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[21]~q ),
	.prn(vcc));
defparam \rdata_p_ams[21] .is_wysiwyg = "true";
defparam \rdata_p_ams[21] .power_up = "low";

arriaii_lcell_comb \dio_rdata_h_2x[21]~21 (
	.dataa(!\rdata_p_ams[21]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_h_2x[21]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_h_2x[21]~21 .extended_lut = "off";
defparam \dio_rdata_h_2x[21]~21 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_h_2x[21]~21 .shared_arith = "off";

arriaii_lcell_comb \rdata_p_ams[22]~22 (
	.dataa(!\dqs_group[2].dq_dqs|wire_bidir_dq_6_ddio_in_inst_regoutlo ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_p_ams[22]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_p_ams[22]~22 .extended_lut = "off";
defparam \rdata_p_ams[22]~22 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_p_ams[22]~22 .shared_arith = "off";

dffeas \rdata_p_ams[22] (
	.clk(resync_clk_2x),
	.d(\rdata_p_ams[22]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[22]~q ),
	.prn(vcc));
defparam \rdata_p_ams[22] .is_wysiwyg = "true";
defparam \rdata_p_ams[22] .power_up = "low";

arriaii_lcell_comb \dio_rdata_h_2x[22]~22 (
	.dataa(!\rdata_p_ams[22]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_h_2x[22]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_h_2x[22]~22 .extended_lut = "off";
defparam \dio_rdata_h_2x[22]~22 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_h_2x[22]~22 .shared_arith = "off";

arriaii_lcell_comb \rdata_p_ams[23]~23 (
	.dataa(!\dqs_group[2].dq_dqs|wire_bidir_dq_7_ddio_in_inst_regoutlo ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_p_ams[23]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_p_ams[23]~23 .extended_lut = "off";
defparam \rdata_p_ams[23]~23 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_p_ams[23]~23 .shared_arith = "off";

dffeas \rdata_p_ams[23] (
	.clk(resync_clk_2x),
	.d(\rdata_p_ams[23]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[23]~q ),
	.prn(vcc));
defparam \rdata_p_ams[23] .is_wysiwyg = "true";
defparam \rdata_p_ams[23] .power_up = "low";

arriaii_lcell_comb \dio_rdata_h_2x[23]~23 (
	.dataa(!\rdata_p_ams[23]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_h_2x[23]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_h_2x[23]~23 .extended_lut = "off";
defparam \dio_rdata_h_2x[23]~23 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_h_2x[23]~23 .shared_arith = "off";

arriaii_lcell_comb \rdata_p_ams[24]~24 (
	.dataa(!\dqs_group[3].dq_dqs|wire_bidir_dq_0_ddio_in_inst_regoutlo ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_p_ams[24]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_p_ams[24]~24 .extended_lut = "off";
defparam \rdata_p_ams[24]~24 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_p_ams[24]~24 .shared_arith = "off";

dffeas \rdata_p_ams[24] (
	.clk(resync_clk_2x),
	.d(\rdata_p_ams[24]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[24]~q ),
	.prn(vcc));
defparam \rdata_p_ams[24] .is_wysiwyg = "true";
defparam \rdata_p_ams[24] .power_up = "low";

arriaii_lcell_comb \dio_rdata_h_2x[24]~24 (
	.dataa(!\rdata_p_ams[24]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_h_2x[24]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_h_2x[24]~24 .extended_lut = "off";
defparam \dio_rdata_h_2x[24]~24 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_h_2x[24]~24 .shared_arith = "off";

arriaii_lcell_comb \rdata_p_ams[25]~25 (
	.dataa(!\dqs_group[3].dq_dqs|wire_bidir_dq_1_ddio_in_inst_regoutlo ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_p_ams[25]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_p_ams[25]~25 .extended_lut = "off";
defparam \rdata_p_ams[25]~25 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_p_ams[25]~25 .shared_arith = "off";

dffeas \rdata_p_ams[25] (
	.clk(resync_clk_2x),
	.d(\rdata_p_ams[25]~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[25]~q ),
	.prn(vcc));
defparam \rdata_p_ams[25] .is_wysiwyg = "true";
defparam \rdata_p_ams[25] .power_up = "low";

arriaii_lcell_comb \dio_rdata_h_2x[25]~25 (
	.dataa(!\rdata_p_ams[25]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_h_2x[25]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_h_2x[25]~25 .extended_lut = "off";
defparam \dio_rdata_h_2x[25]~25 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_h_2x[25]~25 .shared_arith = "off";

arriaii_lcell_comb \rdata_p_ams[26]~26 (
	.dataa(!\dqs_group[3].dq_dqs|wire_bidir_dq_2_ddio_in_inst_regoutlo ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_p_ams[26]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_p_ams[26]~26 .extended_lut = "off";
defparam \rdata_p_ams[26]~26 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_p_ams[26]~26 .shared_arith = "off";

dffeas \rdata_p_ams[26] (
	.clk(resync_clk_2x),
	.d(\rdata_p_ams[26]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[26]~q ),
	.prn(vcc));
defparam \rdata_p_ams[26] .is_wysiwyg = "true";
defparam \rdata_p_ams[26] .power_up = "low";

arriaii_lcell_comb \dio_rdata_h_2x[26]~26 (
	.dataa(!\rdata_p_ams[26]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_h_2x[26]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_h_2x[26]~26 .extended_lut = "off";
defparam \dio_rdata_h_2x[26]~26 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_h_2x[26]~26 .shared_arith = "off";

arriaii_lcell_comb \rdata_p_ams[27]~27 (
	.dataa(!\dqs_group[3].dq_dqs|wire_bidir_dq_3_ddio_in_inst_regoutlo ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_p_ams[27]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_p_ams[27]~27 .extended_lut = "off";
defparam \rdata_p_ams[27]~27 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_p_ams[27]~27 .shared_arith = "off";

dffeas \rdata_p_ams[27] (
	.clk(resync_clk_2x),
	.d(\rdata_p_ams[27]~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[27]~q ),
	.prn(vcc));
defparam \rdata_p_ams[27] .is_wysiwyg = "true";
defparam \rdata_p_ams[27] .power_up = "low";

arriaii_lcell_comb \dio_rdata_h_2x[27]~27 (
	.dataa(!\rdata_p_ams[27]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_h_2x[27]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_h_2x[27]~27 .extended_lut = "off";
defparam \dio_rdata_h_2x[27]~27 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_h_2x[27]~27 .shared_arith = "off";

arriaii_lcell_comb \rdata_p_ams[28]~28 (
	.dataa(!\dqs_group[3].dq_dqs|wire_bidir_dq_4_ddio_in_inst_regoutlo ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_p_ams[28]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_p_ams[28]~28 .extended_lut = "off";
defparam \rdata_p_ams[28]~28 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_p_ams[28]~28 .shared_arith = "off";

dffeas \rdata_p_ams[28] (
	.clk(resync_clk_2x),
	.d(\rdata_p_ams[28]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[28]~q ),
	.prn(vcc));
defparam \rdata_p_ams[28] .is_wysiwyg = "true";
defparam \rdata_p_ams[28] .power_up = "low";

arriaii_lcell_comb \dio_rdata_h_2x[28]~28 (
	.dataa(!\rdata_p_ams[28]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_h_2x[28]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_h_2x[28]~28 .extended_lut = "off";
defparam \dio_rdata_h_2x[28]~28 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_h_2x[28]~28 .shared_arith = "off";

arriaii_lcell_comb \rdata_p_ams[29]~29 (
	.dataa(!\dqs_group[3].dq_dqs|wire_bidir_dq_5_ddio_in_inst_regoutlo ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_p_ams[29]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_p_ams[29]~29 .extended_lut = "off";
defparam \rdata_p_ams[29]~29 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_p_ams[29]~29 .shared_arith = "off";

dffeas \rdata_p_ams[29] (
	.clk(resync_clk_2x),
	.d(\rdata_p_ams[29]~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[29]~q ),
	.prn(vcc));
defparam \rdata_p_ams[29] .is_wysiwyg = "true";
defparam \rdata_p_ams[29] .power_up = "low";

arriaii_lcell_comb \dio_rdata_h_2x[29]~29 (
	.dataa(!\rdata_p_ams[29]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_h_2x[29]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_h_2x[29]~29 .extended_lut = "off";
defparam \dio_rdata_h_2x[29]~29 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_h_2x[29]~29 .shared_arith = "off";

arriaii_lcell_comb \rdata_p_ams[30]~30 (
	.dataa(!\dqs_group[3].dq_dqs|wire_bidir_dq_6_ddio_in_inst_regoutlo ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_p_ams[30]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_p_ams[30]~30 .extended_lut = "off";
defparam \rdata_p_ams[30]~30 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_p_ams[30]~30 .shared_arith = "off";

dffeas \rdata_p_ams[30] (
	.clk(resync_clk_2x),
	.d(\rdata_p_ams[30]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[30]~q ),
	.prn(vcc));
defparam \rdata_p_ams[30] .is_wysiwyg = "true";
defparam \rdata_p_ams[30] .power_up = "low";

arriaii_lcell_comb \dio_rdata_h_2x[30]~30 (
	.dataa(!\rdata_p_ams[30]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_h_2x[30]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_h_2x[30]~30 .extended_lut = "off";
defparam \dio_rdata_h_2x[30]~30 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_h_2x[30]~30 .shared_arith = "off";

arriaii_lcell_comb \rdata_p_ams[31]~31 (
	.dataa(!\dqs_group[3].dq_dqs|wire_bidir_dq_7_ddio_in_inst_regoutlo ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_p_ams[31]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_p_ams[31]~31 .extended_lut = "off";
defparam \rdata_p_ams[31]~31 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_p_ams[31]~31 .shared_arith = "off";

dffeas \rdata_p_ams[31] (
	.clk(resync_clk_2x),
	.d(\rdata_p_ams[31]~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_p_ams[31]~q ),
	.prn(vcc));
defparam \rdata_p_ams[31] .is_wysiwyg = "true";
defparam \rdata_p_ams[31] .power_up = "low";

arriaii_lcell_comb \dio_rdata_h_2x[31]~31 (
	.dataa(!\rdata_p_ams[31]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_h_2x[31]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_h_2x[31]~31 .extended_lut = "off";
defparam \dio_rdata_h_2x[31]~31 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_h_2x[31]~31 .shared_arith = "off";

arriaii_lcell_comb \rdata_n_ams[0]~0 (
	.dataa(!\dqs_group[0].dq_dqs|wire_bidir_dq_0_ddio_in_inst_regouthi ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_n_ams[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_n_ams[0]~0 .extended_lut = "off";
defparam \rdata_n_ams[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_n_ams[0]~0 .shared_arith = "off";

dffeas \rdata_n_ams[0] (
	.clk(resync_clk_2x),
	.d(\rdata_n_ams[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[0]~q ),
	.prn(vcc));
defparam \rdata_n_ams[0] .is_wysiwyg = "true";
defparam \rdata_n_ams[0] .power_up = "low";

arriaii_lcell_comb \dio_rdata_l_2x[0]~0 (
	.dataa(!\rdata_n_ams[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_l_2x[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_l_2x[0]~0 .extended_lut = "off";
defparam \dio_rdata_l_2x[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_l_2x[0]~0 .shared_arith = "off";

arriaii_lcell_comb \rdata_n_ams[1]~1 (
	.dataa(!\dqs_group[0].dq_dqs|wire_bidir_dq_1_ddio_in_inst_regouthi ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_n_ams[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_n_ams[1]~1 .extended_lut = "off";
defparam \rdata_n_ams[1]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_n_ams[1]~1 .shared_arith = "off";

dffeas \rdata_n_ams[1] (
	.clk(resync_clk_2x),
	.d(\rdata_n_ams[1]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[1]~q ),
	.prn(vcc));
defparam \rdata_n_ams[1] .is_wysiwyg = "true";
defparam \rdata_n_ams[1] .power_up = "low";

arriaii_lcell_comb \dio_rdata_l_2x[1]~1 (
	.dataa(!\rdata_n_ams[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_l_2x[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_l_2x[1]~1 .extended_lut = "off";
defparam \dio_rdata_l_2x[1]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_l_2x[1]~1 .shared_arith = "off";

arriaii_lcell_comb \rdata_n_ams[2]~2 (
	.dataa(!\dqs_group[0].dq_dqs|wire_bidir_dq_2_ddio_in_inst_regouthi ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_n_ams[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_n_ams[2]~2 .extended_lut = "off";
defparam \rdata_n_ams[2]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_n_ams[2]~2 .shared_arith = "off";

dffeas \rdata_n_ams[2] (
	.clk(resync_clk_2x),
	.d(\rdata_n_ams[2]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[2]~q ),
	.prn(vcc));
defparam \rdata_n_ams[2] .is_wysiwyg = "true";
defparam \rdata_n_ams[2] .power_up = "low";

arriaii_lcell_comb \dio_rdata_l_2x[2]~2 (
	.dataa(!\rdata_n_ams[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_l_2x[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_l_2x[2]~2 .extended_lut = "off";
defparam \dio_rdata_l_2x[2]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_l_2x[2]~2 .shared_arith = "off";

arriaii_lcell_comb \rdata_n_ams[3]~3 (
	.dataa(!\dqs_group[0].dq_dqs|wire_bidir_dq_3_ddio_in_inst_regouthi ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_n_ams[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_n_ams[3]~3 .extended_lut = "off";
defparam \rdata_n_ams[3]~3 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_n_ams[3]~3 .shared_arith = "off";

dffeas \rdata_n_ams[3] (
	.clk(resync_clk_2x),
	.d(\rdata_n_ams[3]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[3]~q ),
	.prn(vcc));
defparam \rdata_n_ams[3] .is_wysiwyg = "true";
defparam \rdata_n_ams[3] .power_up = "low";

arriaii_lcell_comb \dio_rdata_l_2x[3]~3 (
	.dataa(!\rdata_n_ams[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_l_2x[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_l_2x[3]~3 .extended_lut = "off";
defparam \dio_rdata_l_2x[3]~3 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_l_2x[3]~3 .shared_arith = "off";

arriaii_lcell_comb \rdata_n_ams[4]~4 (
	.dataa(!\dqs_group[0].dq_dqs|wire_bidir_dq_4_ddio_in_inst_regouthi ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_n_ams[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_n_ams[4]~4 .extended_lut = "off";
defparam \rdata_n_ams[4]~4 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_n_ams[4]~4 .shared_arith = "off";

dffeas \rdata_n_ams[4] (
	.clk(resync_clk_2x),
	.d(\rdata_n_ams[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[4]~q ),
	.prn(vcc));
defparam \rdata_n_ams[4] .is_wysiwyg = "true";
defparam \rdata_n_ams[4] .power_up = "low";

arriaii_lcell_comb \dio_rdata_l_2x[4]~4 (
	.dataa(!\rdata_n_ams[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_l_2x[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_l_2x[4]~4 .extended_lut = "off";
defparam \dio_rdata_l_2x[4]~4 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_l_2x[4]~4 .shared_arith = "off";

arriaii_lcell_comb \rdata_n_ams[5]~5 (
	.dataa(!\dqs_group[0].dq_dqs|wire_bidir_dq_5_ddio_in_inst_regouthi ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_n_ams[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_n_ams[5]~5 .extended_lut = "off";
defparam \rdata_n_ams[5]~5 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_n_ams[5]~5 .shared_arith = "off";

dffeas \rdata_n_ams[5] (
	.clk(resync_clk_2x),
	.d(\rdata_n_ams[5]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[5]~q ),
	.prn(vcc));
defparam \rdata_n_ams[5] .is_wysiwyg = "true";
defparam \rdata_n_ams[5] .power_up = "low";

arriaii_lcell_comb \dio_rdata_l_2x[5]~5 (
	.dataa(!\rdata_n_ams[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_l_2x[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_l_2x[5]~5 .extended_lut = "off";
defparam \dio_rdata_l_2x[5]~5 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_l_2x[5]~5 .shared_arith = "off";

arriaii_lcell_comb \rdata_n_ams[6]~6 (
	.dataa(!\dqs_group[0].dq_dqs|wire_bidir_dq_6_ddio_in_inst_regouthi ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_n_ams[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_n_ams[6]~6 .extended_lut = "off";
defparam \rdata_n_ams[6]~6 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_n_ams[6]~6 .shared_arith = "off";

dffeas \rdata_n_ams[6] (
	.clk(resync_clk_2x),
	.d(\rdata_n_ams[6]~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[6]~q ),
	.prn(vcc));
defparam \rdata_n_ams[6] .is_wysiwyg = "true";
defparam \rdata_n_ams[6] .power_up = "low";

arriaii_lcell_comb \dio_rdata_l_2x[6]~6 (
	.dataa(!\rdata_n_ams[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_l_2x[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_l_2x[6]~6 .extended_lut = "off";
defparam \dio_rdata_l_2x[6]~6 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_l_2x[6]~6 .shared_arith = "off";

arriaii_lcell_comb \rdata_n_ams[7]~7 (
	.dataa(!\dqs_group[0].dq_dqs|wire_bidir_dq_7_ddio_in_inst_regouthi ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_n_ams[7]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_n_ams[7]~7 .extended_lut = "off";
defparam \rdata_n_ams[7]~7 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_n_ams[7]~7 .shared_arith = "off";

dffeas \rdata_n_ams[7] (
	.clk(resync_clk_2x),
	.d(\rdata_n_ams[7]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[7]~q ),
	.prn(vcc));
defparam \rdata_n_ams[7] .is_wysiwyg = "true";
defparam \rdata_n_ams[7] .power_up = "low";

arriaii_lcell_comb \dio_rdata_l_2x[7]~7 (
	.dataa(!\rdata_n_ams[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_l_2x[7]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_l_2x[7]~7 .extended_lut = "off";
defparam \dio_rdata_l_2x[7]~7 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_l_2x[7]~7 .shared_arith = "off";

arriaii_lcell_comb \rdata_n_ams[8]~8 (
	.dataa(!\dqs_group[1].dq_dqs|wire_bidir_dq_0_ddio_in_inst_regouthi ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_n_ams[8]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_n_ams[8]~8 .extended_lut = "off";
defparam \rdata_n_ams[8]~8 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_n_ams[8]~8 .shared_arith = "off";

dffeas \rdata_n_ams[8] (
	.clk(resync_clk_2x),
	.d(\rdata_n_ams[8]~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[8]~q ),
	.prn(vcc));
defparam \rdata_n_ams[8] .is_wysiwyg = "true";
defparam \rdata_n_ams[8] .power_up = "low";

arriaii_lcell_comb \dio_rdata_l_2x[8]~8 (
	.dataa(!\rdata_n_ams[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_l_2x[8]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_l_2x[8]~8 .extended_lut = "off";
defparam \dio_rdata_l_2x[8]~8 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_l_2x[8]~8 .shared_arith = "off";

arriaii_lcell_comb \rdata_n_ams[9]~9 (
	.dataa(!\dqs_group[1].dq_dqs|wire_bidir_dq_1_ddio_in_inst_regouthi ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_n_ams[9]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_n_ams[9]~9 .extended_lut = "off";
defparam \rdata_n_ams[9]~9 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_n_ams[9]~9 .shared_arith = "off";

dffeas \rdata_n_ams[9] (
	.clk(resync_clk_2x),
	.d(\rdata_n_ams[9]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[9]~q ),
	.prn(vcc));
defparam \rdata_n_ams[9] .is_wysiwyg = "true";
defparam \rdata_n_ams[9] .power_up = "low";

arriaii_lcell_comb \dio_rdata_l_2x[9]~9 (
	.dataa(!\rdata_n_ams[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_l_2x[9]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_l_2x[9]~9 .extended_lut = "off";
defparam \dio_rdata_l_2x[9]~9 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_l_2x[9]~9 .shared_arith = "off";

arriaii_lcell_comb \rdata_n_ams[10]~10 (
	.dataa(!\dqs_group[1].dq_dqs|wire_bidir_dq_2_ddio_in_inst_regouthi ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_n_ams[10]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_n_ams[10]~10 .extended_lut = "off";
defparam \rdata_n_ams[10]~10 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_n_ams[10]~10 .shared_arith = "off";

dffeas \rdata_n_ams[10] (
	.clk(resync_clk_2x),
	.d(\rdata_n_ams[10]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[10]~q ),
	.prn(vcc));
defparam \rdata_n_ams[10] .is_wysiwyg = "true";
defparam \rdata_n_ams[10] .power_up = "low";

arriaii_lcell_comb \dio_rdata_l_2x[10]~10 (
	.dataa(!\rdata_n_ams[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_l_2x[10]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_l_2x[10]~10 .extended_lut = "off";
defparam \dio_rdata_l_2x[10]~10 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_l_2x[10]~10 .shared_arith = "off";

arriaii_lcell_comb \rdata_n_ams[11]~11 (
	.dataa(!\dqs_group[1].dq_dqs|wire_bidir_dq_3_ddio_in_inst_regouthi ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_n_ams[11]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_n_ams[11]~11 .extended_lut = "off";
defparam \rdata_n_ams[11]~11 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_n_ams[11]~11 .shared_arith = "off";

dffeas \rdata_n_ams[11] (
	.clk(resync_clk_2x),
	.d(\rdata_n_ams[11]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[11]~q ),
	.prn(vcc));
defparam \rdata_n_ams[11] .is_wysiwyg = "true";
defparam \rdata_n_ams[11] .power_up = "low";

arriaii_lcell_comb \dio_rdata_l_2x[11]~11 (
	.dataa(!\rdata_n_ams[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_l_2x[11]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_l_2x[11]~11 .extended_lut = "off";
defparam \dio_rdata_l_2x[11]~11 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_l_2x[11]~11 .shared_arith = "off";

arriaii_lcell_comb \rdata_n_ams[12]~12 (
	.dataa(!\dqs_group[1].dq_dqs|wire_bidir_dq_4_ddio_in_inst_regouthi ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_n_ams[12]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_n_ams[12]~12 .extended_lut = "off";
defparam \rdata_n_ams[12]~12 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_n_ams[12]~12 .shared_arith = "off";

dffeas \rdata_n_ams[12] (
	.clk(resync_clk_2x),
	.d(\rdata_n_ams[12]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[12]~q ),
	.prn(vcc));
defparam \rdata_n_ams[12] .is_wysiwyg = "true";
defparam \rdata_n_ams[12] .power_up = "low";

arriaii_lcell_comb \dio_rdata_l_2x[12]~12 (
	.dataa(!\rdata_n_ams[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_l_2x[12]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_l_2x[12]~12 .extended_lut = "off";
defparam \dio_rdata_l_2x[12]~12 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_l_2x[12]~12 .shared_arith = "off";

arriaii_lcell_comb \rdata_n_ams[13]~13 (
	.dataa(!\dqs_group[1].dq_dqs|wire_bidir_dq_5_ddio_in_inst_regouthi ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_n_ams[13]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_n_ams[13]~13 .extended_lut = "off";
defparam \rdata_n_ams[13]~13 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_n_ams[13]~13 .shared_arith = "off";

dffeas \rdata_n_ams[13] (
	.clk(resync_clk_2x),
	.d(\rdata_n_ams[13]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[13]~q ),
	.prn(vcc));
defparam \rdata_n_ams[13] .is_wysiwyg = "true";
defparam \rdata_n_ams[13] .power_up = "low";

arriaii_lcell_comb \dio_rdata_l_2x[13]~13 (
	.dataa(!\rdata_n_ams[13]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_l_2x[13]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_l_2x[13]~13 .extended_lut = "off";
defparam \dio_rdata_l_2x[13]~13 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_l_2x[13]~13 .shared_arith = "off";

arriaii_lcell_comb \rdata_n_ams[14]~14 (
	.dataa(!\dqs_group[1].dq_dqs|wire_bidir_dq_6_ddio_in_inst_regouthi ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_n_ams[14]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_n_ams[14]~14 .extended_lut = "off";
defparam \rdata_n_ams[14]~14 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_n_ams[14]~14 .shared_arith = "off";

dffeas \rdata_n_ams[14] (
	.clk(resync_clk_2x),
	.d(\rdata_n_ams[14]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[14]~q ),
	.prn(vcc));
defparam \rdata_n_ams[14] .is_wysiwyg = "true";
defparam \rdata_n_ams[14] .power_up = "low";

arriaii_lcell_comb \dio_rdata_l_2x[14]~14 (
	.dataa(!\rdata_n_ams[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_l_2x[14]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_l_2x[14]~14 .extended_lut = "off";
defparam \dio_rdata_l_2x[14]~14 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_l_2x[14]~14 .shared_arith = "off";

arriaii_lcell_comb \rdata_n_ams[15]~15 (
	.dataa(!\dqs_group[1].dq_dqs|wire_bidir_dq_7_ddio_in_inst_regouthi ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_n_ams[15]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_n_ams[15]~15 .extended_lut = "off";
defparam \rdata_n_ams[15]~15 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_n_ams[15]~15 .shared_arith = "off";

dffeas \rdata_n_ams[15] (
	.clk(resync_clk_2x),
	.d(\rdata_n_ams[15]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[15]~q ),
	.prn(vcc));
defparam \rdata_n_ams[15] .is_wysiwyg = "true";
defparam \rdata_n_ams[15] .power_up = "low";

arriaii_lcell_comb \dio_rdata_l_2x[15]~15 (
	.dataa(!\rdata_n_ams[15]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_l_2x[15]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_l_2x[15]~15 .extended_lut = "off";
defparam \dio_rdata_l_2x[15]~15 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_l_2x[15]~15 .shared_arith = "off";

arriaii_lcell_comb \rdata_n_ams[16]~16 (
	.dataa(!\dqs_group[2].dq_dqs|wire_bidir_dq_0_ddio_in_inst_regouthi ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_n_ams[16]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_n_ams[16]~16 .extended_lut = "off";
defparam \rdata_n_ams[16]~16 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_n_ams[16]~16 .shared_arith = "off";

dffeas \rdata_n_ams[16] (
	.clk(resync_clk_2x),
	.d(\rdata_n_ams[16]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[16]~q ),
	.prn(vcc));
defparam \rdata_n_ams[16] .is_wysiwyg = "true";
defparam \rdata_n_ams[16] .power_up = "low";

arriaii_lcell_comb \dio_rdata_l_2x[16]~16 (
	.dataa(!\rdata_n_ams[16]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_l_2x[16]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_l_2x[16]~16 .extended_lut = "off";
defparam \dio_rdata_l_2x[16]~16 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_l_2x[16]~16 .shared_arith = "off";

arriaii_lcell_comb \rdata_n_ams[17]~17 (
	.dataa(!\dqs_group[2].dq_dqs|wire_bidir_dq_1_ddio_in_inst_regouthi ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_n_ams[17]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_n_ams[17]~17 .extended_lut = "off";
defparam \rdata_n_ams[17]~17 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_n_ams[17]~17 .shared_arith = "off";

dffeas \rdata_n_ams[17] (
	.clk(resync_clk_2x),
	.d(\rdata_n_ams[17]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[17]~q ),
	.prn(vcc));
defparam \rdata_n_ams[17] .is_wysiwyg = "true";
defparam \rdata_n_ams[17] .power_up = "low";

arriaii_lcell_comb \dio_rdata_l_2x[17]~17 (
	.dataa(!\rdata_n_ams[17]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_l_2x[17]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_l_2x[17]~17 .extended_lut = "off";
defparam \dio_rdata_l_2x[17]~17 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_l_2x[17]~17 .shared_arith = "off";

arriaii_lcell_comb \rdata_n_ams[18]~18 (
	.dataa(!\dqs_group[2].dq_dqs|wire_bidir_dq_2_ddio_in_inst_regouthi ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_n_ams[18]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_n_ams[18]~18 .extended_lut = "off";
defparam \rdata_n_ams[18]~18 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_n_ams[18]~18 .shared_arith = "off";

dffeas \rdata_n_ams[18] (
	.clk(resync_clk_2x),
	.d(\rdata_n_ams[18]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[18]~q ),
	.prn(vcc));
defparam \rdata_n_ams[18] .is_wysiwyg = "true";
defparam \rdata_n_ams[18] .power_up = "low";

arriaii_lcell_comb \dio_rdata_l_2x[18]~18 (
	.dataa(!\rdata_n_ams[18]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_l_2x[18]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_l_2x[18]~18 .extended_lut = "off";
defparam \dio_rdata_l_2x[18]~18 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_l_2x[18]~18 .shared_arith = "off";

arriaii_lcell_comb \rdata_n_ams[19]~19 (
	.dataa(!\dqs_group[2].dq_dqs|wire_bidir_dq_3_ddio_in_inst_regouthi ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_n_ams[19]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_n_ams[19]~19 .extended_lut = "off";
defparam \rdata_n_ams[19]~19 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_n_ams[19]~19 .shared_arith = "off";

dffeas \rdata_n_ams[19] (
	.clk(resync_clk_2x),
	.d(\rdata_n_ams[19]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[19]~q ),
	.prn(vcc));
defparam \rdata_n_ams[19] .is_wysiwyg = "true";
defparam \rdata_n_ams[19] .power_up = "low";

arriaii_lcell_comb \dio_rdata_l_2x[19]~19 (
	.dataa(!\rdata_n_ams[19]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_l_2x[19]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_l_2x[19]~19 .extended_lut = "off";
defparam \dio_rdata_l_2x[19]~19 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_l_2x[19]~19 .shared_arith = "off";

arriaii_lcell_comb \rdata_n_ams[20]~20 (
	.dataa(!\dqs_group[2].dq_dqs|wire_bidir_dq_4_ddio_in_inst_regouthi ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_n_ams[20]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_n_ams[20]~20 .extended_lut = "off";
defparam \rdata_n_ams[20]~20 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_n_ams[20]~20 .shared_arith = "off";

dffeas \rdata_n_ams[20] (
	.clk(resync_clk_2x),
	.d(\rdata_n_ams[20]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[20]~q ),
	.prn(vcc));
defparam \rdata_n_ams[20] .is_wysiwyg = "true";
defparam \rdata_n_ams[20] .power_up = "low";

arriaii_lcell_comb \dio_rdata_l_2x[20]~20 (
	.dataa(!\rdata_n_ams[20]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_l_2x[20]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_l_2x[20]~20 .extended_lut = "off";
defparam \dio_rdata_l_2x[20]~20 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_l_2x[20]~20 .shared_arith = "off";

arriaii_lcell_comb \rdata_n_ams[21]~21 (
	.dataa(!\dqs_group[2].dq_dqs|wire_bidir_dq_5_ddio_in_inst_regouthi ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_n_ams[21]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_n_ams[21]~21 .extended_lut = "off";
defparam \rdata_n_ams[21]~21 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_n_ams[21]~21 .shared_arith = "off";

dffeas \rdata_n_ams[21] (
	.clk(resync_clk_2x),
	.d(\rdata_n_ams[21]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[21]~q ),
	.prn(vcc));
defparam \rdata_n_ams[21] .is_wysiwyg = "true";
defparam \rdata_n_ams[21] .power_up = "low";

arriaii_lcell_comb \dio_rdata_l_2x[21]~21 (
	.dataa(!\rdata_n_ams[21]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_l_2x[21]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_l_2x[21]~21 .extended_lut = "off";
defparam \dio_rdata_l_2x[21]~21 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_l_2x[21]~21 .shared_arith = "off";

arriaii_lcell_comb \rdata_n_ams[22]~22 (
	.dataa(!\dqs_group[2].dq_dqs|wire_bidir_dq_6_ddio_in_inst_regouthi ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_n_ams[22]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_n_ams[22]~22 .extended_lut = "off";
defparam \rdata_n_ams[22]~22 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_n_ams[22]~22 .shared_arith = "off";

dffeas \rdata_n_ams[22] (
	.clk(resync_clk_2x),
	.d(\rdata_n_ams[22]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[22]~q ),
	.prn(vcc));
defparam \rdata_n_ams[22] .is_wysiwyg = "true";
defparam \rdata_n_ams[22] .power_up = "low";

arriaii_lcell_comb \dio_rdata_l_2x[22]~22 (
	.dataa(!\rdata_n_ams[22]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_l_2x[22]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_l_2x[22]~22 .extended_lut = "off";
defparam \dio_rdata_l_2x[22]~22 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_l_2x[22]~22 .shared_arith = "off";

arriaii_lcell_comb \rdata_n_ams[23]~23 (
	.dataa(!\dqs_group[2].dq_dqs|wire_bidir_dq_7_ddio_in_inst_regouthi ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_n_ams[23]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_n_ams[23]~23 .extended_lut = "off";
defparam \rdata_n_ams[23]~23 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_n_ams[23]~23 .shared_arith = "off";

dffeas \rdata_n_ams[23] (
	.clk(resync_clk_2x),
	.d(\rdata_n_ams[23]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[23]~q ),
	.prn(vcc));
defparam \rdata_n_ams[23] .is_wysiwyg = "true";
defparam \rdata_n_ams[23] .power_up = "low";

arriaii_lcell_comb \dio_rdata_l_2x[23]~23 (
	.dataa(!\rdata_n_ams[23]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_l_2x[23]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_l_2x[23]~23 .extended_lut = "off";
defparam \dio_rdata_l_2x[23]~23 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_l_2x[23]~23 .shared_arith = "off";

arriaii_lcell_comb \rdata_n_ams[24]~24 (
	.dataa(!\dqs_group[3].dq_dqs|wire_bidir_dq_0_ddio_in_inst_regouthi ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_n_ams[24]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_n_ams[24]~24 .extended_lut = "off";
defparam \rdata_n_ams[24]~24 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_n_ams[24]~24 .shared_arith = "off";

dffeas \rdata_n_ams[24] (
	.clk(resync_clk_2x),
	.d(\rdata_n_ams[24]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[24]~q ),
	.prn(vcc));
defparam \rdata_n_ams[24] .is_wysiwyg = "true";
defparam \rdata_n_ams[24] .power_up = "low";

arriaii_lcell_comb \dio_rdata_l_2x[24]~24 (
	.dataa(!\rdata_n_ams[24]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_l_2x[24]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_l_2x[24]~24 .extended_lut = "off";
defparam \dio_rdata_l_2x[24]~24 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_l_2x[24]~24 .shared_arith = "off";

arriaii_lcell_comb \rdata_n_ams[25]~25 (
	.dataa(!\dqs_group[3].dq_dqs|wire_bidir_dq_1_ddio_in_inst_regouthi ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_n_ams[25]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_n_ams[25]~25 .extended_lut = "off";
defparam \rdata_n_ams[25]~25 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_n_ams[25]~25 .shared_arith = "off";

dffeas \rdata_n_ams[25] (
	.clk(resync_clk_2x),
	.d(\rdata_n_ams[25]~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[25]~q ),
	.prn(vcc));
defparam \rdata_n_ams[25] .is_wysiwyg = "true";
defparam \rdata_n_ams[25] .power_up = "low";

arriaii_lcell_comb \dio_rdata_l_2x[25]~25 (
	.dataa(!\rdata_n_ams[25]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_l_2x[25]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_l_2x[25]~25 .extended_lut = "off";
defparam \dio_rdata_l_2x[25]~25 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_l_2x[25]~25 .shared_arith = "off";

arriaii_lcell_comb \rdata_n_ams[26]~26 (
	.dataa(!\dqs_group[3].dq_dqs|wire_bidir_dq_2_ddio_in_inst_regouthi ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_n_ams[26]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_n_ams[26]~26 .extended_lut = "off";
defparam \rdata_n_ams[26]~26 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_n_ams[26]~26 .shared_arith = "off";

dffeas \rdata_n_ams[26] (
	.clk(resync_clk_2x),
	.d(\rdata_n_ams[26]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[26]~q ),
	.prn(vcc));
defparam \rdata_n_ams[26] .is_wysiwyg = "true";
defparam \rdata_n_ams[26] .power_up = "low";

arriaii_lcell_comb \dio_rdata_l_2x[26]~26 (
	.dataa(!\rdata_n_ams[26]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_l_2x[26]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_l_2x[26]~26 .extended_lut = "off";
defparam \dio_rdata_l_2x[26]~26 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_l_2x[26]~26 .shared_arith = "off";

arriaii_lcell_comb \rdata_n_ams[27]~27 (
	.dataa(!\dqs_group[3].dq_dqs|wire_bidir_dq_3_ddio_in_inst_regouthi ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_n_ams[27]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_n_ams[27]~27 .extended_lut = "off";
defparam \rdata_n_ams[27]~27 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_n_ams[27]~27 .shared_arith = "off";

dffeas \rdata_n_ams[27] (
	.clk(resync_clk_2x),
	.d(\rdata_n_ams[27]~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[27]~q ),
	.prn(vcc));
defparam \rdata_n_ams[27] .is_wysiwyg = "true";
defparam \rdata_n_ams[27] .power_up = "low";

arriaii_lcell_comb \dio_rdata_l_2x[27]~27 (
	.dataa(!\rdata_n_ams[27]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_l_2x[27]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_l_2x[27]~27 .extended_lut = "off";
defparam \dio_rdata_l_2x[27]~27 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_l_2x[27]~27 .shared_arith = "off";

arriaii_lcell_comb \rdata_n_ams[28]~28 (
	.dataa(!\dqs_group[3].dq_dqs|wire_bidir_dq_4_ddio_in_inst_regouthi ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_n_ams[28]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_n_ams[28]~28 .extended_lut = "off";
defparam \rdata_n_ams[28]~28 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_n_ams[28]~28 .shared_arith = "off";

dffeas \rdata_n_ams[28] (
	.clk(resync_clk_2x),
	.d(\rdata_n_ams[28]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[28]~q ),
	.prn(vcc));
defparam \rdata_n_ams[28] .is_wysiwyg = "true";
defparam \rdata_n_ams[28] .power_up = "low";

arriaii_lcell_comb \dio_rdata_l_2x[28]~28 (
	.dataa(!\rdata_n_ams[28]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_l_2x[28]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_l_2x[28]~28 .extended_lut = "off";
defparam \dio_rdata_l_2x[28]~28 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_l_2x[28]~28 .shared_arith = "off";

arriaii_lcell_comb \rdata_n_ams[29]~29 (
	.dataa(!\dqs_group[3].dq_dqs|wire_bidir_dq_5_ddio_in_inst_regouthi ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_n_ams[29]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_n_ams[29]~29 .extended_lut = "off";
defparam \rdata_n_ams[29]~29 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_n_ams[29]~29 .shared_arith = "off";

dffeas \rdata_n_ams[29] (
	.clk(resync_clk_2x),
	.d(\rdata_n_ams[29]~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[29]~q ),
	.prn(vcc));
defparam \rdata_n_ams[29] .is_wysiwyg = "true";
defparam \rdata_n_ams[29] .power_up = "low";

arriaii_lcell_comb \dio_rdata_l_2x[29]~29 (
	.dataa(!\rdata_n_ams[29]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_l_2x[29]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_l_2x[29]~29 .extended_lut = "off";
defparam \dio_rdata_l_2x[29]~29 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_l_2x[29]~29 .shared_arith = "off";

arriaii_lcell_comb \rdata_n_ams[30]~30 (
	.dataa(!\dqs_group[3].dq_dqs|wire_bidir_dq_6_ddio_in_inst_regouthi ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_n_ams[30]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_n_ams[30]~30 .extended_lut = "off";
defparam \rdata_n_ams[30]~30 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_n_ams[30]~30 .shared_arith = "off";

dffeas \rdata_n_ams[30] (
	.clk(resync_clk_2x),
	.d(\rdata_n_ams[30]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[30]~q ),
	.prn(vcc));
defparam \rdata_n_ams[30] .is_wysiwyg = "true";
defparam \rdata_n_ams[30] .power_up = "low";

arriaii_lcell_comb \dio_rdata_l_2x[30]~30 (
	.dataa(!\rdata_n_ams[30]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_l_2x[30]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_l_2x[30]~30 .extended_lut = "off";
defparam \dio_rdata_l_2x[30]~30 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_l_2x[30]~30 .shared_arith = "off";

arriaii_lcell_comb \rdata_n_ams[31]~31 (
	.dataa(!\dqs_group[3].dq_dqs|wire_bidir_dq_7_ddio_in_inst_regouthi ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rdata_n_ams[31]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rdata_n_ams[31]~31 .extended_lut = "off";
defparam \rdata_n_ams[31]~31 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rdata_n_ams[31]~31 .shared_arith = "off";

dffeas \rdata_n_ams[31] (
	.clk(resync_clk_2x),
	.d(\rdata_n_ams[31]~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rdata_n_ams[31]~q ),
	.prn(vcc));
defparam \rdata_n_ams[31] .is_wysiwyg = "true";
defparam \rdata_n_ams[31] .power_up = "low";

arriaii_lcell_comb \dio_rdata_l_2x[31]~31 (
	.dataa(!\rdata_n_ams[31]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dio_rdata_l_2x[31]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dio_rdata_l_2x[31]~31 .extended_lut = "off";
defparam \dio_rdata_l_2x[31]~31 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dio_rdata_l_2x[31]~31 .shared_arith = "off";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_dq_dqs (
	dqs_output_reg_clk,
	dq_output_reg_clk,
	dqs_enable_ctrl_clk,
	dll_delayctrlin,
	output_dq_output_data_out,
	output_dq_output_data_in_low,
	output_dq_output_data_in_high,
	bidir_dq_output_data_out,
	bidir_dq_input_data_out_low,
	bidir_dq_input_data_out_high,
	bidir_dq_output_data_in_low,
	bidir_dq_output_data_in_high,
	dq_oe_2x_0,
	dq_oe_2x_1,
	dqs_output_data_out,
	bidir_dq_input_data_in,
	dqs_input_data_in,
	bidir_dq_0_oe_ff_inst1,
	bidir_dq_1_oe_ff_inst1,
	bidir_dq_2_oe_ff_inst1,
	bidir_dq_3_oe_ff_inst1,
	bidir_dq_4_oe_ff_inst1,
	bidir_dq_5_oe_ff_inst1,
	bidir_dq_6_oe_ff_inst1,
	bidir_dq_7_oe_ff_inst1,
	dqs_0_oe_ff_inst1,
	dqsn_0_oe_ff_inst1,
	bidir_dq_areset,
	dqs_output_data_in_high,
	dqs_enable_ctrl_in)/* synthesis synthesis_greybox=0 */;
input 	dqs_output_reg_clk;
input 	dq_output_reg_clk;
input 	dqs_enable_ctrl_clk;
input 	[5:0] dll_delayctrlin;
output 	[0:0] output_dq_output_data_out;
input 	[0:0] output_dq_output_data_in_low;
input 	[0:0] output_dq_output_data_in_high;
output 	[7:0] bidir_dq_output_data_out;
output 	[7:0] bidir_dq_input_data_out_low;
output 	[7:0] bidir_dq_input_data_out_high;
input 	[7:0] bidir_dq_output_data_in_low;
input 	[7:0] bidir_dq_output_data_in_high;
input 	dq_oe_2x_0;
input 	dq_oe_2x_1;
output 	[0:0] dqs_output_data_out;
input 	[7:0] bidir_dq_input_data_in;
input 	[0:0] dqs_input_data_in;
output 	bidir_dq_0_oe_ff_inst1;
output 	bidir_dq_1_oe_ff_inst1;
output 	bidir_dq_2_oe_ff_inst1;
output 	bidir_dq_3_oe_ff_inst1;
output 	bidir_dq_4_oe_ff_inst1;
output 	bidir_dq_5_oe_ff_inst1;
output 	bidir_dq_6_oe_ff_inst1;
output 	bidir_dq_7_oe_ff_inst1;
output 	dqs_0_oe_ff_inst1;
output 	dqsn_0_oe_ff_inst1;
input 	[7:0] bidir_dq_areset;
input 	[0:0] dqs_output_data_in_high;
input 	dqs_enable_ctrl_in;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire wire_dqs_0_delay_chain_inst_dqsbusout;
wire wire_dqs_0_enable_ctrl_inst_dqsenableout;
wire wire_dqs_0_enable_inst_dqsbusout;
wire \bidir_dq_0_oe_ff_inst~0_combout ;
wire \bidir_dq_1_oe_ff_inst~0_combout ;
wire \bidir_dq_2_oe_ff_inst~0_combout ;
wire \bidir_dq_3_oe_ff_inst~0_combout ;
wire \bidir_dq_4_oe_ff_inst~0_combout ;
wire \bidir_dq_5_oe_ff_inst~0_combout ;
wire \bidir_dq_6_oe_ff_inst~0_combout ;
wire \bidir_dq_7_oe_ff_inst~0_combout ;
wire \dqs_0_oe_ff_inst~0_combout ;
wire \dqsn_0_oe_ff_inst~0_combout ;


arriaii_ddio_out output_dq_0_output_ddio_out_inst(
	.datainlo(output_dq_output_data_in_low[0]),
	.datainhi(output_dq_output_data_in_high[0]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.clk(gnd),
	.dataout(output_dq_output_data_out[0]),
	.dfflo(),
	.dffhi());
defparam output_dq_0_output_ddio_out_inst.async_mode = "clear";
defparam output_dq_0_output_ddio_out_inst.power_up = "low";
defparam output_dq_0_output_ddio_out_inst.sync_mode = "none";
defparam output_dq_0_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_out bidir_dq_0_output_ddio_out_inst(
	.datainlo(bidir_dq_output_data_in_low[0]),
	.datainhi(bidir_dq_output_data_in_high[0]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(!bidir_dq_areset[1]),
	.sreset(gnd),
	.clk(gnd),
	.dataout(bidir_dq_output_data_out[0]),
	.dfflo(),
	.dffhi());
defparam bidir_dq_0_output_ddio_out_inst.async_mode = "clear";
defparam bidir_dq_0_output_ddio_out_inst.power_up = "low";
defparam bidir_dq_0_output_ddio_out_inst.sync_mode = "none";
defparam bidir_dq_0_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_out bidir_dq_1_output_ddio_out_inst(
	.datainlo(bidir_dq_output_data_in_low[1]),
	.datainhi(bidir_dq_output_data_in_high[1]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(!bidir_dq_areset[1]),
	.sreset(gnd),
	.clk(gnd),
	.dataout(bidir_dq_output_data_out[1]),
	.dfflo(),
	.dffhi());
defparam bidir_dq_1_output_ddio_out_inst.async_mode = "clear";
defparam bidir_dq_1_output_ddio_out_inst.power_up = "low";
defparam bidir_dq_1_output_ddio_out_inst.sync_mode = "none";
defparam bidir_dq_1_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_out bidir_dq_2_output_ddio_out_inst(
	.datainlo(bidir_dq_output_data_in_low[2]),
	.datainhi(bidir_dq_output_data_in_high[2]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(!bidir_dq_areset[1]),
	.sreset(gnd),
	.clk(gnd),
	.dataout(bidir_dq_output_data_out[2]),
	.dfflo(),
	.dffhi());
defparam bidir_dq_2_output_ddio_out_inst.async_mode = "clear";
defparam bidir_dq_2_output_ddio_out_inst.power_up = "low";
defparam bidir_dq_2_output_ddio_out_inst.sync_mode = "none";
defparam bidir_dq_2_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_out bidir_dq_3_output_ddio_out_inst(
	.datainlo(bidir_dq_output_data_in_low[3]),
	.datainhi(bidir_dq_output_data_in_high[3]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(!bidir_dq_areset[1]),
	.sreset(gnd),
	.clk(gnd),
	.dataout(bidir_dq_output_data_out[3]),
	.dfflo(),
	.dffhi());
defparam bidir_dq_3_output_ddio_out_inst.async_mode = "clear";
defparam bidir_dq_3_output_ddio_out_inst.power_up = "low";
defparam bidir_dq_3_output_ddio_out_inst.sync_mode = "none";
defparam bidir_dq_3_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_out bidir_dq_4_output_ddio_out_inst(
	.datainlo(bidir_dq_output_data_in_low[4]),
	.datainhi(bidir_dq_output_data_in_high[4]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(!bidir_dq_areset[1]),
	.sreset(gnd),
	.clk(gnd),
	.dataout(bidir_dq_output_data_out[4]),
	.dfflo(),
	.dffhi());
defparam bidir_dq_4_output_ddio_out_inst.async_mode = "clear";
defparam bidir_dq_4_output_ddio_out_inst.power_up = "low";
defparam bidir_dq_4_output_ddio_out_inst.sync_mode = "none";
defparam bidir_dq_4_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_out bidir_dq_5_output_ddio_out_inst(
	.datainlo(bidir_dq_output_data_in_low[5]),
	.datainhi(bidir_dq_output_data_in_high[5]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(!bidir_dq_areset[1]),
	.sreset(gnd),
	.clk(gnd),
	.dataout(bidir_dq_output_data_out[5]),
	.dfflo(),
	.dffhi());
defparam bidir_dq_5_output_ddio_out_inst.async_mode = "clear";
defparam bidir_dq_5_output_ddio_out_inst.power_up = "low";
defparam bidir_dq_5_output_ddio_out_inst.sync_mode = "none";
defparam bidir_dq_5_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_out bidir_dq_6_output_ddio_out_inst(
	.datainlo(bidir_dq_output_data_in_low[6]),
	.datainhi(bidir_dq_output_data_in_high[6]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(!bidir_dq_areset[1]),
	.sreset(gnd),
	.clk(gnd),
	.dataout(bidir_dq_output_data_out[6]),
	.dfflo(),
	.dffhi());
defparam bidir_dq_6_output_ddio_out_inst.async_mode = "clear";
defparam bidir_dq_6_output_ddio_out_inst.power_up = "low";
defparam bidir_dq_6_output_ddio_out_inst.sync_mode = "none";
defparam bidir_dq_6_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_out bidir_dq_7_output_ddio_out_inst(
	.datainlo(bidir_dq_output_data_in_low[7]),
	.datainhi(bidir_dq_output_data_in_high[7]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(!bidir_dq_areset[1]),
	.sreset(gnd),
	.clk(gnd),
	.dataout(bidir_dq_output_data_out[7]),
	.dfflo(),
	.dffhi());
defparam bidir_dq_7_output_ddio_out_inst.async_mode = "clear";
defparam bidir_dq_7_output_ddio_out_inst.power_up = "low";
defparam bidir_dq_7_output_ddio_out_inst.sync_mode = "none";
defparam bidir_dq_7_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_in bidir_dq_0_ddio_in_inst(
	.datain(bidir_dq_input_data_in[0]),
	.clk(!wire_dqs_0_enable_inst_dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(bidir_dq_input_data_out_low[0]),
	.regouthi(bidir_dq_input_data_out_high[0]),
	.dfflo());
defparam bidir_dq_0_ddio_in_inst.async_mode = "none";
defparam bidir_dq_0_ddio_in_inst.power_up = "low";
defparam bidir_dq_0_ddio_in_inst.sync_mode = "none";
defparam bidir_dq_0_ddio_in_inst.use_clkn = "false";

arriaii_ddio_in bidir_dq_1_ddio_in_inst(
	.datain(bidir_dq_input_data_in[1]),
	.clk(!wire_dqs_0_enable_inst_dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(bidir_dq_input_data_out_low[1]),
	.regouthi(bidir_dq_input_data_out_high[1]),
	.dfflo());
defparam bidir_dq_1_ddio_in_inst.async_mode = "none";
defparam bidir_dq_1_ddio_in_inst.power_up = "low";
defparam bidir_dq_1_ddio_in_inst.sync_mode = "none";
defparam bidir_dq_1_ddio_in_inst.use_clkn = "false";

arriaii_ddio_in bidir_dq_2_ddio_in_inst(
	.datain(bidir_dq_input_data_in[2]),
	.clk(!wire_dqs_0_enable_inst_dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(bidir_dq_input_data_out_low[2]),
	.regouthi(bidir_dq_input_data_out_high[2]),
	.dfflo());
defparam bidir_dq_2_ddio_in_inst.async_mode = "none";
defparam bidir_dq_2_ddio_in_inst.power_up = "low";
defparam bidir_dq_2_ddio_in_inst.sync_mode = "none";
defparam bidir_dq_2_ddio_in_inst.use_clkn = "false";

arriaii_ddio_in bidir_dq_3_ddio_in_inst(
	.datain(bidir_dq_input_data_in[3]),
	.clk(!wire_dqs_0_enable_inst_dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(bidir_dq_input_data_out_low[3]),
	.regouthi(bidir_dq_input_data_out_high[3]),
	.dfflo());
defparam bidir_dq_3_ddio_in_inst.async_mode = "none";
defparam bidir_dq_3_ddio_in_inst.power_up = "low";
defparam bidir_dq_3_ddio_in_inst.sync_mode = "none";
defparam bidir_dq_3_ddio_in_inst.use_clkn = "false";

arriaii_ddio_in bidir_dq_4_ddio_in_inst(
	.datain(bidir_dq_input_data_in[4]),
	.clk(!wire_dqs_0_enable_inst_dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(bidir_dq_input_data_out_low[4]),
	.regouthi(bidir_dq_input_data_out_high[4]),
	.dfflo());
defparam bidir_dq_4_ddio_in_inst.async_mode = "none";
defparam bidir_dq_4_ddio_in_inst.power_up = "low";
defparam bidir_dq_4_ddio_in_inst.sync_mode = "none";
defparam bidir_dq_4_ddio_in_inst.use_clkn = "false";

arriaii_ddio_in bidir_dq_5_ddio_in_inst(
	.datain(bidir_dq_input_data_in[5]),
	.clk(!wire_dqs_0_enable_inst_dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(bidir_dq_input_data_out_low[5]),
	.regouthi(bidir_dq_input_data_out_high[5]),
	.dfflo());
defparam bidir_dq_5_ddio_in_inst.async_mode = "none";
defparam bidir_dq_5_ddio_in_inst.power_up = "low";
defparam bidir_dq_5_ddio_in_inst.sync_mode = "none";
defparam bidir_dq_5_ddio_in_inst.use_clkn = "false";

arriaii_ddio_in bidir_dq_6_ddio_in_inst(
	.datain(bidir_dq_input_data_in[6]),
	.clk(!wire_dqs_0_enable_inst_dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(bidir_dq_input_data_out_low[6]),
	.regouthi(bidir_dq_input_data_out_high[6]),
	.dfflo());
defparam bidir_dq_6_ddio_in_inst.async_mode = "none";
defparam bidir_dq_6_ddio_in_inst.power_up = "low";
defparam bidir_dq_6_ddio_in_inst.sync_mode = "none";
defparam bidir_dq_6_ddio_in_inst.use_clkn = "false";

arriaii_ddio_in bidir_dq_7_ddio_in_inst(
	.datain(bidir_dq_input_data_in[7]),
	.clk(!wire_dqs_0_enable_inst_dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(bidir_dq_input_data_out_low[7]),
	.regouthi(bidir_dq_input_data_out_high[7]),
	.dfflo());
defparam bidir_dq_7_ddio_in_inst.async_mode = "none";
defparam bidir_dq_7_ddio_in_inst.power_up = "low";
defparam bidir_dq_7_ddio_in_inst.sync_mode = "none";
defparam bidir_dq_7_ddio_in_inst.use_clkn = "false";

arriaii_ddio_out dqs_0_output_ddio_out_inst(
	.datainlo(gnd),
	.datainhi(dqs_output_data_in_high[0]),
	.clkhi(dqs_output_reg_clk),
	.clklo(dqs_output_reg_clk),
	.muxsel(dqs_output_reg_clk),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.clk(gnd),
	.dataout(dqs_output_data_out[0]),
	.dfflo(),
	.dffhi());
defparam dqs_0_output_ddio_out_inst.async_mode = "none";
defparam dqs_0_output_ddio_out_inst.power_up = "low";
defparam dqs_0_output_ddio_out_inst.sync_mode = "none";
defparam dqs_0_output_ddio_out_inst.use_new_clocking_model = "true";

dffeas bidir_dq_0_oe_ff_inst(
	.clk(dq_output_reg_clk),
	.d(\bidir_dq_0_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(bidir_dq_0_oe_ff_inst1),
	.prn(vcc));
defparam bidir_dq_0_oe_ff_inst.is_wysiwyg = "true";
defparam bidir_dq_0_oe_ff_inst.power_up = "low";

dffeas bidir_dq_1_oe_ff_inst(
	.clk(dq_output_reg_clk),
	.d(\bidir_dq_1_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(bidir_dq_1_oe_ff_inst1),
	.prn(vcc));
defparam bidir_dq_1_oe_ff_inst.is_wysiwyg = "true";
defparam bidir_dq_1_oe_ff_inst.power_up = "low";

dffeas bidir_dq_2_oe_ff_inst(
	.clk(dq_output_reg_clk),
	.d(\bidir_dq_2_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(bidir_dq_2_oe_ff_inst1),
	.prn(vcc));
defparam bidir_dq_2_oe_ff_inst.is_wysiwyg = "true";
defparam bidir_dq_2_oe_ff_inst.power_up = "low";

dffeas bidir_dq_3_oe_ff_inst(
	.clk(dq_output_reg_clk),
	.d(\bidir_dq_3_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(bidir_dq_3_oe_ff_inst1),
	.prn(vcc));
defparam bidir_dq_3_oe_ff_inst.is_wysiwyg = "true";
defparam bidir_dq_3_oe_ff_inst.power_up = "low";

dffeas bidir_dq_4_oe_ff_inst(
	.clk(dq_output_reg_clk),
	.d(\bidir_dq_4_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(bidir_dq_4_oe_ff_inst1),
	.prn(vcc));
defparam bidir_dq_4_oe_ff_inst.is_wysiwyg = "true";
defparam bidir_dq_4_oe_ff_inst.power_up = "low";

dffeas bidir_dq_5_oe_ff_inst(
	.clk(dq_output_reg_clk),
	.d(\bidir_dq_5_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(bidir_dq_5_oe_ff_inst1),
	.prn(vcc));
defparam bidir_dq_5_oe_ff_inst.is_wysiwyg = "true";
defparam bidir_dq_5_oe_ff_inst.power_up = "low";

dffeas bidir_dq_6_oe_ff_inst(
	.clk(dq_output_reg_clk),
	.d(\bidir_dq_6_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(bidir_dq_6_oe_ff_inst1),
	.prn(vcc));
defparam bidir_dq_6_oe_ff_inst.is_wysiwyg = "true";
defparam bidir_dq_6_oe_ff_inst.power_up = "low";

dffeas bidir_dq_7_oe_ff_inst(
	.clk(dq_output_reg_clk),
	.d(\bidir_dq_7_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(bidir_dq_7_oe_ff_inst1),
	.prn(vcc));
defparam bidir_dq_7_oe_ff_inst.is_wysiwyg = "true";
defparam bidir_dq_7_oe_ff_inst.power_up = "low";

dffeas dqs_0_oe_ff_inst(
	.clk(dqs_output_reg_clk),
	.d(\dqs_0_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dqs_0_oe_ff_inst1),
	.prn(vcc));
defparam dqs_0_oe_ff_inst.is_wysiwyg = "true";
defparam dqs_0_oe_ff_inst.power_up = "low";

dffeas dqsn_0_oe_ff_inst(
	.clk(dqs_output_reg_clk),
	.d(\dqsn_0_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dqsn_0_oe_ff_inst1),
	.prn(vcc));
defparam dqsn_0_oe_ff_inst.is_wysiwyg = "true";
defparam dqsn_0_oe_ff_inst.power_up = "low";

arriaii_dqs_delay_chain dqs_0_delay_chain_inst(
	.dqsin(dqs_input_data_in[0]),
	.dqsupdateen(gnd),
	.delayctrlin({dll_delayctrlin[5],dll_delayctrlin[4],dll_delayctrlin[3],dll_delayctrlin[2],dll_delayctrlin[1],dll_delayctrlin[0]}),
	.offsetctrlin(6'b000000),
	.dqsbusout(wire_dqs_0_delay_chain_inst_dqsbusout));
defparam dqs_0_delay_chain_inst.delay_buffer_mode = "high";
defparam dqs_0_delay_chain_inst.dqs_ctrl_latches_enable = "false";
defparam dqs_0_delay_chain_inst.dqs_input_frequency = "3333ps";
defparam dqs_0_delay_chain_inst.dqs_offsetctrl_enable = "false";
defparam dqs_0_delay_chain_inst.dqs_phase_shift = 7200;
defparam dqs_0_delay_chain_inst.phase_setting = 2;
defparam dqs_0_delay_chain_inst.sim_buffer_delay_increment = 10;
defparam dqs_0_delay_chain_inst.sim_high_buffer_intrinsic_delay = 175;
defparam dqs_0_delay_chain_inst.sim_low_buffer_intrinsic_delay = 350;
defparam dqs_0_delay_chain_inst.test_enable = "false";
defparam dqs_0_delay_chain_inst.test_select = 0;

arriaii_dqs_enable_ctrl dqs_0_enable_ctrl_inst(
	.dqsenablein(dqs_enable_ctrl_in),
	.clk(dqs_enable_ctrl_clk),
	.dqsenableout(wire_dqs_0_enable_ctrl_inst_dqsenableout));
defparam dqs_0_enable_ctrl_inst.delay_dqs_enable_by_half_cycle = "true";

arriaii_dqs_enable dqs_0_enable_inst(
	.dqsin(wire_dqs_0_delay_chain_inst_dqsbusout),
	.dqsenable(wire_dqs_0_enable_ctrl_inst_dqsenableout),
	.dqsbusout(wire_dqs_0_enable_inst_dqsbusout));

arriaii_lcell_comb \bidir_dq_0_oe_ff_inst~0 (
	.dataa(!dq_oe_2x_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bidir_dq_0_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bidir_dq_0_oe_ff_inst~0 .extended_lut = "off";
defparam \bidir_dq_0_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \bidir_dq_0_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \bidir_dq_1_oe_ff_inst~0 (
	.dataa(!dq_oe_2x_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bidir_dq_1_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bidir_dq_1_oe_ff_inst~0 .extended_lut = "off";
defparam \bidir_dq_1_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \bidir_dq_1_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \bidir_dq_2_oe_ff_inst~0 (
	.dataa(!dq_oe_2x_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bidir_dq_2_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bidir_dq_2_oe_ff_inst~0 .extended_lut = "off";
defparam \bidir_dq_2_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \bidir_dq_2_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \bidir_dq_3_oe_ff_inst~0 (
	.dataa(!dq_oe_2x_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bidir_dq_3_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bidir_dq_3_oe_ff_inst~0 .extended_lut = "off";
defparam \bidir_dq_3_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \bidir_dq_3_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \bidir_dq_4_oe_ff_inst~0 (
	.dataa(!dq_oe_2x_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bidir_dq_4_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bidir_dq_4_oe_ff_inst~0 .extended_lut = "off";
defparam \bidir_dq_4_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \bidir_dq_4_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \bidir_dq_5_oe_ff_inst~0 (
	.dataa(!dq_oe_2x_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bidir_dq_5_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bidir_dq_5_oe_ff_inst~0 .extended_lut = "off";
defparam \bidir_dq_5_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \bidir_dq_5_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \bidir_dq_6_oe_ff_inst~0 (
	.dataa(!dq_oe_2x_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bidir_dq_6_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bidir_dq_6_oe_ff_inst~0 .extended_lut = "off";
defparam \bidir_dq_6_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \bidir_dq_6_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \bidir_dq_7_oe_ff_inst~0 (
	.dataa(!dq_oe_2x_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bidir_dq_7_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bidir_dq_7_oe_ff_inst~0 .extended_lut = "off";
defparam \bidir_dq_7_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \bidir_dq_7_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \dqs_0_oe_ff_inst~0 (
	.dataa(!dqs_output_data_in_high[0]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dqs_0_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dqs_0_oe_ff_inst~0 .extended_lut = "off";
defparam \dqs_0_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dqs_0_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \dqsn_0_oe_ff_inst~0 (
	.dataa(!dqs_output_data_in_high[0]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dqsn_0_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dqsn_0_oe_ff_inst~0 .extended_lut = "off";
defparam \dqsn_0_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dqsn_0_oe_ff_inst~0 .shared_arith = "off";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_dq_dqs_1 (
	dqs_output_reg_clk,
	dq_output_reg_clk,
	dqs_enable_ctrl_clk,
	dll_delayctrlin,
	output_dq_output_data_out,
	output_dq_output_data_in_low,
	output_dq_output_data_in_high,
	bidir_dq_output_data_out,
	bidir_dq_input_data_out_low,
	bidir_dq_input_data_out_high,
	bidir_dq_output_data_in_low,
	bidir_dq_output_data_in_high,
	dq_oe_2x_2,
	dq_oe_2x_3,
	dqs_output_data_out,
	bidir_dq_input_data_in,
	dqs_input_data_in,
	bidir_dq_0_oe_ff_inst1,
	bidir_dq_1_oe_ff_inst1,
	bidir_dq_2_oe_ff_inst1,
	bidir_dq_3_oe_ff_inst1,
	bidir_dq_4_oe_ff_inst1,
	bidir_dq_5_oe_ff_inst1,
	bidir_dq_6_oe_ff_inst1,
	bidir_dq_7_oe_ff_inst1,
	dqs_0_oe_ff_inst1,
	dqsn_0_oe_ff_inst1,
	bidir_dq_areset,
	dqs_output_data_in_high,
	dqs_enable_ctrl_in)/* synthesis synthesis_greybox=0 */;
input 	dqs_output_reg_clk;
input 	dq_output_reg_clk;
input 	dqs_enable_ctrl_clk;
input 	[5:0] dll_delayctrlin;
output 	[0:0] output_dq_output_data_out;
input 	[0:0] output_dq_output_data_in_low;
input 	[0:0] output_dq_output_data_in_high;
output 	[7:0] bidir_dq_output_data_out;
output 	[7:0] bidir_dq_input_data_out_low;
output 	[7:0] bidir_dq_input_data_out_high;
input 	[7:0] bidir_dq_output_data_in_low;
input 	[7:0] bidir_dq_output_data_in_high;
input 	dq_oe_2x_2;
input 	dq_oe_2x_3;
output 	[0:0] dqs_output_data_out;
input 	[7:0] bidir_dq_input_data_in;
input 	[0:0] dqs_input_data_in;
output 	bidir_dq_0_oe_ff_inst1;
output 	bidir_dq_1_oe_ff_inst1;
output 	bidir_dq_2_oe_ff_inst1;
output 	bidir_dq_3_oe_ff_inst1;
output 	bidir_dq_4_oe_ff_inst1;
output 	bidir_dq_5_oe_ff_inst1;
output 	bidir_dq_6_oe_ff_inst1;
output 	bidir_dq_7_oe_ff_inst1;
output 	dqs_0_oe_ff_inst1;
output 	dqsn_0_oe_ff_inst1;
input 	[7:0] bidir_dq_areset;
input 	[0:0] dqs_output_data_in_high;
input 	dqs_enable_ctrl_in;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire wire_dqs_0_delay_chain_inst_dqsbusout;
wire wire_dqs_0_enable_ctrl_inst_dqsenableout;
wire wire_dqs_0_enable_inst_dqsbusout;
wire \bidir_dq_0_oe_ff_inst~0_combout ;
wire \bidir_dq_1_oe_ff_inst~0_combout ;
wire \bidir_dq_2_oe_ff_inst~0_combout ;
wire \bidir_dq_3_oe_ff_inst~0_combout ;
wire \bidir_dq_4_oe_ff_inst~0_combout ;
wire \bidir_dq_5_oe_ff_inst~0_combout ;
wire \bidir_dq_6_oe_ff_inst~0_combout ;
wire \bidir_dq_7_oe_ff_inst~0_combout ;
wire \dqs_0_oe_ff_inst~0_combout ;
wire \dqsn_0_oe_ff_inst~0_combout ;


arriaii_ddio_out output_dq_0_output_ddio_out_inst(
	.datainlo(output_dq_output_data_in_low[0]),
	.datainhi(output_dq_output_data_in_high[0]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.clk(gnd),
	.dataout(output_dq_output_data_out[0]),
	.dfflo(),
	.dffhi());
defparam output_dq_0_output_ddio_out_inst.async_mode = "clear";
defparam output_dq_0_output_ddio_out_inst.power_up = "low";
defparam output_dq_0_output_ddio_out_inst.sync_mode = "none";
defparam output_dq_0_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_out bidir_dq_0_output_ddio_out_inst(
	.datainlo(bidir_dq_output_data_in_low[0]),
	.datainhi(bidir_dq_output_data_in_high[0]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(!bidir_dq_areset[1]),
	.sreset(gnd),
	.clk(gnd),
	.dataout(bidir_dq_output_data_out[0]),
	.dfflo(),
	.dffhi());
defparam bidir_dq_0_output_ddio_out_inst.async_mode = "clear";
defparam bidir_dq_0_output_ddio_out_inst.power_up = "low";
defparam bidir_dq_0_output_ddio_out_inst.sync_mode = "none";
defparam bidir_dq_0_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_out bidir_dq_1_output_ddio_out_inst(
	.datainlo(bidir_dq_output_data_in_low[1]),
	.datainhi(bidir_dq_output_data_in_high[1]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(!bidir_dq_areset[1]),
	.sreset(gnd),
	.clk(gnd),
	.dataout(bidir_dq_output_data_out[1]),
	.dfflo(),
	.dffhi());
defparam bidir_dq_1_output_ddio_out_inst.async_mode = "clear";
defparam bidir_dq_1_output_ddio_out_inst.power_up = "low";
defparam bidir_dq_1_output_ddio_out_inst.sync_mode = "none";
defparam bidir_dq_1_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_out bidir_dq_2_output_ddio_out_inst(
	.datainlo(bidir_dq_output_data_in_low[2]),
	.datainhi(bidir_dq_output_data_in_high[2]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(!bidir_dq_areset[1]),
	.sreset(gnd),
	.clk(gnd),
	.dataout(bidir_dq_output_data_out[2]),
	.dfflo(),
	.dffhi());
defparam bidir_dq_2_output_ddio_out_inst.async_mode = "clear";
defparam bidir_dq_2_output_ddio_out_inst.power_up = "low";
defparam bidir_dq_2_output_ddio_out_inst.sync_mode = "none";
defparam bidir_dq_2_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_out bidir_dq_3_output_ddio_out_inst(
	.datainlo(bidir_dq_output_data_in_low[3]),
	.datainhi(bidir_dq_output_data_in_high[3]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(!bidir_dq_areset[1]),
	.sreset(gnd),
	.clk(gnd),
	.dataout(bidir_dq_output_data_out[3]),
	.dfflo(),
	.dffhi());
defparam bidir_dq_3_output_ddio_out_inst.async_mode = "clear";
defparam bidir_dq_3_output_ddio_out_inst.power_up = "low";
defparam bidir_dq_3_output_ddio_out_inst.sync_mode = "none";
defparam bidir_dq_3_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_out bidir_dq_4_output_ddio_out_inst(
	.datainlo(bidir_dq_output_data_in_low[4]),
	.datainhi(bidir_dq_output_data_in_high[4]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(!bidir_dq_areset[1]),
	.sreset(gnd),
	.clk(gnd),
	.dataout(bidir_dq_output_data_out[4]),
	.dfflo(),
	.dffhi());
defparam bidir_dq_4_output_ddio_out_inst.async_mode = "clear";
defparam bidir_dq_4_output_ddio_out_inst.power_up = "low";
defparam bidir_dq_4_output_ddio_out_inst.sync_mode = "none";
defparam bidir_dq_4_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_out bidir_dq_5_output_ddio_out_inst(
	.datainlo(bidir_dq_output_data_in_low[5]),
	.datainhi(bidir_dq_output_data_in_high[5]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(!bidir_dq_areset[1]),
	.sreset(gnd),
	.clk(gnd),
	.dataout(bidir_dq_output_data_out[5]),
	.dfflo(),
	.dffhi());
defparam bidir_dq_5_output_ddio_out_inst.async_mode = "clear";
defparam bidir_dq_5_output_ddio_out_inst.power_up = "low";
defparam bidir_dq_5_output_ddio_out_inst.sync_mode = "none";
defparam bidir_dq_5_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_out bidir_dq_6_output_ddio_out_inst(
	.datainlo(bidir_dq_output_data_in_low[6]),
	.datainhi(bidir_dq_output_data_in_high[6]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(!bidir_dq_areset[1]),
	.sreset(gnd),
	.clk(gnd),
	.dataout(bidir_dq_output_data_out[6]),
	.dfflo(),
	.dffhi());
defparam bidir_dq_6_output_ddio_out_inst.async_mode = "clear";
defparam bidir_dq_6_output_ddio_out_inst.power_up = "low";
defparam bidir_dq_6_output_ddio_out_inst.sync_mode = "none";
defparam bidir_dq_6_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_out bidir_dq_7_output_ddio_out_inst(
	.datainlo(bidir_dq_output_data_in_low[7]),
	.datainhi(bidir_dq_output_data_in_high[7]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(!bidir_dq_areset[1]),
	.sreset(gnd),
	.clk(gnd),
	.dataout(bidir_dq_output_data_out[7]),
	.dfflo(),
	.dffhi());
defparam bidir_dq_7_output_ddio_out_inst.async_mode = "clear";
defparam bidir_dq_7_output_ddio_out_inst.power_up = "low";
defparam bidir_dq_7_output_ddio_out_inst.sync_mode = "none";
defparam bidir_dq_7_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_in bidir_dq_0_ddio_in_inst(
	.datain(bidir_dq_input_data_in[0]),
	.clk(!wire_dqs_0_enable_inst_dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(bidir_dq_input_data_out_low[0]),
	.regouthi(bidir_dq_input_data_out_high[0]),
	.dfflo());
defparam bidir_dq_0_ddio_in_inst.async_mode = "none";
defparam bidir_dq_0_ddio_in_inst.power_up = "low";
defparam bidir_dq_0_ddio_in_inst.sync_mode = "none";
defparam bidir_dq_0_ddio_in_inst.use_clkn = "false";

arriaii_ddio_in bidir_dq_1_ddio_in_inst(
	.datain(bidir_dq_input_data_in[1]),
	.clk(!wire_dqs_0_enable_inst_dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(bidir_dq_input_data_out_low[1]),
	.regouthi(bidir_dq_input_data_out_high[1]),
	.dfflo());
defparam bidir_dq_1_ddio_in_inst.async_mode = "none";
defparam bidir_dq_1_ddio_in_inst.power_up = "low";
defparam bidir_dq_1_ddio_in_inst.sync_mode = "none";
defparam bidir_dq_1_ddio_in_inst.use_clkn = "false";

arriaii_ddio_in bidir_dq_2_ddio_in_inst(
	.datain(bidir_dq_input_data_in[2]),
	.clk(!wire_dqs_0_enable_inst_dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(bidir_dq_input_data_out_low[2]),
	.regouthi(bidir_dq_input_data_out_high[2]),
	.dfflo());
defparam bidir_dq_2_ddio_in_inst.async_mode = "none";
defparam bidir_dq_2_ddio_in_inst.power_up = "low";
defparam bidir_dq_2_ddio_in_inst.sync_mode = "none";
defparam bidir_dq_2_ddio_in_inst.use_clkn = "false";

arriaii_ddio_in bidir_dq_3_ddio_in_inst(
	.datain(bidir_dq_input_data_in[3]),
	.clk(!wire_dqs_0_enable_inst_dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(bidir_dq_input_data_out_low[3]),
	.regouthi(bidir_dq_input_data_out_high[3]),
	.dfflo());
defparam bidir_dq_3_ddio_in_inst.async_mode = "none";
defparam bidir_dq_3_ddio_in_inst.power_up = "low";
defparam bidir_dq_3_ddio_in_inst.sync_mode = "none";
defparam bidir_dq_3_ddio_in_inst.use_clkn = "false";

arriaii_ddio_in bidir_dq_4_ddio_in_inst(
	.datain(bidir_dq_input_data_in[4]),
	.clk(!wire_dqs_0_enable_inst_dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(bidir_dq_input_data_out_low[4]),
	.regouthi(bidir_dq_input_data_out_high[4]),
	.dfflo());
defparam bidir_dq_4_ddio_in_inst.async_mode = "none";
defparam bidir_dq_4_ddio_in_inst.power_up = "low";
defparam bidir_dq_4_ddio_in_inst.sync_mode = "none";
defparam bidir_dq_4_ddio_in_inst.use_clkn = "false";

arriaii_ddio_in bidir_dq_5_ddio_in_inst(
	.datain(bidir_dq_input_data_in[5]),
	.clk(!wire_dqs_0_enable_inst_dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(bidir_dq_input_data_out_low[5]),
	.regouthi(bidir_dq_input_data_out_high[5]),
	.dfflo());
defparam bidir_dq_5_ddio_in_inst.async_mode = "none";
defparam bidir_dq_5_ddio_in_inst.power_up = "low";
defparam bidir_dq_5_ddio_in_inst.sync_mode = "none";
defparam bidir_dq_5_ddio_in_inst.use_clkn = "false";

arriaii_ddio_in bidir_dq_6_ddio_in_inst(
	.datain(bidir_dq_input_data_in[6]),
	.clk(!wire_dqs_0_enable_inst_dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(bidir_dq_input_data_out_low[6]),
	.regouthi(bidir_dq_input_data_out_high[6]),
	.dfflo());
defparam bidir_dq_6_ddio_in_inst.async_mode = "none";
defparam bidir_dq_6_ddio_in_inst.power_up = "low";
defparam bidir_dq_6_ddio_in_inst.sync_mode = "none";
defparam bidir_dq_6_ddio_in_inst.use_clkn = "false";

arriaii_ddio_in bidir_dq_7_ddio_in_inst(
	.datain(bidir_dq_input_data_in[7]),
	.clk(!wire_dqs_0_enable_inst_dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(bidir_dq_input_data_out_low[7]),
	.regouthi(bidir_dq_input_data_out_high[7]),
	.dfflo());
defparam bidir_dq_7_ddio_in_inst.async_mode = "none";
defparam bidir_dq_7_ddio_in_inst.power_up = "low";
defparam bidir_dq_7_ddio_in_inst.sync_mode = "none";
defparam bidir_dq_7_ddio_in_inst.use_clkn = "false";

arriaii_ddio_out dqs_0_output_ddio_out_inst(
	.datainlo(gnd),
	.datainhi(dqs_output_data_in_high[0]),
	.clkhi(dqs_output_reg_clk),
	.clklo(dqs_output_reg_clk),
	.muxsel(dqs_output_reg_clk),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.clk(gnd),
	.dataout(dqs_output_data_out[0]),
	.dfflo(),
	.dffhi());
defparam dqs_0_output_ddio_out_inst.async_mode = "none";
defparam dqs_0_output_ddio_out_inst.power_up = "low";
defparam dqs_0_output_ddio_out_inst.sync_mode = "none";
defparam dqs_0_output_ddio_out_inst.use_new_clocking_model = "true";

dffeas bidir_dq_0_oe_ff_inst(
	.clk(dq_output_reg_clk),
	.d(\bidir_dq_0_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(bidir_dq_0_oe_ff_inst1),
	.prn(vcc));
defparam bidir_dq_0_oe_ff_inst.is_wysiwyg = "true";
defparam bidir_dq_0_oe_ff_inst.power_up = "low";

dffeas bidir_dq_1_oe_ff_inst(
	.clk(dq_output_reg_clk),
	.d(\bidir_dq_1_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(bidir_dq_1_oe_ff_inst1),
	.prn(vcc));
defparam bidir_dq_1_oe_ff_inst.is_wysiwyg = "true";
defparam bidir_dq_1_oe_ff_inst.power_up = "low";

dffeas bidir_dq_2_oe_ff_inst(
	.clk(dq_output_reg_clk),
	.d(\bidir_dq_2_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(bidir_dq_2_oe_ff_inst1),
	.prn(vcc));
defparam bidir_dq_2_oe_ff_inst.is_wysiwyg = "true";
defparam bidir_dq_2_oe_ff_inst.power_up = "low";

dffeas bidir_dq_3_oe_ff_inst(
	.clk(dq_output_reg_clk),
	.d(\bidir_dq_3_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(bidir_dq_3_oe_ff_inst1),
	.prn(vcc));
defparam bidir_dq_3_oe_ff_inst.is_wysiwyg = "true";
defparam bidir_dq_3_oe_ff_inst.power_up = "low";

dffeas bidir_dq_4_oe_ff_inst(
	.clk(dq_output_reg_clk),
	.d(\bidir_dq_4_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(bidir_dq_4_oe_ff_inst1),
	.prn(vcc));
defparam bidir_dq_4_oe_ff_inst.is_wysiwyg = "true";
defparam bidir_dq_4_oe_ff_inst.power_up = "low";

dffeas bidir_dq_5_oe_ff_inst(
	.clk(dq_output_reg_clk),
	.d(\bidir_dq_5_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(bidir_dq_5_oe_ff_inst1),
	.prn(vcc));
defparam bidir_dq_5_oe_ff_inst.is_wysiwyg = "true";
defparam bidir_dq_5_oe_ff_inst.power_up = "low";

dffeas bidir_dq_6_oe_ff_inst(
	.clk(dq_output_reg_clk),
	.d(\bidir_dq_6_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(bidir_dq_6_oe_ff_inst1),
	.prn(vcc));
defparam bidir_dq_6_oe_ff_inst.is_wysiwyg = "true";
defparam bidir_dq_6_oe_ff_inst.power_up = "low";

dffeas bidir_dq_7_oe_ff_inst(
	.clk(dq_output_reg_clk),
	.d(\bidir_dq_7_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(bidir_dq_7_oe_ff_inst1),
	.prn(vcc));
defparam bidir_dq_7_oe_ff_inst.is_wysiwyg = "true";
defparam bidir_dq_7_oe_ff_inst.power_up = "low";

dffeas dqs_0_oe_ff_inst(
	.clk(dqs_output_reg_clk),
	.d(\dqs_0_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dqs_0_oe_ff_inst1),
	.prn(vcc));
defparam dqs_0_oe_ff_inst.is_wysiwyg = "true";
defparam dqs_0_oe_ff_inst.power_up = "low";

dffeas dqsn_0_oe_ff_inst(
	.clk(dqs_output_reg_clk),
	.d(\dqsn_0_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dqsn_0_oe_ff_inst1),
	.prn(vcc));
defparam dqsn_0_oe_ff_inst.is_wysiwyg = "true";
defparam dqsn_0_oe_ff_inst.power_up = "low";

arriaii_dqs_delay_chain dqs_0_delay_chain_inst(
	.dqsin(dqs_input_data_in[0]),
	.dqsupdateen(gnd),
	.delayctrlin({dll_delayctrlin[5],dll_delayctrlin[4],dll_delayctrlin[3],dll_delayctrlin[2],dll_delayctrlin[1],dll_delayctrlin[0]}),
	.offsetctrlin(6'b000000),
	.dqsbusout(wire_dqs_0_delay_chain_inst_dqsbusout));
defparam dqs_0_delay_chain_inst.delay_buffer_mode = "high";
defparam dqs_0_delay_chain_inst.dqs_ctrl_latches_enable = "false";
defparam dqs_0_delay_chain_inst.dqs_input_frequency = "3333ps";
defparam dqs_0_delay_chain_inst.dqs_offsetctrl_enable = "false";
defparam dqs_0_delay_chain_inst.dqs_phase_shift = 7200;
defparam dqs_0_delay_chain_inst.phase_setting = 2;
defparam dqs_0_delay_chain_inst.sim_buffer_delay_increment = 10;
defparam dqs_0_delay_chain_inst.sim_high_buffer_intrinsic_delay = 175;
defparam dqs_0_delay_chain_inst.sim_low_buffer_intrinsic_delay = 350;
defparam dqs_0_delay_chain_inst.test_enable = "false";
defparam dqs_0_delay_chain_inst.test_select = 0;

arriaii_dqs_enable_ctrl dqs_0_enable_ctrl_inst(
	.dqsenablein(dqs_enable_ctrl_in),
	.clk(dqs_enable_ctrl_clk),
	.dqsenableout(wire_dqs_0_enable_ctrl_inst_dqsenableout));
defparam dqs_0_enable_ctrl_inst.delay_dqs_enable_by_half_cycle = "true";

arriaii_dqs_enable dqs_0_enable_inst(
	.dqsin(wire_dqs_0_delay_chain_inst_dqsbusout),
	.dqsenable(wire_dqs_0_enable_ctrl_inst_dqsenableout),
	.dqsbusout(wire_dqs_0_enable_inst_dqsbusout));

arriaii_lcell_comb \bidir_dq_0_oe_ff_inst~0 (
	.dataa(!dq_oe_2x_2),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bidir_dq_0_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bidir_dq_0_oe_ff_inst~0 .extended_lut = "off";
defparam \bidir_dq_0_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \bidir_dq_0_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \bidir_dq_1_oe_ff_inst~0 (
	.dataa(!dq_oe_2x_2),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bidir_dq_1_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bidir_dq_1_oe_ff_inst~0 .extended_lut = "off";
defparam \bidir_dq_1_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \bidir_dq_1_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \bidir_dq_2_oe_ff_inst~0 (
	.dataa(!dq_oe_2x_2),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bidir_dq_2_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bidir_dq_2_oe_ff_inst~0 .extended_lut = "off";
defparam \bidir_dq_2_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \bidir_dq_2_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \bidir_dq_3_oe_ff_inst~0 (
	.dataa(!dq_oe_2x_2),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bidir_dq_3_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bidir_dq_3_oe_ff_inst~0 .extended_lut = "off";
defparam \bidir_dq_3_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \bidir_dq_3_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \bidir_dq_4_oe_ff_inst~0 (
	.dataa(!dq_oe_2x_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bidir_dq_4_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bidir_dq_4_oe_ff_inst~0 .extended_lut = "off";
defparam \bidir_dq_4_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \bidir_dq_4_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \bidir_dq_5_oe_ff_inst~0 (
	.dataa(!dq_oe_2x_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bidir_dq_5_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bidir_dq_5_oe_ff_inst~0 .extended_lut = "off";
defparam \bidir_dq_5_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \bidir_dq_5_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \bidir_dq_6_oe_ff_inst~0 (
	.dataa(!dq_oe_2x_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bidir_dq_6_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bidir_dq_6_oe_ff_inst~0 .extended_lut = "off";
defparam \bidir_dq_6_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \bidir_dq_6_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \bidir_dq_7_oe_ff_inst~0 (
	.dataa(!dq_oe_2x_3),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bidir_dq_7_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bidir_dq_7_oe_ff_inst~0 .extended_lut = "off";
defparam \bidir_dq_7_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \bidir_dq_7_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \dqs_0_oe_ff_inst~0 (
	.dataa(!dqs_output_data_in_high[0]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dqs_0_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dqs_0_oe_ff_inst~0 .extended_lut = "off";
defparam \dqs_0_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dqs_0_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \dqsn_0_oe_ff_inst~0 (
	.dataa(!dqs_output_data_in_high[0]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dqsn_0_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dqsn_0_oe_ff_inst~0 .extended_lut = "off";
defparam \dqsn_0_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dqsn_0_oe_ff_inst~0 .shared_arith = "off";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_dq_dqs_2 (
	dqs_output_reg_clk,
	dq_output_reg_clk,
	dqs_enable_ctrl_clk,
	dll_delayctrlin,
	output_dq_output_data_out,
	output_dq_output_data_in_low,
	output_dq_output_data_in_high,
	bidir_dq_output_data_out,
	bidir_dq_input_data_out_low,
	bidir_dq_input_data_out_high,
	bidir_dq_output_data_in_low,
	bidir_dq_output_data_in_high,
	dq_oe_2x_4,
	dq_oe_2x_5,
	dqs_output_data_out,
	bidir_dq_input_data_in,
	dqs_input_data_in,
	bidir_dq_0_oe_ff_inst1,
	bidir_dq_1_oe_ff_inst1,
	bidir_dq_2_oe_ff_inst1,
	bidir_dq_3_oe_ff_inst1,
	bidir_dq_4_oe_ff_inst1,
	bidir_dq_5_oe_ff_inst1,
	bidir_dq_6_oe_ff_inst1,
	bidir_dq_7_oe_ff_inst1,
	dqs_0_oe_ff_inst1,
	dqsn_0_oe_ff_inst1,
	bidir_dq_areset,
	dqs_output_data_in_high,
	dqs_enable_ctrl_in)/* synthesis synthesis_greybox=0 */;
input 	dqs_output_reg_clk;
input 	dq_output_reg_clk;
input 	dqs_enable_ctrl_clk;
input 	[5:0] dll_delayctrlin;
output 	[0:0] output_dq_output_data_out;
input 	[0:0] output_dq_output_data_in_low;
input 	[0:0] output_dq_output_data_in_high;
output 	[7:0] bidir_dq_output_data_out;
output 	[7:0] bidir_dq_input_data_out_low;
output 	[7:0] bidir_dq_input_data_out_high;
input 	[7:0] bidir_dq_output_data_in_low;
input 	[7:0] bidir_dq_output_data_in_high;
input 	dq_oe_2x_4;
input 	dq_oe_2x_5;
output 	[0:0] dqs_output_data_out;
input 	[7:0] bidir_dq_input_data_in;
input 	[0:0] dqs_input_data_in;
output 	bidir_dq_0_oe_ff_inst1;
output 	bidir_dq_1_oe_ff_inst1;
output 	bidir_dq_2_oe_ff_inst1;
output 	bidir_dq_3_oe_ff_inst1;
output 	bidir_dq_4_oe_ff_inst1;
output 	bidir_dq_5_oe_ff_inst1;
output 	bidir_dq_6_oe_ff_inst1;
output 	bidir_dq_7_oe_ff_inst1;
output 	dqs_0_oe_ff_inst1;
output 	dqsn_0_oe_ff_inst1;
input 	[7:0] bidir_dq_areset;
input 	[0:0] dqs_output_data_in_high;
input 	dqs_enable_ctrl_in;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire wire_dqs_0_delay_chain_inst_dqsbusout;
wire wire_dqs_0_enable_ctrl_inst_dqsenableout;
wire wire_dqs_0_enable_inst_dqsbusout;
wire \bidir_dq_0_oe_ff_inst~0_combout ;
wire \bidir_dq_1_oe_ff_inst~0_combout ;
wire \bidir_dq_2_oe_ff_inst~0_combout ;
wire \bidir_dq_3_oe_ff_inst~0_combout ;
wire \bidir_dq_4_oe_ff_inst~0_combout ;
wire \bidir_dq_5_oe_ff_inst~0_combout ;
wire \bidir_dq_6_oe_ff_inst~0_combout ;
wire \bidir_dq_7_oe_ff_inst~0_combout ;
wire \dqs_0_oe_ff_inst~0_combout ;
wire \dqsn_0_oe_ff_inst~0_combout ;


arriaii_ddio_out output_dq_0_output_ddio_out_inst(
	.datainlo(output_dq_output_data_in_low[0]),
	.datainhi(output_dq_output_data_in_high[0]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.clk(gnd),
	.dataout(output_dq_output_data_out[0]),
	.dfflo(),
	.dffhi());
defparam output_dq_0_output_ddio_out_inst.async_mode = "clear";
defparam output_dq_0_output_ddio_out_inst.power_up = "low";
defparam output_dq_0_output_ddio_out_inst.sync_mode = "none";
defparam output_dq_0_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_out bidir_dq_0_output_ddio_out_inst(
	.datainlo(bidir_dq_output_data_in_low[0]),
	.datainhi(bidir_dq_output_data_in_high[0]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(!bidir_dq_areset[1]),
	.sreset(gnd),
	.clk(gnd),
	.dataout(bidir_dq_output_data_out[0]),
	.dfflo(),
	.dffhi());
defparam bidir_dq_0_output_ddio_out_inst.async_mode = "clear";
defparam bidir_dq_0_output_ddio_out_inst.power_up = "low";
defparam bidir_dq_0_output_ddio_out_inst.sync_mode = "none";
defparam bidir_dq_0_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_out bidir_dq_1_output_ddio_out_inst(
	.datainlo(bidir_dq_output_data_in_low[1]),
	.datainhi(bidir_dq_output_data_in_high[1]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(!bidir_dq_areset[1]),
	.sreset(gnd),
	.clk(gnd),
	.dataout(bidir_dq_output_data_out[1]),
	.dfflo(),
	.dffhi());
defparam bidir_dq_1_output_ddio_out_inst.async_mode = "clear";
defparam bidir_dq_1_output_ddio_out_inst.power_up = "low";
defparam bidir_dq_1_output_ddio_out_inst.sync_mode = "none";
defparam bidir_dq_1_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_out bidir_dq_2_output_ddio_out_inst(
	.datainlo(bidir_dq_output_data_in_low[2]),
	.datainhi(bidir_dq_output_data_in_high[2]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(!bidir_dq_areset[1]),
	.sreset(gnd),
	.clk(gnd),
	.dataout(bidir_dq_output_data_out[2]),
	.dfflo(),
	.dffhi());
defparam bidir_dq_2_output_ddio_out_inst.async_mode = "clear";
defparam bidir_dq_2_output_ddio_out_inst.power_up = "low";
defparam bidir_dq_2_output_ddio_out_inst.sync_mode = "none";
defparam bidir_dq_2_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_out bidir_dq_3_output_ddio_out_inst(
	.datainlo(bidir_dq_output_data_in_low[3]),
	.datainhi(bidir_dq_output_data_in_high[3]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(!bidir_dq_areset[1]),
	.sreset(gnd),
	.clk(gnd),
	.dataout(bidir_dq_output_data_out[3]),
	.dfflo(),
	.dffhi());
defparam bidir_dq_3_output_ddio_out_inst.async_mode = "clear";
defparam bidir_dq_3_output_ddio_out_inst.power_up = "low";
defparam bidir_dq_3_output_ddio_out_inst.sync_mode = "none";
defparam bidir_dq_3_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_out bidir_dq_4_output_ddio_out_inst(
	.datainlo(bidir_dq_output_data_in_low[4]),
	.datainhi(bidir_dq_output_data_in_high[4]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(!bidir_dq_areset[1]),
	.sreset(gnd),
	.clk(gnd),
	.dataout(bidir_dq_output_data_out[4]),
	.dfflo(),
	.dffhi());
defparam bidir_dq_4_output_ddio_out_inst.async_mode = "clear";
defparam bidir_dq_4_output_ddio_out_inst.power_up = "low";
defparam bidir_dq_4_output_ddio_out_inst.sync_mode = "none";
defparam bidir_dq_4_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_out bidir_dq_5_output_ddio_out_inst(
	.datainlo(bidir_dq_output_data_in_low[5]),
	.datainhi(bidir_dq_output_data_in_high[5]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(!bidir_dq_areset[1]),
	.sreset(gnd),
	.clk(gnd),
	.dataout(bidir_dq_output_data_out[5]),
	.dfflo(),
	.dffhi());
defparam bidir_dq_5_output_ddio_out_inst.async_mode = "clear";
defparam bidir_dq_5_output_ddio_out_inst.power_up = "low";
defparam bidir_dq_5_output_ddio_out_inst.sync_mode = "none";
defparam bidir_dq_5_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_out bidir_dq_6_output_ddio_out_inst(
	.datainlo(bidir_dq_output_data_in_low[6]),
	.datainhi(bidir_dq_output_data_in_high[6]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(!bidir_dq_areset[1]),
	.sreset(gnd),
	.clk(gnd),
	.dataout(bidir_dq_output_data_out[6]),
	.dfflo(),
	.dffhi());
defparam bidir_dq_6_output_ddio_out_inst.async_mode = "clear";
defparam bidir_dq_6_output_ddio_out_inst.power_up = "low";
defparam bidir_dq_6_output_ddio_out_inst.sync_mode = "none";
defparam bidir_dq_6_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_out bidir_dq_7_output_ddio_out_inst(
	.datainlo(bidir_dq_output_data_in_low[7]),
	.datainhi(bidir_dq_output_data_in_high[7]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(!bidir_dq_areset[1]),
	.sreset(gnd),
	.clk(gnd),
	.dataout(bidir_dq_output_data_out[7]),
	.dfflo(),
	.dffhi());
defparam bidir_dq_7_output_ddio_out_inst.async_mode = "clear";
defparam bidir_dq_7_output_ddio_out_inst.power_up = "low";
defparam bidir_dq_7_output_ddio_out_inst.sync_mode = "none";
defparam bidir_dq_7_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_in bidir_dq_0_ddio_in_inst(
	.datain(bidir_dq_input_data_in[0]),
	.clk(!wire_dqs_0_enable_inst_dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(bidir_dq_input_data_out_low[0]),
	.regouthi(bidir_dq_input_data_out_high[0]),
	.dfflo());
defparam bidir_dq_0_ddio_in_inst.async_mode = "none";
defparam bidir_dq_0_ddio_in_inst.power_up = "low";
defparam bidir_dq_0_ddio_in_inst.sync_mode = "none";
defparam bidir_dq_0_ddio_in_inst.use_clkn = "false";

arriaii_ddio_in bidir_dq_1_ddio_in_inst(
	.datain(bidir_dq_input_data_in[1]),
	.clk(!wire_dqs_0_enable_inst_dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(bidir_dq_input_data_out_low[1]),
	.regouthi(bidir_dq_input_data_out_high[1]),
	.dfflo());
defparam bidir_dq_1_ddio_in_inst.async_mode = "none";
defparam bidir_dq_1_ddio_in_inst.power_up = "low";
defparam bidir_dq_1_ddio_in_inst.sync_mode = "none";
defparam bidir_dq_1_ddio_in_inst.use_clkn = "false";

arriaii_ddio_in bidir_dq_2_ddio_in_inst(
	.datain(bidir_dq_input_data_in[2]),
	.clk(!wire_dqs_0_enable_inst_dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(bidir_dq_input_data_out_low[2]),
	.regouthi(bidir_dq_input_data_out_high[2]),
	.dfflo());
defparam bidir_dq_2_ddio_in_inst.async_mode = "none";
defparam bidir_dq_2_ddio_in_inst.power_up = "low";
defparam bidir_dq_2_ddio_in_inst.sync_mode = "none";
defparam bidir_dq_2_ddio_in_inst.use_clkn = "false";

arriaii_ddio_in bidir_dq_3_ddio_in_inst(
	.datain(bidir_dq_input_data_in[3]),
	.clk(!wire_dqs_0_enable_inst_dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(bidir_dq_input_data_out_low[3]),
	.regouthi(bidir_dq_input_data_out_high[3]),
	.dfflo());
defparam bidir_dq_3_ddio_in_inst.async_mode = "none";
defparam bidir_dq_3_ddio_in_inst.power_up = "low";
defparam bidir_dq_3_ddio_in_inst.sync_mode = "none";
defparam bidir_dq_3_ddio_in_inst.use_clkn = "false";

arriaii_ddio_in bidir_dq_4_ddio_in_inst(
	.datain(bidir_dq_input_data_in[4]),
	.clk(!wire_dqs_0_enable_inst_dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(bidir_dq_input_data_out_low[4]),
	.regouthi(bidir_dq_input_data_out_high[4]),
	.dfflo());
defparam bidir_dq_4_ddio_in_inst.async_mode = "none";
defparam bidir_dq_4_ddio_in_inst.power_up = "low";
defparam bidir_dq_4_ddio_in_inst.sync_mode = "none";
defparam bidir_dq_4_ddio_in_inst.use_clkn = "false";

arriaii_ddio_in bidir_dq_5_ddio_in_inst(
	.datain(bidir_dq_input_data_in[5]),
	.clk(!wire_dqs_0_enable_inst_dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(bidir_dq_input_data_out_low[5]),
	.regouthi(bidir_dq_input_data_out_high[5]),
	.dfflo());
defparam bidir_dq_5_ddio_in_inst.async_mode = "none";
defparam bidir_dq_5_ddio_in_inst.power_up = "low";
defparam bidir_dq_5_ddio_in_inst.sync_mode = "none";
defparam bidir_dq_5_ddio_in_inst.use_clkn = "false";

arriaii_ddio_in bidir_dq_6_ddio_in_inst(
	.datain(bidir_dq_input_data_in[6]),
	.clk(!wire_dqs_0_enable_inst_dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(bidir_dq_input_data_out_low[6]),
	.regouthi(bidir_dq_input_data_out_high[6]),
	.dfflo());
defparam bidir_dq_6_ddio_in_inst.async_mode = "none";
defparam bidir_dq_6_ddio_in_inst.power_up = "low";
defparam bidir_dq_6_ddio_in_inst.sync_mode = "none";
defparam bidir_dq_6_ddio_in_inst.use_clkn = "false";

arriaii_ddio_in bidir_dq_7_ddio_in_inst(
	.datain(bidir_dq_input_data_in[7]),
	.clk(!wire_dqs_0_enable_inst_dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(bidir_dq_input_data_out_low[7]),
	.regouthi(bidir_dq_input_data_out_high[7]),
	.dfflo());
defparam bidir_dq_7_ddio_in_inst.async_mode = "none";
defparam bidir_dq_7_ddio_in_inst.power_up = "low";
defparam bidir_dq_7_ddio_in_inst.sync_mode = "none";
defparam bidir_dq_7_ddio_in_inst.use_clkn = "false";

arriaii_ddio_out dqs_0_output_ddio_out_inst(
	.datainlo(gnd),
	.datainhi(dqs_output_data_in_high[0]),
	.clkhi(dqs_output_reg_clk),
	.clklo(dqs_output_reg_clk),
	.muxsel(dqs_output_reg_clk),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.clk(gnd),
	.dataout(dqs_output_data_out[0]),
	.dfflo(),
	.dffhi());
defparam dqs_0_output_ddio_out_inst.async_mode = "none";
defparam dqs_0_output_ddio_out_inst.power_up = "low";
defparam dqs_0_output_ddio_out_inst.sync_mode = "none";
defparam dqs_0_output_ddio_out_inst.use_new_clocking_model = "true";

dffeas bidir_dq_0_oe_ff_inst(
	.clk(dq_output_reg_clk),
	.d(\bidir_dq_0_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(bidir_dq_0_oe_ff_inst1),
	.prn(vcc));
defparam bidir_dq_0_oe_ff_inst.is_wysiwyg = "true";
defparam bidir_dq_0_oe_ff_inst.power_up = "low";

dffeas bidir_dq_1_oe_ff_inst(
	.clk(dq_output_reg_clk),
	.d(\bidir_dq_1_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(bidir_dq_1_oe_ff_inst1),
	.prn(vcc));
defparam bidir_dq_1_oe_ff_inst.is_wysiwyg = "true";
defparam bidir_dq_1_oe_ff_inst.power_up = "low";

dffeas bidir_dq_2_oe_ff_inst(
	.clk(dq_output_reg_clk),
	.d(\bidir_dq_2_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(bidir_dq_2_oe_ff_inst1),
	.prn(vcc));
defparam bidir_dq_2_oe_ff_inst.is_wysiwyg = "true";
defparam bidir_dq_2_oe_ff_inst.power_up = "low";

dffeas bidir_dq_3_oe_ff_inst(
	.clk(dq_output_reg_clk),
	.d(\bidir_dq_3_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(bidir_dq_3_oe_ff_inst1),
	.prn(vcc));
defparam bidir_dq_3_oe_ff_inst.is_wysiwyg = "true";
defparam bidir_dq_3_oe_ff_inst.power_up = "low";

dffeas bidir_dq_4_oe_ff_inst(
	.clk(dq_output_reg_clk),
	.d(\bidir_dq_4_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(bidir_dq_4_oe_ff_inst1),
	.prn(vcc));
defparam bidir_dq_4_oe_ff_inst.is_wysiwyg = "true";
defparam bidir_dq_4_oe_ff_inst.power_up = "low";

dffeas bidir_dq_5_oe_ff_inst(
	.clk(dq_output_reg_clk),
	.d(\bidir_dq_5_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(bidir_dq_5_oe_ff_inst1),
	.prn(vcc));
defparam bidir_dq_5_oe_ff_inst.is_wysiwyg = "true";
defparam bidir_dq_5_oe_ff_inst.power_up = "low";

dffeas bidir_dq_6_oe_ff_inst(
	.clk(dq_output_reg_clk),
	.d(\bidir_dq_6_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(bidir_dq_6_oe_ff_inst1),
	.prn(vcc));
defparam bidir_dq_6_oe_ff_inst.is_wysiwyg = "true";
defparam bidir_dq_6_oe_ff_inst.power_up = "low";

dffeas bidir_dq_7_oe_ff_inst(
	.clk(dq_output_reg_clk),
	.d(\bidir_dq_7_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(bidir_dq_7_oe_ff_inst1),
	.prn(vcc));
defparam bidir_dq_7_oe_ff_inst.is_wysiwyg = "true";
defparam bidir_dq_7_oe_ff_inst.power_up = "low";

dffeas dqs_0_oe_ff_inst(
	.clk(dqs_output_reg_clk),
	.d(\dqs_0_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dqs_0_oe_ff_inst1),
	.prn(vcc));
defparam dqs_0_oe_ff_inst.is_wysiwyg = "true";
defparam dqs_0_oe_ff_inst.power_up = "low";

dffeas dqsn_0_oe_ff_inst(
	.clk(dqs_output_reg_clk),
	.d(\dqsn_0_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dqsn_0_oe_ff_inst1),
	.prn(vcc));
defparam dqsn_0_oe_ff_inst.is_wysiwyg = "true";
defparam dqsn_0_oe_ff_inst.power_up = "low";

arriaii_dqs_delay_chain dqs_0_delay_chain_inst(
	.dqsin(dqs_input_data_in[0]),
	.dqsupdateen(gnd),
	.delayctrlin({dll_delayctrlin[5],dll_delayctrlin[4],dll_delayctrlin[3],dll_delayctrlin[2],dll_delayctrlin[1],dll_delayctrlin[0]}),
	.offsetctrlin(6'b000000),
	.dqsbusout(wire_dqs_0_delay_chain_inst_dqsbusout));
defparam dqs_0_delay_chain_inst.delay_buffer_mode = "high";
defparam dqs_0_delay_chain_inst.dqs_ctrl_latches_enable = "false";
defparam dqs_0_delay_chain_inst.dqs_input_frequency = "3333ps";
defparam dqs_0_delay_chain_inst.dqs_offsetctrl_enable = "false";
defparam dqs_0_delay_chain_inst.dqs_phase_shift = 7200;
defparam dqs_0_delay_chain_inst.phase_setting = 2;
defparam dqs_0_delay_chain_inst.sim_buffer_delay_increment = 10;
defparam dqs_0_delay_chain_inst.sim_high_buffer_intrinsic_delay = 175;
defparam dqs_0_delay_chain_inst.sim_low_buffer_intrinsic_delay = 350;
defparam dqs_0_delay_chain_inst.test_enable = "false";
defparam dqs_0_delay_chain_inst.test_select = 0;

arriaii_dqs_enable_ctrl dqs_0_enable_ctrl_inst(
	.dqsenablein(dqs_enable_ctrl_in),
	.clk(dqs_enable_ctrl_clk),
	.dqsenableout(wire_dqs_0_enable_ctrl_inst_dqsenableout));
defparam dqs_0_enable_ctrl_inst.delay_dqs_enable_by_half_cycle = "true";

arriaii_dqs_enable dqs_0_enable_inst(
	.dqsin(wire_dqs_0_delay_chain_inst_dqsbusout),
	.dqsenable(wire_dqs_0_enable_ctrl_inst_dqsenableout),
	.dqsbusout(wire_dqs_0_enable_inst_dqsbusout));

arriaii_lcell_comb \bidir_dq_0_oe_ff_inst~0 (
	.dataa(!dq_oe_2x_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bidir_dq_0_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bidir_dq_0_oe_ff_inst~0 .extended_lut = "off";
defparam \bidir_dq_0_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \bidir_dq_0_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \bidir_dq_1_oe_ff_inst~0 (
	.dataa(!dq_oe_2x_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bidir_dq_1_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bidir_dq_1_oe_ff_inst~0 .extended_lut = "off";
defparam \bidir_dq_1_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \bidir_dq_1_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \bidir_dq_2_oe_ff_inst~0 (
	.dataa(!dq_oe_2x_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bidir_dq_2_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bidir_dq_2_oe_ff_inst~0 .extended_lut = "off";
defparam \bidir_dq_2_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \bidir_dq_2_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \bidir_dq_3_oe_ff_inst~0 (
	.dataa(!dq_oe_2x_4),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bidir_dq_3_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bidir_dq_3_oe_ff_inst~0 .extended_lut = "off";
defparam \bidir_dq_3_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \bidir_dq_3_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \bidir_dq_4_oe_ff_inst~0 (
	.dataa(!dq_oe_2x_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bidir_dq_4_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bidir_dq_4_oe_ff_inst~0 .extended_lut = "off";
defparam \bidir_dq_4_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \bidir_dq_4_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \bidir_dq_5_oe_ff_inst~0 (
	.dataa(!dq_oe_2x_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bidir_dq_5_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bidir_dq_5_oe_ff_inst~0 .extended_lut = "off";
defparam \bidir_dq_5_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \bidir_dq_5_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \bidir_dq_6_oe_ff_inst~0 (
	.dataa(!dq_oe_2x_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bidir_dq_6_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bidir_dq_6_oe_ff_inst~0 .extended_lut = "off";
defparam \bidir_dq_6_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \bidir_dq_6_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \bidir_dq_7_oe_ff_inst~0 (
	.dataa(!dq_oe_2x_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bidir_dq_7_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bidir_dq_7_oe_ff_inst~0 .extended_lut = "off";
defparam \bidir_dq_7_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \bidir_dq_7_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \dqs_0_oe_ff_inst~0 (
	.dataa(!dqs_output_data_in_high[0]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dqs_0_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dqs_0_oe_ff_inst~0 .extended_lut = "off";
defparam \dqs_0_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dqs_0_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \dqsn_0_oe_ff_inst~0 (
	.dataa(!dqs_output_data_in_high[0]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dqsn_0_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dqsn_0_oe_ff_inst~0 .extended_lut = "off";
defparam \dqsn_0_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dqsn_0_oe_ff_inst~0 .shared_arith = "off";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_dq_dqs_3 (
	dqs_output_reg_clk,
	dq_output_reg_clk,
	dqs_enable_ctrl_clk,
	dll_delayctrlin,
	output_dq_output_data_out,
	output_dq_output_data_in_low,
	output_dq_output_data_in_high,
	bidir_dq_output_data_out,
	bidir_dq_input_data_out_low,
	bidir_dq_input_data_out_high,
	bidir_dq_output_data_in_low,
	bidir_dq_output_data_in_high,
	dq_oe_2x_6,
	dq_oe_2x_7,
	dqs_output_data_out,
	bidir_dq_input_data_in,
	dqs_input_data_in,
	bidir_dq_0_oe_ff_inst1,
	bidir_dq_1_oe_ff_inst1,
	bidir_dq_2_oe_ff_inst1,
	bidir_dq_3_oe_ff_inst1,
	bidir_dq_4_oe_ff_inst1,
	bidir_dq_5_oe_ff_inst1,
	bidir_dq_6_oe_ff_inst1,
	bidir_dq_7_oe_ff_inst1,
	dqs_0_oe_ff_inst1,
	dqsn_0_oe_ff_inst1,
	bidir_dq_areset,
	dqs_output_data_in_high,
	dqs_enable_ctrl_in)/* synthesis synthesis_greybox=0 */;
input 	dqs_output_reg_clk;
input 	dq_output_reg_clk;
input 	dqs_enable_ctrl_clk;
input 	[5:0] dll_delayctrlin;
output 	[0:0] output_dq_output_data_out;
input 	[0:0] output_dq_output_data_in_low;
input 	[0:0] output_dq_output_data_in_high;
output 	[7:0] bidir_dq_output_data_out;
output 	[7:0] bidir_dq_input_data_out_low;
output 	[7:0] bidir_dq_input_data_out_high;
input 	[7:0] bidir_dq_output_data_in_low;
input 	[7:0] bidir_dq_output_data_in_high;
input 	dq_oe_2x_6;
input 	dq_oe_2x_7;
output 	[0:0] dqs_output_data_out;
input 	[7:0] bidir_dq_input_data_in;
input 	[0:0] dqs_input_data_in;
output 	bidir_dq_0_oe_ff_inst1;
output 	bidir_dq_1_oe_ff_inst1;
output 	bidir_dq_2_oe_ff_inst1;
output 	bidir_dq_3_oe_ff_inst1;
output 	bidir_dq_4_oe_ff_inst1;
output 	bidir_dq_5_oe_ff_inst1;
output 	bidir_dq_6_oe_ff_inst1;
output 	bidir_dq_7_oe_ff_inst1;
output 	dqs_0_oe_ff_inst1;
output 	dqsn_0_oe_ff_inst1;
input 	[7:0] bidir_dq_areset;
input 	[0:0] dqs_output_data_in_high;
input 	dqs_enable_ctrl_in;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire wire_dqs_0_delay_chain_inst_dqsbusout;
wire wire_dqs_0_enable_ctrl_inst_dqsenableout;
wire wire_dqs_0_enable_inst_dqsbusout;
wire \bidir_dq_0_oe_ff_inst~0_combout ;
wire \bidir_dq_1_oe_ff_inst~0_combout ;
wire \bidir_dq_2_oe_ff_inst~0_combout ;
wire \bidir_dq_3_oe_ff_inst~0_combout ;
wire \bidir_dq_4_oe_ff_inst~0_combout ;
wire \bidir_dq_5_oe_ff_inst~0_combout ;
wire \bidir_dq_6_oe_ff_inst~0_combout ;
wire \bidir_dq_7_oe_ff_inst~0_combout ;
wire \dqs_0_oe_ff_inst~0_combout ;
wire \dqsn_0_oe_ff_inst~0_combout ;


arriaii_ddio_out output_dq_0_output_ddio_out_inst(
	.datainlo(output_dq_output_data_in_low[0]),
	.datainhi(output_dq_output_data_in_high[0]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.clk(gnd),
	.dataout(output_dq_output_data_out[0]),
	.dfflo(),
	.dffhi());
defparam output_dq_0_output_ddio_out_inst.async_mode = "clear";
defparam output_dq_0_output_ddio_out_inst.power_up = "low";
defparam output_dq_0_output_ddio_out_inst.sync_mode = "none";
defparam output_dq_0_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_out bidir_dq_0_output_ddio_out_inst(
	.datainlo(bidir_dq_output_data_in_low[0]),
	.datainhi(bidir_dq_output_data_in_high[0]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(!bidir_dq_areset[1]),
	.sreset(gnd),
	.clk(gnd),
	.dataout(bidir_dq_output_data_out[0]),
	.dfflo(),
	.dffhi());
defparam bidir_dq_0_output_ddio_out_inst.async_mode = "clear";
defparam bidir_dq_0_output_ddio_out_inst.power_up = "low";
defparam bidir_dq_0_output_ddio_out_inst.sync_mode = "none";
defparam bidir_dq_0_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_out bidir_dq_1_output_ddio_out_inst(
	.datainlo(bidir_dq_output_data_in_low[1]),
	.datainhi(bidir_dq_output_data_in_high[1]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(!bidir_dq_areset[1]),
	.sreset(gnd),
	.clk(gnd),
	.dataout(bidir_dq_output_data_out[1]),
	.dfflo(),
	.dffhi());
defparam bidir_dq_1_output_ddio_out_inst.async_mode = "clear";
defparam bidir_dq_1_output_ddio_out_inst.power_up = "low";
defparam bidir_dq_1_output_ddio_out_inst.sync_mode = "none";
defparam bidir_dq_1_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_out bidir_dq_2_output_ddio_out_inst(
	.datainlo(bidir_dq_output_data_in_low[2]),
	.datainhi(bidir_dq_output_data_in_high[2]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(!bidir_dq_areset[1]),
	.sreset(gnd),
	.clk(gnd),
	.dataout(bidir_dq_output_data_out[2]),
	.dfflo(),
	.dffhi());
defparam bidir_dq_2_output_ddio_out_inst.async_mode = "clear";
defparam bidir_dq_2_output_ddio_out_inst.power_up = "low";
defparam bidir_dq_2_output_ddio_out_inst.sync_mode = "none";
defparam bidir_dq_2_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_out bidir_dq_3_output_ddio_out_inst(
	.datainlo(bidir_dq_output_data_in_low[3]),
	.datainhi(bidir_dq_output_data_in_high[3]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(!bidir_dq_areset[1]),
	.sreset(gnd),
	.clk(gnd),
	.dataout(bidir_dq_output_data_out[3]),
	.dfflo(),
	.dffhi());
defparam bidir_dq_3_output_ddio_out_inst.async_mode = "clear";
defparam bidir_dq_3_output_ddio_out_inst.power_up = "low";
defparam bidir_dq_3_output_ddio_out_inst.sync_mode = "none";
defparam bidir_dq_3_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_out bidir_dq_4_output_ddio_out_inst(
	.datainlo(bidir_dq_output_data_in_low[4]),
	.datainhi(bidir_dq_output_data_in_high[4]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(!bidir_dq_areset[1]),
	.sreset(gnd),
	.clk(gnd),
	.dataout(bidir_dq_output_data_out[4]),
	.dfflo(),
	.dffhi());
defparam bidir_dq_4_output_ddio_out_inst.async_mode = "clear";
defparam bidir_dq_4_output_ddio_out_inst.power_up = "low";
defparam bidir_dq_4_output_ddio_out_inst.sync_mode = "none";
defparam bidir_dq_4_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_out bidir_dq_5_output_ddio_out_inst(
	.datainlo(bidir_dq_output_data_in_low[5]),
	.datainhi(bidir_dq_output_data_in_high[5]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(!bidir_dq_areset[1]),
	.sreset(gnd),
	.clk(gnd),
	.dataout(bidir_dq_output_data_out[5]),
	.dfflo(),
	.dffhi());
defparam bidir_dq_5_output_ddio_out_inst.async_mode = "clear";
defparam bidir_dq_5_output_ddio_out_inst.power_up = "low";
defparam bidir_dq_5_output_ddio_out_inst.sync_mode = "none";
defparam bidir_dq_5_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_out bidir_dq_6_output_ddio_out_inst(
	.datainlo(bidir_dq_output_data_in_low[6]),
	.datainhi(bidir_dq_output_data_in_high[6]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(!bidir_dq_areset[1]),
	.sreset(gnd),
	.clk(gnd),
	.dataout(bidir_dq_output_data_out[6]),
	.dfflo(),
	.dffhi());
defparam bidir_dq_6_output_ddio_out_inst.async_mode = "clear";
defparam bidir_dq_6_output_ddio_out_inst.power_up = "low";
defparam bidir_dq_6_output_ddio_out_inst.sync_mode = "none";
defparam bidir_dq_6_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_out bidir_dq_7_output_ddio_out_inst(
	.datainlo(bidir_dq_output_data_in_low[7]),
	.datainhi(bidir_dq_output_data_in_high[7]),
	.clkhi(dq_output_reg_clk),
	.clklo(dq_output_reg_clk),
	.muxsel(dq_output_reg_clk),
	.ena(vcc),
	.areset(!bidir_dq_areset[1]),
	.sreset(gnd),
	.clk(gnd),
	.dataout(bidir_dq_output_data_out[7]),
	.dfflo(),
	.dffhi());
defparam bidir_dq_7_output_ddio_out_inst.async_mode = "clear";
defparam bidir_dq_7_output_ddio_out_inst.power_up = "low";
defparam bidir_dq_7_output_ddio_out_inst.sync_mode = "none";
defparam bidir_dq_7_output_ddio_out_inst.use_new_clocking_model = "true";

arriaii_ddio_in bidir_dq_0_ddio_in_inst(
	.datain(bidir_dq_input_data_in[0]),
	.clk(!wire_dqs_0_enable_inst_dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(bidir_dq_input_data_out_low[0]),
	.regouthi(bidir_dq_input_data_out_high[0]),
	.dfflo());
defparam bidir_dq_0_ddio_in_inst.async_mode = "none";
defparam bidir_dq_0_ddio_in_inst.power_up = "low";
defparam bidir_dq_0_ddio_in_inst.sync_mode = "none";
defparam bidir_dq_0_ddio_in_inst.use_clkn = "false";

arriaii_ddio_in bidir_dq_1_ddio_in_inst(
	.datain(bidir_dq_input_data_in[1]),
	.clk(!wire_dqs_0_enable_inst_dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(bidir_dq_input_data_out_low[1]),
	.regouthi(bidir_dq_input_data_out_high[1]),
	.dfflo());
defparam bidir_dq_1_ddio_in_inst.async_mode = "none";
defparam bidir_dq_1_ddio_in_inst.power_up = "low";
defparam bidir_dq_1_ddio_in_inst.sync_mode = "none";
defparam bidir_dq_1_ddio_in_inst.use_clkn = "false";

arriaii_ddio_in bidir_dq_2_ddio_in_inst(
	.datain(bidir_dq_input_data_in[2]),
	.clk(!wire_dqs_0_enable_inst_dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(bidir_dq_input_data_out_low[2]),
	.regouthi(bidir_dq_input_data_out_high[2]),
	.dfflo());
defparam bidir_dq_2_ddio_in_inst.async_mode = "none";
defparam bidir_dq_2_ddio_in_inst.power_up = "low";
defparam bidir_dq_2_ddio_in_inst.sync_mode = "none";
defparam bidir_dq_2_ddio_in_inst.use_clkn = "false";

arriaii_ddio_in bidir_dq_3_ddio_in_inst(
	.datain(bidir_dq_input_data_in[3]),
	.clk(!wire_dqs_0_enable_inst_dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(bidir_dq_input_data_out_low[3]),
	.regouthi(bidir_dq_input_data_out_high[3]),
	.dfflo());
defparam bidir_dq_3_ddio_in_inst.async_mode = "none";
defparam bidir_dq_3_ddio_in_inst.power_up = "low";
defparam bidir_dq_3_ddio_in_inst.sync_mode = "none";
defparam bidir_dq_3_ddio_in_inst.use_clkn = "false";

arriaii_ddio_in bidir_dq_4_ddio_in_inst(
	.datain(bidir_dq_input_data_in[4]),
	.clk(!wire_dqs_0_enable_inst_dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(bidir_dq_input_data_out_low[4]),
	.regouthi(bidir_dq_input_data_out_high[4]),
	.dfflo());
defparam bidir_dq_4_ddio_in_inst.async_mode = "none";
defparam bidir_dq_4_ddio_in_inst.power_up = "low";
defparam bidir_dq_4_ddio_in_inst.sync_mode = "none";
defparam bidir_dq_4_ddio_in_inst.use_clkn = "false";

arriaii_ddio_in bidir_dq_5_ddio_in_inst(
	.datain(bidir_dq_input_data_in[5]),
	.clk(!wire_dqs_0_enable_inst_dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(bidir_dq_input_data_out_low[5]),
	.regouthi(bidir_dq_input_data_out_high[5]),
	.dfflo());
defparam bidir_dq_5_ddio_in_inst.async_mode = "none";
defparam bidir_dq_5_ddio_in_inst.power_up = "low";
defparam bidir_dq_5_ddio_in_inst.sync_mode = "none";
defparam bidir_dq_5_ddio_in_inst.use_clkn = "false";

arriaii_ddio_in bidir_dq_6_ddio_in_inst(
	.datain(bidir_dq_input_data_in[6]),
	.clk(!wire_dqs_0_enable_inst_dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(bidir_dq_input_data_out_low[6]),
	.regouthi(bidir_dq_input_data_out_high[6]),
	.dfflo());
defparam bidir_dq_6_ddio_in_inst.async_mode = "none";
defparam bidir_dq_6_ddio_in_inst.power_up = "low";
defparam bidir_dq_6_ddio_in_inst.sync_mode = "none";
defparam bidir_dq_6_ddio_in_inst.use_clkn = "false";

arriaii_ddio_in bidir_dq_7_ddio_in_inst(
	.datain(bidir_dq_input_data_in[7]),
	.clk(!wire_dqs_0_enable_inst_dqsbusout),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(bidir_dq_input_data_out_low[7]),
	.regouthi(bidir_dq_input_data_out_high[7]),
	.dfflo());
defparam bidir_dq_7_ddio_in_inst.async_mode = "none";
defparam bidir_dq_7_ddio_in_inst.power_up = "low";
defparam bidir_dq_7_ddio_in_inst.sync_mode = "none";
defparam bidir_dq_7_ddio_in_inst.use_clkn = "false";

arriaii_ddio_out dqs_0_output_ddio_out_inst(
	.datainlo(gnd),
	.datainhi(dqs_output_data_in_high[0]),
	.clkhi(dqs_output_reg_clk),
	.clklo(dqs_output_reg_clk),
	.muxsel(dqs_output_reg_clk),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.clk(gnd),
	.dataout(dqs_output_data_out[0]),
	.dfflo(),
	.dffhi());
defparam dqs_0_output_ddio_out_inst.async_mode = "none";
defparam dqs_0_output_ddio_out_inst.power_up = "low";
defparam dqs_0_output_ddio_out_inst.sync_mode = "none";
defparam dqs_0_output_ddio_out_inst.use_new_clocking_model = "true";

dffeas bidir_dq_0_oe_ff_inst(
	.clk(dq_output_reg_clk),
	.d(\bidir_dq_0_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(bidir_dq_0_oe_ff_inst1),
	.prn(vcc));
defparam bidir_dq_0_oe_ff_inst.is_wysiwyg = "true";
defparam bidir_dq_0_oe_ff_inst.power_up = "low";

dffeas bidir_dq_1_oe_ff_inst(
	.clk(dq_output_reg_clk),
	.d(\bidir_dq_1_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(bidir_dq_1_oe_ff_inst1),
	.prn(vcc));
defparam bidir_dq_1_oe_ff_inst.is_wysiwyg = "true";
defparam bidir_dq_1_oe_ff_inst.power_up = "low";

dffeas bidir_dq_2_oe_ff_inst(
	.clk(dq_output_reg_clk),
	.d(\bidir_dq_2_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(bidir_dq_2_oe_ff_inst1),
	.prn(vcc));
defparam bidir_dq_2_oe_ff_inst.is_wysiwyg = "true";
defparam bidir_dq_2_oe_ff_inst.power_up = "low";

dffeas bidir_dq_3_oe_ff_inst(
	.clk(dq_output_reg_clk),
	.d(\bidir_dq_3_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(bidir_dq_3_oe_ff_inst1),
	.prn(vcc));
defparam bidir_dq_3_oe_ff_inst.is_wysiwyg = "true";
defparam bidir_dq_3_oe_ff_inst.power_up = "low";

dffeas bidir_dq_4_oe_ff_inst(
	.clk(dq_output_reg_clk),
	.d(\bidir_dq_4_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(bidir_dq_4_oe_ff_inst1),
	.prn(vcc));
defparam bidir_dq_4_oe_ff_inst.is_wysiwyg = "true";
defparam bidir_dq_4_oe_ff_inst.power_up = "low";

dffeas bidir_dq_5_oe_ff_inst(
	.clk(dq_output_reg_clk),
	.d(\bidir_dq_5_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(bidir_dq_5_oe_ff_inst1),
	.prn(vcc));
defparam bidir_dq_5_oe_ff_inst.is_wysiwyg = "true";
defparam bidir_dq_5_oe_ff_inst.power_up = "low";

dffeas bidir_dq_6_oe_ff_inst(
	.clk(dq_output_reg_clk),
	.d(\bidir_dq_6_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(bidir_dq_6_oe_ff_inst1),
	.prn(vcc));
defparam bidir_dq_6_oe_ff_inst.is_wysiwyg = "true";
defparam bidir_dq_6_oe_ff_inst.power_up = "low";

dffeas bidir_dq_7_oe_ff_inst(
	.clk(dq_output_reg_clk),
	.d(\bidir_dq_7_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(bidir_dq_7_oe_ff_inst1),
	.prn(vcc));
defparam bidir_dq_7_oe_ff_inst.is_wysiwyg = "true";
defparam bidir_dq_7_oe_ff_inst.power_up = "low";

dffeas dqs_0_oe_ff_inst(
	.clk(dqs_output_reg_clk),
	.d(\dqs_0_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dqs_0_oe_ff_inst1),
	.prn(vcc));
defparam dqs_0_oe_ff_inst.is_wysiwyg = "true";
defparam dqs_0_oe_ff_inst.power_up = "low";

dffeas dqsn_0_oe_ff_inst(
	.clk(dqs_output_reg_clk),
	.d(\dqsn_0_oe_ff_inst~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dqsn_0_oe_ff_inst1),
	.prn(vcc));
defparam dqsn_0_oe_ff_inst.is_wysiwyg = "true";
defparam dqsn_0_oe_ff_inst.power_up = "low";

arriaii_dqs_delay_chain dqs_0_delay_chain_inst(
	.dqsin(dqs_input_data_in[0]),
	.dqsupdateen(gnd),
	.delayctrlin({dll_delayctrlin[5],dll_delayctrlin[4],dll_delayctrlin[3],dll_delayctrlin[2],dll_delayctrlin[1],dll_delayctrlin[0]}),
	.offsetctrlin(6'b000000),
	.dqsbusout(wire_dqs_0_delay_chain_inst_dqsbusout));
defparam dqs_0_delay_chain_inst.delay_buffer_mode = "high";
defparam dqs_0_delay_chain_inst.dqs_ctrl_latches_enable = "false";
defparam dqs_0_delay_chain_inst.dqs_input_frequency = "3333ps";
defparam dqs_0_delay_chain_inst.dqs_offsetctrl_enable = "false";
defparam dqs_0_delay_chain_inst.dqs_phase_shift = 7200;
defparam dqs_0_delay_chain_inst.phase_setting = 2;
defparam dqs_0_delay_chain_inst.sim_buffer_delay_increment = 10;
defparam dqs_0_delay_chain_inst.sim_high_buffer_intrinsic_delay = 175;
defparam dqs_0_delay_chain_inst.sim_low_buffer_intrinsic_delay = 350;
defparam dqs_0_delay_chain_inst.test_enable = "false";
defparam dqs_0_delay_chain_inst.test_select = 0;

arriaii_dqs_enable_ctrl dqs_0_enable_ctrl_inst(
	.dqsenablein(dqs_enable_ctrl_in),
	.clk(dqs_enable_ctrl_clk),
	.dqsenableout(wire_dqs_0_enable_ctrl_inst_dqsenableout));
defparam dqs_0_enable_ctrl_inst.delay_dqs_enable_by_half_cycle = "true";

arriaii_dqs_enable dqs_0_enable_inst(
	.dqsin(wire_dqs_0_delay_chain_inst_dqsbusout),
	.dqsenable(wire_dqs_0_enable_ctrl_inst_dqsenableout),
	.dqsbusout(wire_dqs_0_enable_inst_dqsbusout));

arriaii_lcell_comb \bidir_dq_0_oe_ff_inst~0 (
	.dataa(!dq_oe_2x_6),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bidir_dq_0_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bidir_dq_0_oe_ff_inst~0 .extended_lut = "off";
defparam \bidir_dq_0_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \bidir_dq_0_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \bidir_dq_1_oe_ff_inst~0 (
	.dataa(!dq_oe_2x_6),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bidir_dq_1_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bidir_dq_1_oe_ff_inst~0 .extended_lut = "off";
defparam \bidir_dq_1_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \bidir_dq_1_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \bidir_dq_2_oe_ff_inst~0 (
	.dataa(!dq_oe_2x_6),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bidir_dq_2_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bidir_dq_2_oe_ff_inst~0 .extended_lut = "off";
defparam \bidir_dq_2_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \bidir_dq_2_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \bidir_dq_3_oe_ff_inst~0 (
	.dataa(!dq_oe_2x_6),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bidir_dq_3_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bidir_dq_3_oe_ff_inst~0 .extended_lut = "off";
defparam \bidir_dq_3_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \bidir_dq_3_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \bidir_dq_4_oe_ff_inst~0 (
	.dataa(!dq_oe_2x_7),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bidir_dq_4_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bidir_dq_4_oe_ff_inst~0 .extended_lut = "off";
defparam \bidir_dq_4_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \bidir_dq_4_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \bidir_dq_5_oe_ff_inst~0 (
	.dataa(!dq_oe_2x_7),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bidir_dq_5_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bidir_dq_5_oe_ff_inst~0 .extended_lut = "off";
defparam \bidir_dq_5_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \bidir_dq_5_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \bidir_dq_6_oe_ff_inst~0 (
	.dataa(!dq_oe_2x_7),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bidir_dq_6_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bidir_dq_6_oe_ff_inst~0 .extended_lut = "off";
defparam \bidir_dq_6_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \bidir_dq_6_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \bidir_dq_7_oe_ff_inst~0 (
	.dataa(!dq_oe_2x_7),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bidir_dq_7_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bidir_dq_7_oe_ff_inst~0 .extended_lut = "off";
defparam \bidir_dq_7_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \bidir_dq_7_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \dqs_0_oe_ff_inst~0 (
	.dataa(!dqs_output_data_in_high[0]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dqs_0_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dqs_0_oe_ff_inst~0 .extended_lut = "off";
defparam \dqs_0_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dqs_0_oe_ff_inst~0 .shared_arith = "off";

arriaii_lcell_comb \dqsn_0_oe_ff_inst~0 (
	.dataa(!dqs_output_data_in_high[0]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dqsn_0_oe_ff_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dqsn_0_oe_ff_inst~0 .extended_lut = "off";
defparam \dqsn_0_oe_ff_inst~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dqsn_0_oe_ff_inst~0 .shared_arith = "off";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_mimic (
	measure_clk,
	mimic_data_in,
	mimic_done_out1,
	reset_measure_clk_n,
	seq_mmc_start,
	mimic_value_captured1)/* synthesis synthesis_greybox=0 */;
input 	measure_clk;
input 	mimic_data_in;
output 	mimic_done_out1;
input 	reset_measure_clk_n;
input 	seq_mmc_start;
output 	mimic_value_captured1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \shift_reg_data_out[2]~q ;
wire \mimic_data_in_metastable[1]~q ;
wire \shift_reg_data_out~3_combout ;
wire \mimic_data_in_metastable[0]~q ;
wire \seq_mmc_start_metastable[0]~q ;
wire \seq_mmc_start_metastable[1]~q ;
wire \seq_mmc_start_metastable[2]~q ;
wire \Selector6~1_combout ;
wire \shift_reg_counter[0]~4_combout ;
wire \shift_reg_counter[0]~q ;
wire \shift_reg_counter[0]~1_combout ;
wire \shift_reg_counter[1]~3_combout ;
wire \shift_reg_counter[1]~q ;
wire \shift_reg_counter[2]~2_combout ;
wire \shift_reg_counter[2]~q ;
wire \Equal0~0_combout ;
wire \Selector7~0_combout ;
wire \mimic_state.001~q ;
wire \Equal0~1_combout ;
wire \shift_reg_counter[3]~0_combout ;
wire \shift_reg_counter[3]~q ;
wire \shift_reg_counter[0]~5_combout ;
wire \mimic_state.010~q ;
wire \mimic_state.011~q ;
wire \mimic_state.100~q ;
wire \Selector6~0_combout ;
wire \mimic_state.000~q ;
wire \Selector4~0_combout ;
wire \shift_reg_s_clr~0_combout ;
wire \shift_reg_s_clr~q ;
wire \shift_reg_data_out~0_combout ;
wire \Selector5~0_combout ;
wire \shift_reg_enable~q ;
wire \shift_reg_data_out[0]~1_combout ;
wire \shift_reg_data_out[0]~q ;
wire \shift_reg_data_out~2_combout ;
wire \shift_reg_data_out[1]~q ;
wire \shift_reg_data_out~4_combout ;
wire \shift_reg_data_out[3]~q ;
wire \shift_reg_data_out~5_combout ;
wire \shift_reg_data_out[5]~q ;
wire \shift_reg_data_out~6_combout ;
wire \shift_reg_data_out[4]~q ;
wire \mimic_value_captured~0_combout ;
wire \mimic_value_captured~1_combout ;


dffeas \shift_reg_data_out[2] (
	.clk(measure_clk),
	.d(\shift_reg_data_out~3_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shift_reg_data_out[0]~1_combout ),
	.q(\shift_reg_data_out[2]~q ),
	.prn(vcc));
defparam \shift_reg_data_out[2] .is_wysiwyg = "true";
defparam \shift_reg_data_out[2] .power_up = "low";

dffeas \mimic_data_in_metastable[1] (
	.clk(measure_clk),
	.d(\mimic_data_in_metastable[0]~q ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mimic_data_in_metastable[1]~q ),
	.prn(vcc));
defparam \mimic_data_in_metastable[1] .is_wysiwyg = "true";
defparam \mimic_data_in_metastable[1] .power_up = "low";

arriaii_lcell_comb \shift_reg_data_out~3 (
	.dataa(!\shift_reg_data_out[1]~q ),
	.datab(!\shift_reg_s_clr~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\shift_reg_data_out~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \shift_reg_data_out~3 .extended_lut = "off";
defparam \shift_reg_data_out~3 .lut_mask = 64'h4444444444444444;
defparam \shift_reg_data_out~3 .shared_arith = "off";

dffeas \mimic_data_in_metastable[0] (
	.clk(measure_clk),
	.d(mimic_data_in),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mimic_data_in_metastable[0]~q ),
	.prn(vcc));
defparam \mimic_data_in_metastable[0] .is_wysiwyg = "true";
defparam \mimic_data_in_metastable[0] .power_up = "low";

dffeas mimic_done_out(
	.clk(measure_clk),
	.d(\Selector4~0_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mimic_done_out1),
	.prn(vcc));
defparam mimic_done_out.is_wysiwyg = "true";
defparam mimic_done_out.power_up = "low";

dffeas mimic_value_captured(
	.clk(measure_clk),
	.d(\mimic_value_captured~1_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mimic_value_captured1),
	.prn(vcc));
defparam mimic_value_captured.is_wysiwyg = "true";
defparam mimic_value_captured.power_up = "low";

dffeas \seq_mmc_start_metastable[0] (
	.clk(measure_clk),
	.d(seq_mmc_start),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_mmc_start_metastable[0]~q ),
	.prn(vcc));
defparam \seq_mmc_start_metastable[0] .is_wysiwyg = "true";
defparam \seq_mmc_start_metastable[0] .power_up = "low";

dffeas \seq_mmc_start_metastable[1] (
	.clk(measure_clk),
	.d(\seq_mmc_start_metastable[0]~q ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_mmc_start_metastable[1]~q ),
	.prn(vcc));
defparam \seq_mmc_start_metastable[1] .is_wysiwyg = "true";
defparam \seq_mmc_start_metastable[1] .power_up = "low";

dffeas \seq_mmc_start_metastable[2] (
	.clk(measure_clk),
	.d(\seq_mmc_start_metastable[1]~q ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_mmc_start_metastable[2]~q ),
	.prn(vcc));
defparam \seq_mmc_start_metastable[2] .is_wysiwyg = "true";
defparam \seq_mmc_start_metastable[2] .power_up = "low";

arriaii_lcell_comb \Selector6~1 (
	.dataa(!\mimic_state.000~q ),
	.datab(!\seq_mmc_start_metastable[2]~q ),
	.datac(!\seq_mmc_start_metastable[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector6~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~1 .extended_lut = "off";
defparam \Selector6~1 .lut_mask = 64'hA2A2A2A2A2A2A2A2;
defparam \Selector6~1 .shared_arith = "off";

arriaii_lcell_comb \shift_reg_counter[0]~4 (
	.dataa(!\mimic_state.000~q ),
	.datab(!\mimic_state.001~q ),
	.datac(!\shift_reg_counter[0]~q ),
	.datad(!\Equal0~0_combout ),
	.datae(!\Selector6~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\shift_reg_counter[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \shift_reg_counter[0]~4 .extended_lut = "off";
defparam \shift_reg_counter[0]~4 .lut_mask = 64'hB4870407B4870407;
defparam \shift_reg_counter[0]~4 .shared_arith = "off";

dffeas \shift_reg_counter[0] (
	.clk(measure_clk),
	.d(\shift_reg_counter[0]~4_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\shift_reg_counter[0]~q ),
	.prn(vcc));
defparam \shift_reg_counter[0] .is_wysiwyg = "true";
defparam \shift_reg_counter[0] .power_up = "low";

arriaii_lcell_comb \shift_reg_counter[0]~1 (
	.dataa(!\mimic_state.000~q ),
	.datab(!\mimic_state.001~q ),
	.datac(!\shift_reg_counter[3]~q ),
	.datad(!\shift_reg_counter[2]~q ),
	.datae(!\shift_reg_counter[1]~q ),
	.dataf(!\shift_reg_counter[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\shift_reg_counter[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \shift_reg_counter[0]~1 .extended_lut = "off";
defparam \shift_reg_counter[0]~1 .lut_mask = 64'h4444444444444474;
defparam \shift_reg_counter[0]~1 .shared_arith = "off";

arriaii_lcell_comb \shift_reg_counter[1]~3 (
	.dataa(!\shift_reg_counter[1]~q ),
	.datab(!\shift_reg_counter[0]~q ),
	.datac(!\Selector6~1_combout ),
	.datad(!\shift_reg_counter[0]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\shift_reg_counter[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \shift_reg_counter[1]~3 .extended_lut = "off";
defparam \shift_reg_counter[1]~3 .lut_mask = 64'h6055605560556055;
defparam \shift_reg_counter[1]~3 .shared_arith = "off";

dffeas \shift_reg_counter[1] (
	.clk(measure_clk),
	.d(\shift_reg_counter[1]~3_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\shift_reg_counter[1]~q ),
	.prn(vcc));
defparam \shift_reg_counter[1] .is_wysiwyg = "true";
defparam \shift_reg_counter[1] .power_up = "low";

arriaii_lcell_comb \shift_reg_counter[2]~2 (
	.dataa(!\shift_reg_counter[2]~q ),
	.datab(!\shift_reg_counter[1]~q ),
	.datac(!\shift_reg_counter[0]~q ),
	.datad(!\Selector6~1_combout ),
	.datae(!\shift_reg_counter[0]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\shift_reg_counter[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \shift_reg_counter[2]~2 .extended_lut = "off";
defparam \shift_reg_counter[2]~2 .lut_mask = 64'h5600555556005555;
defparam \shift_reg_counter[2]~2 .shared_arith = "off";

dffeas \shift_reg_counter[2] (
	.clk(measure_clk),
	.d(\shift_reg_counter[2]~2_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\shift_reg_counter[2]~q ),
	.prn(vcc));
defparam \shift_reg_counter[2] .is_wysiwyg = "true";
defparam \shift_reg_counter[2] .power_up = "low";

arriaii_lcell_comb \Equal0~0 (
	.dataa(!\shift_reg_counter[3]~q ),
	.datab(!\shift_reg_counter[2]~q ),
	.datac(!\shift_reg_counter[1]~q ),
	.datad(!\shift_reg_counter[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h0002000200020002;
defparam \Equal0~0 .shared_arith = "off";

arriaii_lcell_comb \Selector7~0 (
	.dataa(!\mimic_state.000~q ),
	.datab(!\mimic_state.001~q ),
	.datac(!\Equal0~0_combout ),
	.datad(!\seq_mmc_start_metastable[2]~q ),
	.datae(!\seq_mmc_start_metastable[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector7~0 .extended_lut = "off";
defparam \Selector7~0 .lut_mask = 64'h3030BA303030BA30;
defparam \Selector7~0 .shared_arith = "off";

dffeas \mimic_state.001 (
	.clk(measure_clk),
	.d(\Selector7~0_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mimic_state.001~q ),
	.prn(vcc));
defparam \mimic_state.001 .is_wysiwyg = "true";
defparam \mimic_state.001 .power_up = "low";

arriaii_lcell_comb \Equal0~1 (
	.dataa(!\shift_reg_counter[2]~q ),
	.datab(!\shift_reg_counter[1]~q ),
	.datac(!\shift_reg_counter[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~1 .extended_lut = "off";
defparam \Equal0~1 .lut_mask = 64'h0101010101010101;
defparam \Equal0~1 .shared_arith = "off";

arriaii_lcell_comb \shift_reg_counter[3]~0 (
	.dataa(!\mimic_state.000~q ),
	.datab(!\mimic_state.001~q ),
	.datac(!\shift_reg_counter[3]~q ),
	.datad(!\Equal0~1_combout ),
	.datae(!\Selector6~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\shift_reg_counter[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \shift_reg_counter[3]~0 .extended_lut = "off";
defparam \shift_reg_counter[3]~0 .lut_mask = 64'h0F8404040F840404;
defparam \shift_reg_counter[3]~0 .shared_arith = "off";

dffeas \shift_reg_counter[3] (
	.clk(measure_clk),
	.d(\shift_reg_counter[3]~0_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\shift_reg_counter[3]~q ),
	.prn(vcc));
defparam \shift_reg_counter[3] .is_wysiwyg = "true";
defparam \shift_reg_counter[3] .power_up = "low";

arriaii_lcell_comb \shift_reg_counter[0]~5 (
	.dataa(!\mimic_state.001~q ),
	.datab(!\shift_reg_counter[3]~q ),
	.datac(!\shift_reg_counter[2]~q ),
	.datad(!\shift_reg_counter[1]~q ),
	.datae(!\shift_reg_counter[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\shift_reg_counter[0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \shift_reg_counter[0]~5 .extended_lut = "off";
defparam \shift_reg_counter[0]~5 .lut_mask = 64'h0000000400000004;
defparam \shift_reg_counter[0]~5 .shared_arith = "off";

dffeas \mimic_state.010 (
	.clk(measure_clk),
	.d(\shift_reg_counter[0]~5_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mimic_state.010~q ),
	.prn(vcc));
defparam \mimic_state.010 .is_wysiwyg = "true";
defparam \mimic_state.010 .power_up = "low";

dffeas \mimic_state.011 (
	.clk(measure_clk),
	.d(\mimic_state.010~q ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mimic_state.011~q ),
	.prn(vcc));
defparam \mimic_state.011 .is_wysiwyg = "true";
defparam \mimic_state.011 .power_up = "low";

dffeas \mimic_state.100 (
	.clk(measure_clk),
	.d(\mimic_state.011~q ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mimic_state.100~q ),
	.prn(vcc));
defparam \mimic_state.100 .is_wysiwyg = "true";
defparam \mimic_state.100 .power_up = "low";

arriaii_lcell_comb \Selector6~0 (
	.dataa(!\mimic_state.000~q ),
	.datab(!\mimic_state.100~q ),
	.datac(!\seq_mmc_start_metastable[2]~q ),
	.datad(!\seq_mmc_start_metastable[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~0 .extended_lut = "off";
defparam \Selector6~0 .lut_mask = 64'h44C444C444C444C4;
defparam \Selector6~0 .shared_arith = "off";

dffeas \mimic_state.000 (
	.clk(measure_clk),
	.d(\Selector6~0_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mimic_state.000~q ),
	.prn(vcc));
defparam \mimic_state.000 .is_wysiwyg = "true";
defparam \mimic_state.000 .power_up = "low";

arriaii_lcell_comb \Selector4~0 (
	.dataa(!mimic_done_out1),
	.datab(!\mimic_state.000~q ),
	.datac(!\mimic_state.001~q ),
	.datad(!\Equal0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~0 .extended_lut = "off";
defparam \Selector4~0 .lut_mask = 64'h353F353F353F353F;
defparam \Selector4~0 .shared_arith = "off";

arriaii_lcell_comb \shift_reg_s_clr~0 (
	.dataa(!\mimic_state.000~q ),
	.datab(!\seq_mmc_start_metastable[2]~q ),
	.datac(!\seq_mmc_start_metastable[1]~q ),
	.datad(!\shift_reg_s_clr~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\shift_reg_s_clr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \shift_reg_s_clr~0 .extended_lut = "off";
defparam \shift_reg_s_clr~0 .lut_mask = 64'hA2F7A2F7A2F7A2F7;
defparam \shift_reg_s_clr~0 .shared_arith = "off";

dffeas shift_reg_s_clr(
	.clk(measure_clk),
	.d(\shift_reg_s_clr~0_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\shift_reg_s_clr~q ),
	.prn(vcc));
defparam shift_reg_s_clr.is_wysiwyg = "true";
defparam shift_reg_s_clr.power_up = "low";

arriaii_lcell_comb \shift_reg_data_out~0 (
	.dataa(!\mimic_data_in_metastable[1]~q ),
	.datab(!\shift_reg_s_clr~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\shift_reg_data_out~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \shift_reg_data_out~0 .extended_lut = "off";
defparam \shift_reg_data_out~0 .lut_mask = 64'h4444444444444444;
defparam \shift_reg_data_out~0 .shared_arith = "off";

arriaii_lcell_comb \Selector5~0 (
	.dataa(!\mimic_state.000~q ),
	.datab(!\mimic_state.001~q ),
	.datac(!\Equal0~0_combout ),
	.datad(!\shift_reg_enable~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~0 .extended_lut = "off";
defparam \Selector5~0 .lut_mask = 64'h88FC88FC88FC88FC;
defparam \Selector5~0 .shared_arith = "off";

dffeas shift_reg_enable(
	.clk(measure_clk),
	.d(\Selector5~0_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\shift_reg_enable~q ),
	.prn(vcc));
defparam shift_reg_enable.is_wysiwyg = "true";
defparam shift_reg_enable.power_up = "low";

arriaii_lcell_comb \shift_reg_data_out[0]~1 (
	.dataa(!\shift_reg_s_clr~q ),
	.datab(!\shift_reg_enable~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\shift_reg_data_out[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \shift_reg_data_out[0]~1 .extended_lut = "off";
defparam \shift_reg_data_out[0]~1 .lut_mask = 64'h7777777777777777;
defparam \shift_reg_data_out[0]~1 .shared_arith = "off";

dffeas \shift_reg_data_out[0] (
	.clk(measure_clk),
	.d(\shift_reg_data_out~0_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shift_reg_data_out[0]~1_combout ),
	.q(\shift_reg_data_out[0]~q ),
	.prn(vcc));
defparam \shift_reg_data_out[0] .is_wysiwyg = "true";
defparam \shift_reg_data_out[0] .power_up = "low";

arriaii_lcell_comb \shift_reg_data_out~2 (
	.dataa(!\shift_reg_data_out[0]~q ),
	.datab(!\shift_reg_s_clr~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\shift_reg_data_out~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \shift_reg_data_out~2 .extended_lut = "off";
defparam \shift_reg_data_out~2 .lut_mask = 64'h4444444444444444;
defparam \shift_reg_data_out~2 .shared_arith = "off";

dffeas \shift_reg_data_out[1] (
	.clk(measure_clk),
	.d(\shift_reg_data_out~2_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shift_reg_data_out[0]~1_combout ),
	.q(\shift_reg_data_out[1]~q ),
	.prn(vcc));
defparam \shift_reg_data_out[1] .is_wysiwyg = "true";
defparam \shift_reg_data_out[1] .power_up = "low";

arriaii_lcell_comb \shift_reg_data_out~4 (
	.dataa(!\shift_reg_data_out[2]~q ),
	.datab(!\shift_reg_s_clr~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\shift_reg_data_out~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \shift_reg_data_out~4 .extended_lut = "off";
defparam \shift_reg_data_out~4 .lut_mask = 64'h4444444444444444;
defparam \shift_reg_data_out~4 .shared_arith = "off";

dffeas \shift_reg_data_out[3] (
	.clk(measure_clk),
	.d(\shift_reg_data_out~4_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shift_reg_data_out[0]~1_combout ),
	.q(\shift_reg_data_out[3]~q ),
	.prn(vcc));
defparam \shift_reg_data_out[3] .is_wysiwyg = "true";
defparam \shift_reg_data_out[3] .power_up = "low";

arriaii_lcell_comb \shift_reg_data_out~5 (
	.dataa(!\shift_reg_data_out[4]~q ),
	.datab(!\shift_reg_s_clr~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\shift_reg_data_out~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \shift_reg_data_out~5 .extended_lut = "off";
defparam \shift_reg_data_out~5 .lut_mask = 64'h4444444444444444;
defparam \shift_reg_data_out~5 .shared_arith = "off";

dffeas \shift_reg_data_out[5] (
	.clk(measure_clk),
	.d(\shift_reg_data_out~5_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shift_reg_data_out[0]~1_combout ),
	.q(\shift_reg_data_out[5]~q ),
	.prn(vcc));
defparam \shift_reg_data_out[5] .is_wysiwyg = "true";
defparam \shift_reg_data_out[5] .power_up = "low";

arriaii_lcell_comb \shift_reg_data_out~6 (
	.dataa(!\shift_reg_data_out[3]~q ),
	.datab(!\shift_reg_s_clr~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\shift_reg_data_out~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \shift_reg_data_out~6 .extended_lut = "off";
defparam \shift_reg_data_out~6 .lut_mask = 64'h4444444444444444;
defparam \shift_reg_data_out~6 .shared_arith = "off";

dffeas \shift_reg_data_out[4] (
	.clk(measure_clk),
	.d(\shift_reg_data_out~6_combout ),
	.asdata(vcc),
	.clrn(reset_measure_clk_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shift_reg_data_out[0]~1_combout ),
	.q(\shift_reg_data_out[4]~q ),
	.prn(vcc));
defparam \shift_reg_data_out[4] .is_wysiwyg = "true";
defparam \shift_reg_data_out[4] .power_up = "low";

arriaii_lcell_comb \mimic_value_captured~0 (
	.dataa(!\shift_reg_data_out[2]~q ),
	.datab(!\shift_reg_data_out[3]~q ),
	.datac(!\shift_reg_data_out[5]~q ),
	.datad(!\shift_reg_data_out[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mimic_value_captured~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mimic_value_captured~0 .extended_lut = "off";
defparam \mimic_value_captured~0 .lut_mask = 64'h0001000100010001;
defparam \mimic_value_captured~0 .shared_arith = "off";

arriaii_lcell_comb \mimic_value_captured~1 (
	.dataa(!\shift_reg_counter[0]~5_combout ),
	.datab(!mimic_value_captured1),
	.datac(!\shift_reg_data_out[0]~q ),
	.datad(!\shift_reg_data_out[1]~q ),
	.datae(!\mimic_value_captured~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mimic_value_captured~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mimic_value_captured~1 .extended_lut = "off";
defparam \mimic_value_captured~1 .lut_mask = 64'h2222222722222227;
defparam \mimic_value_captured~1 .shared_arith = "off";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_postamble (
	clk_0,
	clk_4,
	rd_addr_2x_0,
	reset_phy_clk_1x_n,
	reset_poa_clk_2x_n,
	seq_rdv_doing_rd_7,
	merged_doing_rd,
	seq_rdv_doing_rd_4,
	postamble_en_pos_2x_0,
	postamble_en_pos_2x_1,
	postamble_en_pos_2x_2,
	postamble_en_pos_2x_3,
	seq_poa_protection_override_1x,
	seq_poa_lat_dec_1x,
	ctl_doing_rd_beat2_1x)/* synthesis synthesis_greybox=0 */;
input 	clk_0;
input 	clk_4;
output 	rd_addr_2x_0;
input 	reset_phy_clk_1x_n;
input 	reset_poa_clk_2x_n;
input 	seq_rdv_doing_rd_7;
input 	merged_doing_rd;
input 	seq_rdv_doing_rd_4;
output 	postamble_en_pos_2x_0;
output 	postamble_en_pos_2x_1;
output 	postamble_en_pos_2x_2;
output 	postamble_en_pos_2x_3;
input 	seq_poa_protection_override_1x;
input 	seq_poa_lat_dec_1x;
input 	ctl_doing_rd_beat2_1x;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \half_rate_ram_gen.altsyncram_inst|auto_generated|q_b[0] ;
wire \Add0~1_sumout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \Add2~1_sumout ;
wire \Add2~2 ;
wire \Add2~5_sumout ;
wire \Add2~6 ;
wire \Add2~9_sumout ;
wire \Add2~10 ;
wire \Add2~13_sumout ;
wire \Add2~14 ;
wire \Add2~17_sumout ;
wire \bit_order_1x~q ;
wire \ctl_doing_rd_beat2_1x_r1~q ;
wire \wr_data_1x[0]~0_combout ;
wire \wr_data_1x[1]~1_combout ;
wire \wr_addr_1x[0]~q ;
wire \wr_addr_1x[1]~q ;
wire \wr_addr_1x[2]~q ;
wire \wr_addr_1x[3]~q ;
wire \wr_addr_1x[4]~q ;
wire \rd_addr_2x[1]~q ;
wire \rd_addr_2x[2]~q ;
wire \rd_addr_2x[3]~q ;
wire \rd_addr_2x[4]~q ;
wire \rd_addr_2x[5]~q ;
wire \seq_poa_lat_dec_1x_1t~q ;
wire \bit_order_1x~0_combout ;
wire \wr_addr_1x[0]~0_combout ;
wire \wr_addr_1x[4]~1_combout ;
wire \wr_addr_1x[4]~_wirecell_combout ;
wire \rd_addr_2x[0]~0_combout ;
wire \postamble_en_2x_r[0]~q ;
wire \postamble_en_2x_r[1]~q ;
wire \postamble_en_2x_r[2]~q ;
wire \postamble_en_2x_r[3]~q ;


ddr3_int_altsyncram_1 \half_rate_ram_gen.altsyncram_inst (
	.clock0(clk_0),
	.clock1(clk_4),
	.q_b({q_b_unconnected_wire_127,q_b_unconnected_wire_126,q_b_unconnected_wire_125,q_b_unconnected_wire_124,q_b_unconnected_wire_123,q_b_unconnected_wire_122,q_b_unconnected_wire_121,q_b_unconnected_wire_120,q_b_unconnected_wire_119,q_b_unconnected_wire_118,
q_b_unconnected_wire_117,q_b_unconnected_wire_116,q_b_unconnected_wire_115,q_b_unconnected_wire_114,q_b_unconnected_wire_113,q_b_unconnected_wire_112,q_b_unconnected_wire_111,q_b_unconnected_wire_110,q_b_unconnected_wire_109,q_b_unconnected_wire_108,
q_b_unconnected_wire_107,q_b_unconnected_wire_106,q_b_unconnected_wire_105,q_b_unconnected_wire_104,q_b_unconnected_wire_103,q_b_unconnected_wire_102,q_b_unconnected_wire_101,q_b_unconnected_wire_100,q_b_unconnected_wire_99,q_b_unconnected_wire_98,
q_b_unconnected_wire_97,q_b_unconnected_wire_96,q_b_unconnected_wire_95,q_b_unconnected_wire_94,q_b_unconnected_wire_93,q_b_unconnected_wire_92,q_b_unconnected_wire_91,q_b_unconnected_wire_90,q_b_unconnected_wire_89,q_b_unconnected_wire_88,q_b_unconnected_wire_87,
q_b_unconnected_wire_86,q_b_unconnected_wire_85,q_b_unconnected_wire_84,q_b_unconnected_wire_83,q_b_unconnected_wire_82,q_b_unconnected_wire_81,q_b_unconnected_wire_80,q_b_unconnected_wire_79,q_b_unconnected_wire_78,q_b_unconnected_wire_77,q_b_unconnected_wire_76,
q_b_unconnected_wire_75,q_b_unconnected_wire_74,q_b_unconnected_wire_73,q_b_unconnected_wire_72,q_b_unconnected_wire_71,q_b_unconnected_wire_70,q_b_unconnected_wire_69,q_b_unconnected_wire_68,q_b_unconnected_wire_67,q_b_unconnected_wire_66,q_b_unconnected_wire_65,
q_b_unconnected_wire_64,q_b_unconnected_wire_63,q_b_unconnected_wire_62,q_b_unconnected_wire_61,q_b_unconnected_wire_60,q_b_unconnected_wire_59,q_b_unconnected_wire_58,q_b_unconnected_wire_57,q_b_unconnected_wire_56,q_b_unconnected_wire_55,q_b_unconnected_wire_54,
q_b_unconnected_wire_53,q_b_unconnected_wire_52,q_b_unconnected_wire_51,q_b_unconnected_wire_50,q_b_unconnected_wire_49,q_b_unconnected_wire_48,q_b_unconnected_wire_47,q_b_unconnected_wire_46,q_b_unconnected_wire_45,q_b_unconnected_wire_44,q_b_unconnected_wire_43,
q_b_unconnected_wire_42,q_b_unconnected_wire_41,q_b_unconnected_wire_40,q_b_unconnected_wire_39,q_b_unconnected_wire_38,q_b_unconnected_wire_37,q_b_unconnected_wire_36,q_b_unconnected_wire_35,q_b_unconnected_wire_34,q_b_unconnected_wire_33,q_b_unconnected_wire_32,
q_b_unconnected_wire_31,q_b_unconnected_wire_30,q_b_unconnected_wire_29,q_b_unconnected_wire_28,q_b_unconnected_wire_27,q_b_unconnected_wire_26,q_b_unconnected_wire_25,q_b_unconnected_wire_24,q_b_unconnected_wire_23,q_b_unconnected_wire_22,q_b_unconnected_wire_21,
q_b_unconnected_wire_20,q_b_unconnected_wire_19,q_b_unconnected_wire_18,q_b_unconnected_wire_17,q_b_unconnected_wire_16,q_b_unconnected_wire_15,q_b_unconnected_wire_14,q_b_unconnected_wire_13,q_b_unconnected_wire_12,q_b_unconnected_wire_11,q_b_unconnected_wire_10,
q_b_unconnected_wire_9,q_b_unconnected_wire_8,q_b_unconnected_wire_7,q_b_unconnected_wire_6,q_b_unconnected_wire_5,q_b_unconnected_wire_4,q_b_unconnected_wire_3,q_b_unconnected_wire_2,q_b_unconnected_wire_1,\half_rate_ram_gen.altsyncram_inst|auto_generated|q_b[0] }),
	.address_b({\rd_addr_2x[5]~q ,\rd_addr_2x[4]~q ,\rd_addr_2x[3]~q ,\rd_addr_2x[2]~q ,\rd_addr_2x[1]~q ,rd_addr_2x_0}),
	.data_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_data_1x[1]~1_combout ,\wr_data_1x[0]~0_combout }),
	.address_a({\wr_addr_1x[4]~_wirecell_combout ,\wr_addr_1x[3]~q ,\wr_addr_1x[2]~q ,\wr_addr_1x[1]~q ,\wr_addr_1x[0]~q }));

arriaii_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\wr_addr_1x[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

arriaii_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\wr_addr_1x[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~5 .shared_arith = "off";

arriaii_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\wr_addr_1x[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~9 .shared_arith = "off";

arriaii_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\wr_addr_1x[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~13 .shared_arith = "off";

arriaii_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\wr_addr_1x[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FFFF0000FF00;
defparam \Add0~17 .shared_arith = "off";

arriaii_lcell_comb \Add2~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!rd_addr_2x_0),
	.datae(gnd),
	.dataf(!\rd_addr_2x[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~1_sumout ),
	.cout(\Add2~2 ),
	.shareout());
defparam \Add2~1 .extended_lut = "off";
defparam \Add2~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add2~1 .shared_arith = "off";

arriaii_lcell_comb \Add2~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\rd_addr_2x[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~5_sumout ),
	.cout(\Add2~6 ),
	.shareout());
defparam \Add2~5 .extended_lut = "off";
defparam \Add2~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add2~5 .shared_arith = "off";

arriaii_lcell_comb \Add2~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\rd_addr_2x[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~9_sumout ),
	.cout(\Add2~10 ),
	.shareout());
defparam \Add2~9 .extended_lut = "off";
defparam \Add2~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add2~9 .shared_arith = "off";

arriaii_lcell_comb \Add2~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\rd_addr_2x[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~13_sumout ),
	.cout(\Add2~14 ),
	.shareout());
defparam \Add2~13 .extended_lut = "off";
defparam \Add2~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add2~13 .shared_arith = "off";

arriaii_lcell_comb \Add2~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\rd_addr_2x[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~17_sumout ),
	.cout(),
	.shareout());
defparam \Add2~17 .extended_lut = "off";
defparam \Add2~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add2~17 .shared_arith = "off";

dffeas bit_order_1x(
	.clk(clk_0),
	.d(\bit_order_1x~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\bit_order_1x~q ),
	.prn(vcc));
defparam bit_order_1x.is_wysiwyg = "true";
defparam bit_order_1x.power_up = "low";

dffeas ctl_doing_rd_beat2_1x_r1(
	.clk(clk_0),
	.d(ctl_doing_rd_beat2_1x),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctl_doing_rd_beat2_1x_r1~q ),
	.prn(vcc));
defparam ctl_doing_rd_beat2_1x_r1.is_wysiwyg = "true";
defparam ctl_doing_rd_beat2_1x_r1.power_up = "low";

arriaii_lcell_comb \wr_data_1x[0]~0 (
	.dataa(!seq_rdv_doing_rd_7),
	.datab(!merged_doing_rd),
	.datac(!\bit_order_1x~q ),
	.datad(!seq_poa_protection_override_1x),
	.datae(!\ctl_doing_rd_beat2_1x_r1~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wr_data_1x[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wr_data_1x[0]~0 .extended_lut = "off";
defparam \wr_data_1x[0]~0 .lut_mask = 64'h70FF7FFF70FF7FFF;
defparam \wr_data_1x[0]~0 .shared_arith = "off";

arriaii_lcell_comb \wr_data_1x[1]~1 (
	.dataa(!seq_rdv_doing_rd_7),
	.datab(!merged_doing_rd),
	.datac(!seq_rdv_doing_rd_4),
	.datad(!\bit_order_1x~q ),
	.datae(!seq_poa_protection_override_1x),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wr_data_1x[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wr_data_1x[1]~1 .extended_lut = "off";
defparam \wr_data_1x[1]~1 .lut_mask = 64'h3F77FFFF3F77FFFF;
defparam \wr_data_1x[1]~1 .shared_arith = "off";

dffeas \wr_addr_1x[0] (
	.clk(clk_0),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_addr_1x[0]~0_combout ),
	.q(\wr_addr_1x[0]~q ),
	.prn(vcc));
defparam \wr_addr_1x[0] .is_wysiwyg = "true";
defparam \wr_addr_1x[0] .power_up = "low";

dffeas \wr_addr_1x[1] (
	.clk(clk_0),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_addr_1x[0]~0_combout ),
	.q(\wr_addr_1x[1]~q ),
	.prn(vcc));
defparam \wr_addr_1x[1] .is_wysiwyg = "true";
defparam \wr_addr_1x[1] .power_up = "low";

dffeas \wr_addr_1x[2] (
	.clk(clk_0),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_addr_1x[0]~0_combout ),
	.q(\wr_addr_1x[2]~q ),
	.prn(vcc));
defparam \wr_addr_1x[2] .is_wysiwyg = "true";
defparam \wr_addr_1x[2] .power_up = "low";

dffeas \wr_addr_1x[3] (
	.clk(clk_0),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_addr_1x[0]~0_combout ),
	.q(\wr_addr_1x[3]~q ),
	.prn(vcc));
defparam \wr_addr_1x[3] .is_wysiwyg = "true";
defparam \wr_addr_1x[3] .power_up = "low";

dffeas \wr_addr_1x[4] (
	.clk(clk_0),
	.d(\wr_addr_1x[4]~1_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_addr_1x[4]~q ),
	.prn(vcc));
defparam \wr_addr_1x[4] .is_wysiwyg = "true";
defparam \wr_addr_1x[4] .power_up = "low";

dffeas \rd_addr_2x[1] (
	.clk(clk_4),
	.d(\Add2~1_sumout ),
	.asdata(vcc),
	.clrn(reset_poa_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_addr_2x[1]~q ),
	.prn(vcc));
defparam \rd_addr_2x[1] .is_wysiwyg = "true";
defparam \rd_addr_2x[1] .power_up = "low";

dffeas \rd_addr_2x[2] (
	.clk(clk_4),
	.d(\Add2~5_sumout ),
	.asdata(vcc),
	.clrn(reset_poa_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_addr_2x[2]~q ),
	.prn(vcc));
defparam \rd_addr_2x[2] .is_wysiwyg = "true";
defparam \rd_addr_2x[2] .power_up = "low";

dffeas \rd_addr_2x[3] (
	.clk(clk_4),
	.d(\Add2~9_sumout ),
	.asdata(vcc),
	.clrn(reset_poa_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_addr_2x[3]~q ),
	.prn(vcc));
defparam \rd_addr_2x[3] .is_wysiwyg = "true";
defparam \rd_addr_2x[3] .power_up = "low";

dffeas \rd_addr_2x[4] (
	.clk(clk_4),
	.d(\Add2~13_sumout ),
	.asdata(vcc),
	.clrn(reset_poa_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_addr_2x[4]~q ),
	.prn(vcc));
defparam \rd_addr_2x[4] .is_wysiwyg = "true";
defparam \rd_addr_2x[4] .power_up = "low";

dffeas \rd_addr_2x[5] (
	.clk(clk_4),
	.d(\Add2~17_sumout ),
	.asdata(vcc),
	.clrn(reset_poa_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_addr_2x[5]~q ),
	.prn(vcc));
defparam \rd_addr_2x[5] .is_wysiwyg = "true";
defparam \rd_addr_2x[5] .power_up = "low";

dffeas seq_poa_lat_dec_1x_1t(
	.clk(clk_0),
	.d(seq_poa_lat_dec_1x),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_poa_lat_dec_1x_1t~q ),
	.prn(vcc));
defparam seq_poa_lat_dec_1x_1t.is_wysiwyg = "true";
defparam seq_poa_lat_dec_1x_1t.power_up = "low";

arriaii_lcell_comb \bit_order_1x~0 (
	.dataa(!\bit_order_1x~q ),
	.datab(!\seq_poa_lat_dec_1x_1t~q ),
	.datac(!seq_poa_lat_dec_1x),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bit_order_1x~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bit_order_1x~0 .extended_lut = "off";
defparam \bit_order_1x~0 .lut_mask = 64'h5959595959595959;
defparam \bit_order_1x~0 .shared_arith = "off";

arriaii_lcell_comb \wr_addr_1x[0]~0 (
	.dataa(!\bit_order_1x~q ),
	.datab(!\seq_poa_lat_dec_1x_1t~q ),
	.datac(!seq_poa_lat_dec_1x),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wr_addr_1x[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wr_addr_1x[0]~0 .extended_lut = "off";
defparam \wr_addr_1x[0]~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \wr_addr_1x[0]~0 .shared_arith = "off";

arriaii_lcell_comb \wr_addr_1x[4]~1 (
	.dataa(!\wr_addr_1x[4]~q ),
	.datab(!\wr_addr_1x[0]~0_combout ),
	.datac(!\Add0~17_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wr_addr_1x[4]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wr_addr_1x[4]~1 .extended_lut = "off";
defparam \wr_addr_1x[4]~1 .lut_mask = 64'h7474747474747474;
defparam \wr_addr_1x[4]~1 .shared_arith = "off";

arriaii_lcell_comb \wr_addr_1x[4]~_wirecell (
	.dataa(!\wr_addr_1x[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wr_addr_1x[4]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wr_addr_1x[4]~_wirecell .extended_lut = "off";
defparam \wr_addr_1x[4]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \wr_addr_1x[4]~_wirecell .shared_arith = "off";

dffeas \rd_addr_2x[0] (
	.clk(clk_4),
	.d(\rd_addr_2x[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_poa_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rd_addr_2x_0),
	.prn(vcc));
defparam \rd_addr_2x[0] .is_wysiwyg = "true";
defparam \rd_addr_2x[0] .power_up = "low";

dffeas \postamble_en_pos_2x[0] (
	.clk(clk_4),
	.d(\postamble_en_2x_r[0]~q ),
	.asdata(vcc),
	.clrn(reset_poa_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(postamble_en_pos_2x_0),
	.prn(vcc));
defparam \postamble_en_pos_2x[0] .is_wysiwyg = "true";
defparam \postamble_en_pos_2x[0] .power_up = "low";

dffeas \postamble_en_pos_2x[1] (
	.clk(clk_4),
	.d(\postamble_en_2x_r[1]~q ),
	.asdata(vcc),
	.clrn(reset_poa_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(postamble_en_pos_2x_1),
	.prn(vcc));
defparam \postamble_en_pos_2x[1] .is_wysiwyg = "true";
defparam \postamble_en_pos_2x[1] .power_up = "low";

dffeas \postamble_en_pos_2x[2] (
	.clk(clk_4),
	.d(\postamble_en_2x_r[2]~q ),
	.asdata(vcc),
	.clrn(reset_poa_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(postamble_en_pos_2x_2),
	.prn(vcc));
defparam \postamble_en_pos_2x[2] .is_wysiwyg = "true";
defparam \postamble_en_pos_2x[2] .power_up = "low";

dffeas \postamble_en_pos_2x[3] (
	.clk(clk_4),
	.d(\postamble_en_2x_r[3]~q ),
	.asdata(vcc),
	.clrn(reset_poa_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(postamble_en_pos_2x_3),
	.prn(vcc));
defparam \postamble_en_pos_2x[3] .is_wysiwyg = "true";
defparam \postamble_en_pos_2x[3] .power_up = "low";

arriaii_lcell_comb \rd_addr_2x[0]~0 (
	.dataa(!rd_addr_2x_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rd_addr_2x[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_addr_2x[0]~0 .extended_lut = "off";
defparam \rd_addr_2x[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rd_addr_2x[0]~0 .shared_arith = "off";

dffeas \postamble_en_2x_r[0] (
	.clk(clk_4),
	.d(\half_rate_ram_gen.altsyncram_inst|auto_generated|q_b[0] ),
	.asdata(vcc),
	.clrn(reset_poa_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\postamble_en_2x_r[0]~q ),
	.prn(vcc));
defparam \postamble_en_2x_r[0] .is_wysiwyg = "true";
defparam \postamble_en_2x_r[0] .power_up = "low";

dffeas \postamble_en_2x_r[1] (
	.clk(clk_4),
	.d(\half_rate_ram_gen.altsyncram_inst|auto_generated|q_b[0] ),
	.asdata(vcc),
	.clrn(reset_poa_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\postamble_en_2x_r[1]~q ),
	.prn(vcc));
defparam \postamble_en_2x_r[1] .is_wysiwyg = "true";
defparam \postamble_en_2x_r[1] .power_up = "low";

dffeas \postamble_en_2x_r[2] (
	.clk(clk_4),
	.d(\half_rate_ram_gen.altsyncram_inst|auto_generated|q_b[0] ),
	.asdata(vcc),
	.clrn(reset_poa_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\postamble_en_2x_r[2]~q ),
	.prn(vcc));
defparam \postamble_en_2x_r[2] .is_wysiwyg = "true";
defparam \postamble_en_2x_r[2] .power_up = "low";

dffeas \postamble_en_2x_r[3] (
	.clk(clk_4),
	.d(\half_rate_ram_gen.altsyncram_inst|auto_generated|q_b[0] ),
	.asdata(vcc),
	.clrn(reset_poa_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\postamble_en_2x_r[3]~q ),
	.prn(vcc));
defparam \postamble_en_2x_r[3] .is_wysiwyg = "true";
defparam \postamble_en_2x_r[3] .power_up = "low";

endmodule

module ddr3_int_altsyncram_1 (
	clock0,
	clock1,
	q_b,
	address_b,
	data_a,
	address_a)/* synthesis synthesis_greybox=0 */;
input 	clock0;
input 	clock1;
output 	[127:0] q_b;
input 	[5:0] address_b;
input 	[63:0] data_a;
input 	[4:0] address_a;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_altsyncram_78h1 auto_generated(
	.clock0(clock0),
	.clock1(clock1),
	.q_b({q_b[0]}),
	.address_b({address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.data_a({data_a[1],data_a[0]}),
	.address_a({address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}));

endmodule

module ddr3_int_altsyncram_78h1 (
	clock0,
	clock1,
	q_b,
	address_b,
	data_a,
	address_a)/* synthesis synthesis_greybox=0 */;
input 	clock0;
input 	clock1;
output 	[0:0] q_b;
input 	[5:0] address_b;
input 	[1:0] data_a;
input 	[4:0] address_a;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

arriaii_ram_block ram_block1a0(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1],data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena2";
defparam ram_block1a0.clk1_core_clock_enable = "ena3";
defparam ram_block1a0.clk1_input_clock_enable = "ena3";
defparam ram_block1a0.clock_duty_cycle_dependence = "on";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_postamble:poa|altsyncram:half_rate_ram_gen.altsyncram_inst|altsyncram_78h1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 5;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 2;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 31;
defparam ram_block1a0.port_a_logical_ram_depth = 32;
defparam ram_block1a0.port_a_logical_ram_width = 2;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 6;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock1";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 63;
defparam ram_block1a0.port_b_logical_ram_depth = 64;
defparam ram_block1a0.port_b_logical_ram_width = 1;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_rdata_valid (
	clk_0,
	do_read_r,
	ctl_rdata_valid_0,
	ctl_init_success,
	rd_addr_0,
	reset_phy_clk_1x_n,
	rdwr_data_valid_r,
	seq_rdv_doing_rd_7,
	doing_read,
	merged_doing_rd,
	seq_rdata_valid_lat_dec,
	seq_rdv_doing_rd_4,
	seq_rdata_valid_0,
	seq_rdata_valid_1)/* synthesis synthesis_greybox=0 */;
input 	clk_0;
input 	do_read_r;
output 	ctl_rdata_valid_0;
input 	ctl_init_success;
output 	rd_addr_0;
input 	reset_phy_clk_1x_n;
input 	rdwr_data_valid_r;
input 	seq_rdv_doing_rd_7;
input 	doing_read;
output 	merged_doing_rd;
input 	seq_rdata_valid_lat_dec;
input 	seq_rdv_doing_rd_4;
output 	seq_rdata_valid_0;
output 	seq_rdata_valid_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altsyncram_component|auto_generated|q_b[0] ;
wire \Add0~1_sumout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \Add2~1_sumout ;
wire \Add2~2 ;
wire \Add2~5_sumout ;
wire \Add2~6 ;
wire \Add2~9_sumout ;
wire \Add2~10 ;
wire \Add2~13_sumout ;
wire \altsyncram_component|auto_generated|q_b[1] ;
wire \bit_order_1x~q ;
wire \rdv_pipe_ip_beat2_r~q ;
wire \wr_data[0]~0_combout ;
wire \wr_addr[0]~q ;
wire \wr_addr[1]~q ;
wire \wr_addr[2]~q ;
wire \wr_addr[3]~q ;
wire \wr_addr[4]~q ;
wire \rd_addr[1]~q ;
wire \rd_addr[2]~q ;
wire \rd_addr[3]~q ;
wire \rd_addr[4]~q ;
wire \seq_rdata_valid_lat_dec_1t~q ;
wire \bit_order_1x~0_combout ;
wire \WideOr1~combout ;
wire \wr_addr[0]~0_combout ;
wire \wr_addr[3]~1_combout ;
wire \wr_data[1]~1_combout ;
wire \wr_addr[0]~2_combout ;
wire \wr_addr[1]~3_combout ;
wire \wr_addr[2]~4_combout ;
wire \wr_addr[4]~5_combout ;
wire \wr_addr[0]~_wirecell_combout ;
wire \wr_addr[1]~_wirecell_combout ;
wire \wr_addr[2]~_wirecell_combout ;
wire \wr_addr[4]~_wirecell_combout ;
wire \ctl_rdata_valid~0_combout ;
wire \rd_addr[0]~0_combout ;


ddr3_int_altsyncram_2 altsyncram_component(
	.clock0(clk_0),
	.q_b({q_b_unconnected_wire_127,q_b_unconnected_wire_126,q_b_unconnected_wire_125,q_b_unconnected_wire_124,q_b_unconnected_wire_123,q_b_unconnected_wire_122,q_b_unconnected_wire_121,q_b_unconnected_wire_120,q_b_unconnected_wire_119,q_b_unconnected_wire_118,
q_b_unconnected_wire_117,q_b_unconnected_wire_116,q_b_unconnected_wire_115,q_b_unconnected_wire_114,q_b_unconnected_wire_113,q_b_unconnected_wire_112,q_b_unconnected_wire_111,q_b_unconnected_wire_110,q_b_unconnected_wire_109,q_b_unconnected_wire_108,
q_b_unconnected_wire_107,q_b_unconnected_wire_106,q_b_unconnected_wire_105,q_b_unconnected_wire_104,q_b_unconnected_wire_103,q_b_unconnected_wire_102,q_b_unconnected_wire_101,q_b_unconnected_wire_100,q_b_unconnected_wire_99,q_b_unconnected_wire_98,
q_b_unconnected_wire_97,q_b_unconnected_wire_96,q_b_unconnected_wire_95,q_b_unconnected_wire_94,q_b_unconnected_wire_93,q_b_unconnected_wire_92,q_b_unconnected_wire_91,q_b_unconnected_wire_90,q_b_unconnected_wire_89,q_b_unconnected_wire_88,q_b_unconnected_wire_87,
q_b_unconnected_wire_86,q_b_unconnected_wire_85,q_b_unconnected_wire_84,q_b_unconnected_wire_83,q_b_unconnected_wire_82,q_b_unconnected_wire_81,q_b_unconnected_wire_80,q_b_unconnected_wire_79,q_b_unconnected_wire_78,q_b_unconnected_wire_77,q_b_unconnected_wire_76,
q_b_unconnected_wire_75,q_b_unconnected_wire_74,q_b_unconnected_wire_73,q_b_unconnected_wire_72,q_b_unconnected_wire_71,q_b_unconnected_wire_70,q_b_unconnected_wire_69,q_b_unconnected_wire_68,q_b_unconnected_wire_67,q_b_unconnected_wire_66,q_b_unconnected_wire_65,
q_b_unconnected_wire_64,q_b_unconnected_wire_63,q_b_unconnected_wire_62,q_b_unconnected_wire_61,q_b_unconnected_wire_60,q_b_unconnected_wire_59,q_b_unconnected_wire_58,q_b_unconnected_wire_57,q_b_unconnected_wire_56,q_b_unconnected_wire_55,q_b_unconnected_wire_54,
q_b_unconnected_wire_53,q_b_unconnected_wire_52,q_b_unconnected_wire_51,q_b_unconnected_wire_50,q_b_unconnected_wire_49,q_b_unconnected_wire_48,q_b_unconnected_wire_47,q_b_unconnected_wire_46,q_b_unconnected_wire_45,q_b_unconnected_wire_44,q_b_unconnected_wire_43,
q_b_unconnected_wire_42,q_b_unconnected_wire_41,q_b_unconnected_wire_40,q_b_unconnected_wire_39,q_b_unconnected_wire_38,q_b_unconnected_wire_37,q_b_unconnected_wire_36,q_b_unconnected_wire_35,q_b_unconnected_wire_34,q_b_unconnected_wire_33,q_b_unconnected_wire_32,
q_b_unconnected_wire_31,q_b_unconnected_wire_30,q_b_unconnected_wire_29,q_b_unconnected_wire_28,q_b_unconnected_wire_27,q_b_unconnected_wire_26,q_b_unconnected_wire_25,q_b_unconnected_wire_24,q_b_unconnected_wire_23,q_b_unconnected_wire_22,q_b_unconnected_wire_21,
q_b_unconnected_wire_20,q_b_unconnected_wire_19,q_b_unconnected_wire_18,q_b_unconnected_wire_17,q_b_unconnected_wire_16,q_b_unconnected_wire_15,q_b_unconnected_wire_14,q_b_unconnected_wire_13,q_b_unconnected_wire_12,q_b_unconnected_wire_11,q_b_unconnected_wire_10,
q_b_unconnected_wire_9,q_b_unconnected_wire_8,q_b_unconnected_wire_7,q_b_unconnected_wire_6,q_b_unconnected_wire_5,q_b_unconnected_wire_4,q_b_unconnected_wire_3,q_b_unconnected_wire_2,\altsyncram_component|auto_generated|q_b[1] ,
\altsyncram_component|auto_generated|q_b[0] }),
	.address_b({gnd,\rd_addr[4]~q ,\rd_addr[3]~q ,\rd_addr[2]~q ,\rd_addr[1]~q ,rd_addr_0}),
	.data_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_data[1]~1_combout ,\wr_data[0]~0_combout }),
	.address_a({\wr_addr[4]~_wirecell_combout ,\wr_addr[3]~q ,\wr_addr[2]~_wirecell_combout ,\wr_addr[1]~_wirecell_combout ,\wr_addr[0]~_wirecell_combout }));

arriaii_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\wr_addr[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "off";

arriaii_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\wr_addr[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FFFF0000FF00;
defparam \Add0~5 .shared_arith = "off";

arriaii_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\wr_addr[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FFFF0000FF00;
defparam \Add0~9 .shared_arith = "off";

arriaii_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\wr_addr[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~13 .shared_arith = "off";

arriaii_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\wr_addr[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FFFF0000FF00;
defparam \Add0~17 .shared_arith = "off";

arriaii_lcell_comb \Add2~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!rd_addr_0),
	.datae(gnd),
	.dataf(!\rd_addr[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~1_sumout ),
	.cout(\Add2~2 ),
	.shareout());
defparam \Add2~1 .extended_lut = "off";
defparam \Add2~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add2~1 .shared_arith = "off";

arriaii_lcell_comb \Add2~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\rd_addr[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~5_sumout ),
	.cout(\Add2~6 ),
	.shareout());
defparam \Add2~5 .extended_lut = "off";
defparam \Add2~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add2~5 .shared_arith = "off";

arriaii_lcell_comb \Add2~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\rd_addr[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~9_sumout ),
	.cout(\Add2~10 ),
	.shareout());
defparam \Add2~9 .extended_lut = "off";
defparam \Add2~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add2~9 .shared_arith = "off";

arriaii_lcell_comb \Add2~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\rd_addr[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~13_sumout ),
	.cout(),
	.shareout());
defparam \Add2~13 .extended_lut = "off";
defparam \Add2~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add2~13 .shared_arith = "off";

dffeas bit_order_1x(
	.clk(clk_0),
	.d(\bit_order_1x~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\bit_order_1x~q ),
	.prn(vcc));
defparam bit_order_1x.is_wysiwyg = "true";
defparam bit_order_1x.power_up = "low";

dffeas rdv_pipe_ip_beat2_r(
	.clk(clk_0),
	.d(\WideOr1~combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(reset_phy_clk_1x_n),
	.q(\rdv_pipe_ip_beat2_r~q ),
	.prn(vcc));
defparam rdv_pipe_ip_beat2_r.is_wysiwyg = "true";
defparam rdv_pipe_ip_beat2_r.power_up = "low";

arriaii_lcell_comb \wr_data[0]~0 (
	.dataa(!\bit_order_1x~q ),
	.datab(!\rdv_pipe_ip_beat2_r~q ),
	.datac(!seq_rdv_doing_rd_7),
	.datad(!merged_doing_rd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wr_data[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wr_data[0]~0 .extended_lut = "off";
defparam \wr_data[0]~0 .lut_mask = 64'h2777277727772777;
defparam \wr_data[0]~0 .shared_arith = "off";

dffeas \wr_addr[0] (
	.clk(clk_0),
	.d(\wr_addr[0]~2_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_addr[0]~0_combout ),
	.q(\wr_addr[0]~q ),
	.prn(vcc));
defparam \wr_addr[0] .is_wysiwyg = "true";
defparam \wr_addr[0] .power_up = "low";

dffeas \wr_addr[1] (
	.clk(clk_0),
	.d(\wr_addr[1]~3_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_addr[0]~0_combout ),
	.q(\wr_addr[1]~q ),
	.prn(vcc));
defparam \wr_addr[1] .is_wysiwyg = "true";
defparam \wr_addr[1] .power_up = "low";

dffeas \wr_addr[2] (
	.clk(clk_0),
	.d(\wr_addr[2]~4_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_addr[0]~0_combout ),
	.q(\wr_addr[2]~q ),
	.prn(vcc));
defparam \wr_addr[2] .is_wysiwyg = "true";
defparam \wr_addr[2] .power_up = "low";

dffeas \wr_addr[3] (
	.clk(clk_0),
	.d(\wr_addr[3]~1_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_addr[3]~q ),
	.prn(vcc));
defparam \wr_addr[3] .is_wysiwyg = "true";
defparam \wr_addr[3] .power_up = "low";

dffeas \wr_addr[4] (
	.clk(clk_0),
	.d(\wr_addr[4]~5_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wr_addr[0]~0_combout ),
	.q(\wr_addr[4]~q ),
	.prn(vcc));
defparam \wr_addr[4] .is_wysiwyg = "true";
defparam \wr_addr[4] .power_up = "low";

dffeas \rd_addr[1] (
	.clk(clk_0),
	.d(\Add2~1_sumout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_addr[1]~q ),
	.prn(vcc));
defparam \rd_addr[1] .is_wysiwyg = "true";
defparam \rd_addr[1] .power_up = "low";

dffeas \rd_addr[2] (
	.clk(clk_0),
	.d(\Add2~5_sumout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_addr[2]~q ),
	.prn(vcc));
defparam \rd_addr[2] .is_wysiwyg = "true";
defparam \rd_addr[2] .power_up = "low";

dffeas \rd_addr[3] (
	.clk(clk_0),
	.d(\Add2~9_sumout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_addr[3]~q ),
	.prn(vcc));
defparam \rd_addr[3] .is_wysiwyg = "true";
defparam \rd_addr[3] .power_up = "low";

dffeas \rd_addr[4] (
	.clk(clk_0),
	.d(\Add2~13_sumout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_addr[4]~q ),
	.prn(vcc));
defparam \rd_addr[4] .is_wysiwyg = "true";
defparam \rd_addr[4] .power_up = "low";

dffeas seq_rdata_valid_lat_dec_1t(
	.clk(clk_0),
	.d(seq_rdata_valid_lat_dec),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_rdata_valid_lat_dec_1t~q ),
	.prn(vcc));
defparam seq_rdata_valid_lat_dec_1t.is_wysiwyg = "true";
defparam seq_rdata_valid_lat_dec_1t.power_up = "low";

arriaii_lcell_comb \bit_order_1x~0 (
	.dataa(!\bit_order_1x~q ),
	.datab(!seq_rdata_valid_lat_dec),
	.datac(!\seq_rdata_valid_lat_dec_1t~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\bit_order_1x~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \bit_order_1x~0 .extended_lut = "off";
defparam \bit_order_1x~0 .lut_mask = 64'h6565656565656565;
defparam \bit_order_1x~0 .shared_arith = "off";

arriaii_lcell_comb WideOr1(
	.dataa(!seq_rdv_doing_rd_7),
	.datab(!merged_doing_rd),
	.datac(!seq_rdv_doing_rd_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam WideOr1.shared_arith = "off";

arriaii_lcell_comb \wr_addr[0]~0 (
	.dataa(!\bit_order_1x~q ),
	.datab(!seq_rdata_valid_lat_dec),
	.datac(!\seq_rdata_valid_lat_dec_1t~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wr_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wr_addr[0]~0 .extended_lut = "off";
defparam \wr_addr[0]~0 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \wr_addr[0]~0 .shared_arith = "off";

arriaii_lcell_comb \wr_addr[3]~1 (
	.dataa(!\wr_addr[3]~q ),
	.datab(!\wr_addr[0]~0_combout ),
	.datac(!\Add0~13_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wr_addr[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wr_addr[3]~1 .extended_lut = "off";
defparam \wr_addr[3]~1 .lut_mask = 64'h4747474747474747;
defparam \wr_addr[3]~1 .shared_arith = "off";

arriaii_lcell_comb \wr_data[1]~1 (
	.dataa(!\bit_order_1x~q ),
	.datab(!seq_rdv_doing_rd_7),
	.datac(!merged_doing_rd),
	.datad(!seq_rdv_doing_rd_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wr_data[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wr_data[1]~1 .extended_lut = "off";
defparam \wr_data[1]~1 .lut_mask = 64'h3F7F3F7F3F7F3F7F;
defparam \wr_data[1]~1 .shared_arith = "off";

arriaii_lcell_comb \wr_addr[0]~2 (
	.dataa(!\Add0~1_sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wr_addr[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wr_addr[0]~2 .extended_lut = "off";
defparam \wr_addr[0]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \wr_addr[0]~2 .shared_arith = "off";

arriaii_lcell_comb \wr_addr[1]~3 (
	.dataa(!\Add0~5_sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wr_addr[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wr_addr[1]~3 .extended_lut = "off";
defparam \wr_addr[1]~3 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \wr_addr[1]~3 .shared_arith = "off";

arriaii_lcell_comb \wr_addr[2]~4 (
	.dataa(!\Add0~9_sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wr_addr[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wr_addr[2]~4 .extended_lut = "off";
defparam \wr_addr[2]~4 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \wr_addr[2]~4 .shared_arith = "off";

arriaii_lcell_comb \wr_addr[4]~5 (
	.dataa(!\Add0~17_sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wr_addr[4]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wr_addr[4]~5 .extended_lut = "off";
defparam \wr_addr[4]~5 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \wr_addr[4]~5 .shared_arith = "off";

arriaii_lcell_comb \wr_addr[0]~_wirecell (
	.dataa(!\wr_addr[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wr_addr[0]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wr_addr[0]~_wirecell .extended_lut = "off";
defparam \wr_addr[0]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \wr_addr[0]~_wirecell .shared_arith = "off";

arriaii_lcell_comb \wr_addr[1]~_wirecell (
	.dataa(!\wr_addr[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wr_addr[1]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wr_addr[1]~_wirecell .extended_lut = "off";
defparam \wr_addr[1]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \wr_addr[1]~_wirecell .shared_arith = "off";

arriaii_lcell_comb \wr_addr[2]~_wirecell (
	.dataa(!\wr_addr[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wr_addr[2]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wr_addr[2]~_wirecell .extended_lut = "off";
defparam \wr_addr[2]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \wr_addr[2]~_wirecell .shared_arith = "off";

arriaii_lcell_comb \wr_addr[4]~_wirecell (
	.dataa(!\wr_addr[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wr_addr[4]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wr_addr[4]~_wirecell .extended_lut = "off";
defparam \wr_addr[4]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \wr_addr[4]~_wirecell .shared_arith = "off";

dffeas \ctl_rdata_valid[0] (
	.clk(clk_0),
	.d(\ctl_rdata_valid~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ctl_rdata_valid_0),
	.prn(vcc));
defparam \ctl_rdata_valid[0] .is_wysiwyg = "true";
defparam \ctl_rdata_valid[0] .power_up = "low";

dffeas \rd_addr[0] (
	.clk(clk_0),
	.d(\rd_addr[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rd_addr_0),
	.prn(vcc));
defparam \rd_addr[0] .is_wysiwyg = "true";
defparam \rd_addr[0] .power_up = "low";

arriaii_lcell_comb \merged_doing_rd~0 (
	.dataa(!ctl_init_success),
	.datab(!do_read_r),
	.datac(!rdwr_data_valid_r),
	.datad(!doing_read),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(merged_doing_rd),
	.sumout(),
	.cout(),
	.shareout());
defparam \merged_doing_rd~0 .extended_lut = "off";
defparam \merged_doing_rd~0 .lut_mask = 64'h0105010501050105;
defparam \merged_doing_rd~0 .shared_arith = "off";

dffeas \seq_rdata_valid[0] (
	.clk(clk_0),
	.d(\altsyncram_component|auto_generated|q_b[0] ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_rdata_valid_0),
	.prn(vcc));
defparam \seq_rdata_valid[0] .is_wysiwyg = "true";
defparam \seq_rdata_valid[0] .power_up = "low";

dffeas \seq_rdata_valid[1] (
	.clk(clk_0),
	.d(\altsyncram_component|auto_generated|q_b[1] ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_rdata_valid_1),
	.prn(vcc));
defparam \seq_rdata_valid[1] .is_wysiwyg = "true";
defparam \seq_rdata_valid[1] .power_up = "low";

arriaii_lcell_comb \ctl_rdata_valid~0 (
	.dataa(!ctl_init_success),
	.datab(!\altsyncram_component|auto_generated|q_b[0] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ctl_rdata_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctl_rdata_valid~0 .extended_lut = "off";
defparam \ctl_rdata_valid~0 .lut_mask = 64'h1111111111111111;
defparam \ctl_rdata_valid~0 .shared_arith = "off";

arriaii_lcell_comb \rd_addr[0]~0 (
	.dataa(!rd_addr_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rd_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_addr[0]~0 .extended_lut = "off";
defparam \rd_addr[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rd_addr[0]~0 .shared_arith = "off";

endmodule

module ddr3_int_altsyncram_2 (
	clock0,
	q_b,
	address_b,
	data_a,
	address_a)/* synthesis synthesis_greybox=0 */;
input 	clock0;
output 	[127:0] q_b;
input 	[5:0] address_b;
input 	[63:0] data_a;
input 	[4:0] address_a;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_altsyncram_ski1 auto_generated(
	.clock0(clock0),
	.q_b({q_b[1],q_b[0]}),
	.address_b({address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.data_a({data_a[1],data_a[0]}),
	.address_a({address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}));

endmodule

module ddr3_int_altsyncram_ski1 (
	clock0,
	q_b,
	address_b,
	data_a,
	address_a)/* synthesis synthesis_greybox=0 */;
input 	clock0;
output 	[1:0] q_b;
input 	[4:0] address_b;
input 	[1:0] data_a;
input 	[4:0] address_a;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

arriaii_ram_block ram_block1a0(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena2";
defparam ram_block1a0.clk0_input_clock_enable = "ena2";
defparam ram_block1a0.clock_duty_cycle_dependence = "on";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_rdata_valid:rdv_pipe|altsyncram:altsyncram_component|altsyncram_ski1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 5;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 31;
defparam ram_block1a0.port_a_logical_ram_depth = 32;
defparam ram_block1a0.port_a_logical_ram_width = 2;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 5;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 31;
defparam ram_block1a0.port_b_logical_ram_depth = 32;
defparam ram_block1a0.port_b_logical_ram_width = 2;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

arriaii_ram_block ram_block1a1(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena2";
defparam ram_block1a1.clk0_input_clock_enable = "ena2";
defparam ram_block1a1.clock_duty_cycle_dependence = "on";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_rdata_valid:rdv_pipe|altsyncram:altsyncram_component|altsyncram_ski1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 5;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 31;
defparam ram_block1a1.port_a_logical_ram_depth = 32;
defparam ram_block1a1.port_a_logical_ram_width = 2;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 5;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 31;
defparam ram_block1a1.port_b_logical_ram_depth = 32;
defparam ram_block1a1.port_b_logical_ram_width = 2;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_read_dp (
	q_b_0,
	q_b_64,
	q_b_1,
	q_b_65,
	q_b_2,
	q_b_66,
	q_b_3,
	q_b_67,
	q_b_4,
	q_b_68,
	q_b_5,
	q_b_69,
	q_b_6,
	q_b_70,
	q_b_7,
	q_b_71,
	q_b_16,
	q_b_80,
	q_b_17,
	q_b_81,
	q_b_18,
	q_b_82,
	q_b_19,
	q_b_83,
	q_b_20,
	q_b_84,
	q_b_21,
	q_b_85,
	q_b_22,
	q_b_86,
	q_b_23,
	q_b_87,
	q_b_32,
	q_b_96,
	q_b_33,
	q_b_97,
	q_b_34,
	q_b_98,
	q_b_35,
	q_b_99,
	q_b_36,
	q_b_100,
	q_b_37,
	q_b_101,
	q_b_38,
	q_b_102,
	q_b_39,
	q_b_103,
	q_b_48,
	q_b_112,
	q_b_49,
	q_b_113,
	q_b_50,
	q_b_114,
	q_b_51,
	q_b_115,
	q_b_52,
	q_b_116,
	q_b_53,
	q_b_117,
	q_b_54,
	q_b_118,
	q_b_55,
	q_b_119,
	q_b_8,
	q_b_72,
	q_b_9,
	q_b_73,
	q_b_10,
	q_b_74,
	q_b_11,
	q_b_75,
	q_b_12,
	q_b_76,
	q_b_13,
	q_b_77,
	q_b_14,
	q_b_78,
	q_b_15,
	q_b_79,
	q_b_24,
	q_b_88,
	q_b_25,
	q_b_89,
	q_b_26,
	q_b_90,
	q_b_27,
	q_b_91,
	q_b_28,
	q_b_92,
	q_b_29,
	q_b_93,
	q_b_30,
	q_b_94,
	q_b_31,
	q_b_95,
	q_b_40,
	q_b_104,
	q_b_41,
	q_b_105,
	q_b_42,
	q_b_106,
	q_b_43,
	q_b_107,
	q_b_44,
	q_b_108,
	q_b_45,
	q_b_109,
	q_b_46,
	q_b_110,
	q_b_47,
	q_b_111,
	q_b_56,
	q_b_120,
	q_b_57,
	q_b_121,
	q_b_58,
	q_b_122,
	q_b_59,
	q_b_123,
	q_b_60,
	q_b_124,
	q_b_61,
	q_b_125,
	q_b_62,
	q_b_126,
	q_b_63,
	q_b_127,
	clk_0,
	clk_4,
	dio_rdata_h_2x_0,
	rd_addr_2x_0,
	rd_addr_0,
	dio_rdata_h_2x_1,
	dio_rdata_h_2x_2,
	dio_rdata_h_2x_3,
	dio_rdata_h_2x_4,
	dio_rdata_h_2x_5,
	dio_rdata_h_2x_6,
	dio_rdata_h_2x_7,
	dio_rdata_h_2x_8,
	dio_rdata_h_2x_9,
	dio_rdata_h_2x_10,
	dio_rdata_h_2x_11,
	dio_rdata_h_2x_12,
	dio_rdata_h_2x_13,
	dio_rdata_h_2x_14,
	dio_rdata_h_2x_15,
	dio_rdata_h_2x_16,
	dio_rdata_h_2x_17,
	dio_rdata_h_2x_18,
	dio_rdata_h_2x_19,
	dio_rdata_h_2x_20,
	dio_rdata_h_2x_21,
	dio_rdata_h_2x_22,
	dio_rdata_h_2x_23,
	dio_rdata_h_2x_24,
	dio_rdata_h_2x_25,
	dio_rdata_h_2x_26,
	dio_rdata_h_2x_27,
	dio_rdata_h_2x_28,
	dio_rdata_h_2x_29,
	dio_rdata_h_2x_30,
	dio_rdata_h_2x_31,
	dio_rdata_l_2x_0,
	dio_rdata_l_2x_1,
	dio_rdata_l_2x_2,
	dio_rdata_l_2x_3,
	dio_rdata_l_2x_4,
	dio_rdata_l_2x_5,
	dio_rdata_l_2x_6,
	dio_rdata_l_2x_7,
	dio_rdata_l_2x_8,
	dio_rdata_l_2x_9,
	dio_rdata_l_2x_10,
	dio_rdata_l_2x_11,
	dio_rdata_l_2x_12,
	dio_rdata_l_2x_13,
	dio_rdata_l_2x_14,
	dio_rdata_l_2x_15,
	dio_rdata_l_2x_16,
	dio_rdata_l_2x_17,
	dio_rdata_l_2x_18,
	dio_rdata_l_2x_19,
	dio_rdata_l_2x_20,
	dio_rdata_l_2x_21,
	dio_rdata_l_2x_22,
	dio_rdata_l_2x_23,
	dio_rdata_l_2x_24,
	dio_rdata_l_2x_25,
	dio_rdata_l_2x_26,
	dio_rdata_l_2x_27,
	dio_rdata_l_2x_28,
	dio_rdata_l_2x_29,
	dio_rdata_l_2x_30,
	dio_rdata_l_2x_31,
	reset_phy_clk_1x_n,
	reset_resync_clk_2x_n)/* synthesis synthesis_greybox=0 */;
output 	q_b_0;
output 	q_b_64;
output 	q_b_1;
output 	q_b_65;
output 	q_b_2;
output 	q_b_66;
output 	q_b_3;
output 	q_b_67;
output 	q_b_4;
output 	q_b_68;
output 	q_b_5;
output 	q_b_69;
output 	q_b_6;
output 	q_b_70;
output 	q_b_7;
output 	q_b_71;
output 	q_b_16;
output 	q_b_80;
output 	q_b_17;
output 	q_b_81;
output 	q_b_18;
output 	q_b_82;
output 	q_b_19;
output 	q_b_83;
output 	q_b_20;
output 	q_b_84;
output 	q_b_21;
output 	q_b_85;
output 	q_b_22;
output 	q_b_86;
output 	q_b_23;
output 	q_b_87;
output 	q_b_32;
output 	q_b_96;
output 	q_b_33;
output 	q_b_97;
output 	q_b_34;
output 	q_b_98;
output 	q_b_35;
output 	q_b_99;
output 	q_b_36;
output 	q_b_100;
output 	q_b_37;
output 	q_b_101;
output 	q_b_38;
output 	q_b_102;
output 	q_b_39;
output 	q_b_103;
output 	q_b_48;
output 	q_b_112;
output 	q_b_49;
output 	q_b_113;
output 	q_b_50;
output 	q_b_114;
output 	q_b_51;
output 	q_b_115;
output 	q_b_52;
output 	q_b_116;
output 	q_b_53;
output 	q_b_117;
output 	q_b_54;
output 	q_b_118;
output 	q_b_55;
output 	q_b_119;
output 	q_b_8;
output 	q_b_72;
output 	q_b_9;
output 	q_b_73;
output 	q_b_10;
output 	q_b_74;
output 	q_b_11;
output 	q_b_75;
output 	q_b_12;
output 	q_b_76;
output 	q_b_13;
output 	q_b_77;
output 	q_b_14;
output 	q_b_78;
output 	q_b_15;
output 	q_b_79;
output 	q_b_24;
output 	q_b_88;
output 	q_b_25;
output 	q_b_89;
output 	q_b_26;
output 	q_b_90;
output 	q_b_27;
output 	q_b_91;
output 	q_b_28;
output 	q_b_92;
output 	q_b_29;
output 	q_b_93;
output 	q_b_30;
output 	q_b_94;
output 	q_b_31;
output 	q_b_95;
output 	q_b_40;
output 	q_b_104;
output 	q_b_41;
output 	q_b_105;
output 	q_b_42;
output 	q_b_106;
output 	q_b_43;
output 	q_b_107;
output 	q_b_44;
output 	q_b_108;
output 	q_b_45;
output 	q_b_109;
output 	q_b_46;
output 	q_b_110;
output 	q_b_47;
output 	q_b_111;
output 	q_b_56;
output 	q_b_120;
output 	q_b_57;
output 	q_b_121;
output 	q_b_58;
output 	q_b_122;
output 	q_b_59;
output 	q_b_123;
output 	q_b_60;
output 	q_b_124;
output 	q_b_61;
output 	q_b_125;
output 	q_b_62;
output 	q_b_126;
output 	q_b_63;
output 	q_b_127;
input 	clk_0;
input 	clk_4;
input 	dio_rdata_h_2x_0;
input 	rd_addr_2x_0;
input 	rd_addr_0;
input 	dio_rdata_h_2x_1;
input 	dio_rdata_h_2x_2;
input 	dio_rdata_h_2x_3;
input 	dio_rdata_h_2x_4;
input 	dio_rdata_h_2x_5;
input 	dio_rdata_h_2x_6;
input 	dio_rdata_h_2x_7;
input 	dio_rdata_h_2x_8;
input 	dio_rdata_h_2x_9;
input 	dio_rdata_h_2x_10;
input 	dio_rdata_h_2x_11;
input 	dio_rdata_h_2x_12;
input 	dio_rdata_h_2x_13;
input 	dio_rdata_h_2x_14;
input 	dio_rdata_h_2x_15;
input 	dio_rdata_h_2x_16;
input 	dio_rdata_h_2x_17;
input 	dio_rdata_h_2x_18;
input 	dio_rdata_h_2x_19;
input 	dio_rdata_h_2x_20;
input 	dio_rdata_h_2x_21;
input 	dio_rdata_h_2x_22;
input 	dio_rdata_h_2x_23;
input 	dio_rdata_h_2x_24;
input 	dio_rdata_h_2x_25;
input 	dio_rdata_h_2x_26;
input 	dio_rdata_h_2x_27;
input 	dio_rdata_h_2x_28;
input 	dio_rdata_h_2x_29;
input 	dio_rdata_h_2x_30;
input 	dio_rdata_h_2x_31;
input 	dio_rdata_l_2x_0;
input 	dio_rdata_l_2x_1;
input 	dio_rdata_l_2x_2;
input 	dio_rdata_l_2x_3;
input 	dio_rdata_l_2x_4;
input 	dio_rdata_l_2x_5;
input 	dio_rdata_l_2x_6;
input 	dio_rdata_l_2x_7;
input 	dio_rdata_l_2x_8;
input 	dio_rdata_l_2x_9;
input 	dio_rdata_l_2x_10;
input 	dio_rdata_l_2x_11;
input 	dio_rdata_l_2x_12;
input 	dio_rdata_l_2x_13;
input 	dio_rdata_l_2x_14;
input 	dio_rdata_l_2x_15;
input 	dio_rdata_l_2x_16;
input 	dio_rdata_l_2x_17;
input 	dio_rdata_l_2x_18;
input 	dio_rdata_l_2x_19;
input 	dio_rdata_l_2x_20;
input 	dio_rdata_l_2x_21;
input 	dio_rdata_l_2x_22;
input 	dio_rdata_l_2x_23;
input 	dio_rdata_l_2x_24;
input 	dio_rdata_l_2x_25;
input 	dio_rdata_l_2x_26;
input 	dio_rdata_l_2x_27;
input 	dio_rdata_l_2x_28;
input 	dio_rdata_l_2x_29;
input 	dio_rdata_l_2x_30;
input 	dio_rdata_l_2x_31;
input 	reset_phy_clk_1x_n;
input 	reset_resync_clk_2x_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \rd_ram_wr_addr[1]~q ;
wire \rd_ram_wr_addr[2]~q ;
wire \rd_ram_wr_addr[3]~q ;
wire \rd_ram_rd_addr[1]~q ;
wire \rd_ram_rd_addr[2]~q ;
wire \rd_ram_wr_addr[1]~0_combout ;
wire \rd_ram_wr_addr[2]~1_combout ;
wire \rd_ram_wr_addr[3]~2_combout ;
wire \rd_ram_rd_addr[1]~0_combout ;
wire \rd_ram_rd_addr[2]~1_combout ;
wire \rd_ram_wr_addr[1]~_wirecell_combout ;
wire \rd_ram_wr_addr[2]~_wirecell_combout ;


ddr3_int_altsyncram_3 \half_rate_ram_gen.altsyncram_component (
	.q_b({q_b_127,q_b_126,q_b_125,q_b_124,q_b_123,q_b_122,q_b_121,q_b_120,q_b_119,q_b_118,q_b_117,q_b_116,q_b_115,q_b_114,q_b_113,q_b_112,q_b_111,q_b_110,q_b_109,q_b_108,q_b_107,q_b_106,q_b_105,q_b_104,q_b_103,q_b_102,q_b_101,q_b_100,q_b_99,q_b_98,q_b_97,q_b_96,q_b_95,q_b_94,q_b_93,q_b_92,q_b_91,q_b_90,
q_b_89,q_b_88,q_b_87,q_b_86,q_b_85,q_b_84,q_b_83,q_b_82,q_b_81,q_b_80,q_b_79,q_b_78,q_b_77,q_b_76,q_b_75,q_b_74,q_b_73,q_b_72,q_b_71,q_b_70,q_b_69,q_b_68,q_b_67,q_b_66,q_b_65,q_b_64,q_b_63,q_b_62,q_b_61,q_b_60,q_b_59,q_b_58,q_b_57,q_b_56,q_b_55,q_b_54,q_b_53,q_b_52,q_b_51,q_b_50,q_b_49,q_b_48,
q_b_47,q_b_46,q_b_45,q_b_44,q_b_43,q_b_42,q_b_41,q_b_40,q_b_39,q_b_38,q_b_37,q_b_36,q_b_35,q_b_34,q_b_33,q_b_32,q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,
q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.clock1(clk_0),
	.clock0(clk_4),
	.data_a({dio_rdata_l_2x_31,dio_rdata_l_2x_30,dio_rdata_l_2x_29,dio_rdata_l_2x_28,dio_rdata_l_2x_27,dio_rdata_l_2x_26,dio_rdata_l_2x_25,dio_rdata_l_2x_24,dio_rdata_h_2x_31,dio_rdata_h_2x_30,dio_rdata_h_2x_29,dio_rdata_h_2x_28,dio_rdata_h_2x_27,dio_rdata_h_2x_26,dio_rdata_h_2x_25,
dio_rdata_h_2x_24,dio_rdata_l_2x_23,dio_rdata_l_2x_22,dio_rdata_l_2x_21,dio_rdata_l_2x_20,dio_rdata_l_2x_19,dio_rdata_l_2x_18,dio_rdata_l_2x_17,dio_rdata_l_2x_16,dio_rdata_h_2x_23,dio_rdata_h_2x_22,dio_rdata_h_2x_21,dio_rdata_h_2x_20,dio_rdata_h_2x_19,dio_rdata_h_2x_18,
dio_rdata_h_2x_17,dio_rdata_h_2x_16,dio_rdata_l_2x_15,dio_rdata_l_2x_14,dio_rdata_l_2x_13,dio_rdata_l_2x_12,dio_rdata_l_2x_11,dio_rdata_l_2x_10,dio_rdata_l_2x_9,dio_rdata_l_2x_8,dio_rdata_h_2x_15,dio_rdata_h_2x_14,dio_rdata_h_2x_13,dio_rdata_h_2x_12,dio_rdata_h_2x_11,
dio_rdata_h_2x_10,dio_rdata_h_2x_9,dio_rdata_h_2x_8,dio_rdata_l_2x_7,dio_rdata_l_2x_6,dio_rdata_l_2x_5,dio_rdata_l_2x_4,dio_rdata_l_2x_3,dio_rdata_l_2x_2,dio_rdata_l_2x_1,dio_rdata_l_2x_0,dio_rdata_h_2x_7,dio_rdata_h_2x_6,dio_rdata_h_2x_5,dio_rdata_h_2x_4,
dio_rdata_h_2x_3,dio_rdata_h_2x_2,dio_rdata_h_2x_1,dio_rdata_h_2x_0}),
	.address_a({gnd,\rd_ram_wr_addr[3]~q ,\rd_ram_wr_addr[2]~_wirecell_combout ,\rd_ram_wr_addr[1]~_wirecell_combout ,rd_addr_2x_0}),
	.address_b({gnd,gnd,gnd,\rd_ram_rd_addr[2]~q ,\rd_ram_rd_addr[1]~q ,rd_addr_0}));

dffeas \rd_ram_wr_addr[1] (
	.clk(clk_4),
	.d(\rd_ram_wr_addr[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset_resync_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_ram_wr_addr[1]~q ),
	.prn(vcc));
defparam \rd_ram_wr_addr[1] .is_wysiwyg = "true";
defparam \rd_ram_wr_addr[1] .power_up = "low";

dffeas \rd_ram_wr_addr[2] (
	.clk(clk_4),
	.d(\rd_ram_wr_addr[2]~1_combout ),
	.asdata(vcc),
	.clrn(reset_resync_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_ram_wr_addr[2]~q ),
	.prn(vcc));
defparam \rd_ram_wr_addr[2] .is_wysiwyg = "true";
defparam \rd_ram_wr_addr[2] .power_up = "low";

dffeas \rd_ram_wr_addr[3] (
	.clk(clk_4),
	.d(\rd_ram_wr_addr[3]~2_combout ),
	.asdata(vcc),
	.clrn(reset_resync_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_ram_wr_addr[3]~q ),
	.prn(vcc));
defparam \rd_ram_wr_addr[3] .is_wysiwyg = "true";
defparam \rd_ram_wr_addr[3] .power_up = "low";

dffeas \rd_ram_rd_addr[1] (
	.clk(clk_0),
	.d(\rd_ram_rd_addr[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_ram_rd_addr[1]~q ),
	.prn(vcc));
defparam \rd_ram_rd_addr[1] .is_wysiwyg = "true";
defparam \rd_ram_rd_addr[1] .power_up = "low";

dffeas \rd_ram_rd_addr[2] (
	.clk(clk_0),
	.d(\rd_ram_rd_addr[2]~1_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_ram_rd_addr[2]~q ),
	.prn(vcc));
defparam \rd_ram_rd_addr[2] .is_wysiwyg = "true";
defparam \rd_ram_rd_addr[2] .power_up = "low";

arriaii_lcell_comb \rd_ram_wr_addr[1]~0 (
	.dataa(!rd_addr_2x_0),
	.datab(!\rd_ram_wr_addr[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rd_ram_wr_addr[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_ram_wr_addr[1]~0 .extended_lut = "off";
defparam \rd_ram_wr_addr[1]~0 .lut_mask = 64'h6666666666666666;
defparam \rd_ram_wr_addr[1]~0 .shared_arith = "off";

arriaii_lcell_comb \rd_ram_wr_addr[2]~1 (
	.dataa(!rd_addr_2x_0),
	.datab(!\rd_ram_wr_addr[1]~q ),
	.datac(!\rd_ram_wr_addr[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rd_ram_wr_addr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_ram_wr_addr[2]~1 .extended_lut = "off";
defparam \rd_ram_wr_addr[2]~1 .lut_mask = 64'h4B4B4B4B4B4B4B4B;
defparam \rd_ram_wr_addr[2]~1 .shared_arith = "off";

arriaii_lcell_comb \rd_ram_wr_addr[3]~2 (
	.dataa(!rd_addr_2x_0),
	.datab(!\rd_ram_wr_addr[1]~q ),
	.datac(!\rd_ram_wr_addr[2]~q ),
	.datad(!\rd_ram_wr_addr[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rd_ram_wr_addr[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_ram_wr_addr[3]~2 .extended_lut = "off";
defparam \rd_ram_wr_addr[3]~2 .lut_mask = 64'h40BF40BF40BF40BF;
defparam \rd_ram_wr_addr[3]~2 .shared_arith = "off";

arriaii_lcell_comb \rd_ram_rd_addr[1]~0 (
	.dataa(!rd_addr_0),
	.datab(!\rd_ram_rd_addr[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rd_ram_rd_addr[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_ram_rd_addr[1]~0 .extended_lut = "off";
defparam \rd_ram_rd_addr[1]~0 .lut_mask = 64'h6666666666666666;
defparam \rd_ram_rd_addr[1]~0 .shared_arith = "off";

arriaii_lcell_comb \rd_ram_rd_addr[2]~1 (
	.dataa(!rd_addr_0),
	.datab(!\rd_ram_rd_addr[1]~q ),
	.datac(!\rd_ram_rd_addr[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rd_ram_rd_addr[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_ram_rd_addr[2]~1 .extended_lut = "off";
defparam \rd_ram_rd_addr[2]~1 .lut_mask = 64'h1E1E1E1E1E1E1E1E;
defparam \rd_ram_rd_addr[2]~1 .shared_arith = "off";

arriaii_lcell_comb \rd_ram_wr_addr[1]~_wirecell (
	.dataa(!\rd_ram_wr_addr[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rd_ram_wr_addr[1]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_ram_wr_addr[1]~_wirecell .extended_lut = "off";
defparam \rd_ram_wr_addr[1]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rd_ram_wr_addr[1]~_wirecell .shared_arith = "off";

arriaii_lcell_comb \rd_ram_wr_addr[2]~_wirecell (
	.dataa(!\rd_ram_wr_addr[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rd_ram_wr_addr[2]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_ram_wr_addr[2]~_wirecell .extended_lut = "off";
defparam \rd_ram_wr_addr[2]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rd_ram_wr_addr[2]~_wirecell .shared_arith = "off";

endmodule

module ddr3_int_altsyncram_3 (
	q_b,
	clock1,
	clock0,
	data_a,
	address_a,
	address_b)/* synthesis synthesis_greybox=0 */;
output 	[127:0] q_b;
input 	clock1;
input 	clock0;
input 	[63:0] data_a;
input 	[4:0] address_a;
input 	[5:0] address_b;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_altsyncram_lbh1 auto_generated(
	.q_b({q_b[127],q_b[126],q_b[125],q_b[124],q_b[123],q_b[122],q_b[121],q_b[120],q_b[119],q_b[118],q_b[117],q_b[116],q_b[115],q_b[114],q_b[113],q_b[112],q_b[111],q_b[110],q_b[109],q_b[108],q_b[107],q_b[106],q_b[105],q_b[104],q_b[103],q_b[102],q_b[101],q_b[100],q_b[99],q_b[98],q_b[97],q_b[96],q_b[95],q_b[94],q_b[93],q_b[92],q_b[91],q_b[90],q_b[89],q_b[88],q_b[87],q_b[86],q_b[85],q_b[84],q_b[83],q_b[82],q_b[81],q_b[80],q_b[79],q_b[78],q_b[77],q_b[76],q_b[75],q_b[74],q_b[73],q_b[72],q_b[71],q_b[70],q_b[69],q_b[68],q_b[67],q_b[66],q_b[65],q_b[64],q_b[63],q_b[62],q_b[61],q_b[60],q_b[59],q_b[58],q_b[57],q_b[56],q_b[55],q_b[54],q_b[53],q_b[52],q_b[51],q_b[50],q_b[49],q_b[48],q_b[47],q_b[46],q_b[45],q_b[44],q_b[43],
q_b[42],q_b[41],q_b[40],q_b[39],q_b[38],q_b[37],q_b[36],q_b[35],q_b[34],q_b[33],q_b[32],q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.clock1(clock1),
	.clock0(clock0),
	.data_a({data_a[63],data_a[62],data_a[61],data_a[60],data_a[59],data_a[58],data_a[57],data_a[56],data_a[55],data_a[54],data_a[53],data_a[52],data_a[51],data_a[50],data_a[49],data_a[48],data_a[47],data_a[46],data_a[45],data_a[44],data_a[43],data_a[42],data_a[41],data_a[40],data_a[39],data_a[38],data_a[37],data_a[36],data_a[35],data_a[34],data_a[33],data_a[32],data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],
data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[2],address_b[1],address_b[0]}));

endmodule

module ddr3_int_altsyncram_lbh1 (
	q_b,
	clock1,
	clock0,
	data_a,
	address_a,
	address_b)/* synthesis synthesis_greybox=0 */;
output 	[127:0] q_b;
input 	clock1;
input 	clock0;
input 	[63:0] data_a;
input 	[3:0] address_a;
input 	[2:0] address_b;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a32_PORTBDATAOUT_bus;
wire [143:0] ram_block1a33_PORTBDATAOUT_bus;
wire [143:0] ram_block1a34_PORTBDATAOUT_bus;
wire [143:0] ram_block1a35_PORTBDATAOUT_bus;
wire [143:0] ram_block1a36_PORTBDATAOUT_bus;
wire [143:0] ram_block1a37_PORTBDATAOUT_bus;
wire [143:0] ram_block1a38_PORTBDATAOUT_bus;
wire [143:0] ram_block1a39_PORTBDATAOUT_bus;
wire [143:0] ram_block1a48_PORTBDATAOUT_bus;
wire [143:0] ram_block1a49_PORTBDATAOUT_bus;
wire [143:0] ram_block1a50_PORTBDATAOUT_bus;
wire [143:0] ram_block1a51_PORTBDATAOUT_bus;
wire [143:0] ram_block1a52_PORTBDATAOUT_bus;
wire [143:0] ram_block1a53_PORTBDATAOUT_bus;
wire [143:0] ram_block1a54_PORTBDATAOUT_bus;
wire [143:0] ram_block1a55_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a40_PORTBDATAOUT_bus;
wire [143:0] ram_block1a41_PORTBDATAOUT_bus;
wire [143:0] ram_block1a42_PORTBDATAOUT_bus;
wire [143:0] ram_block1a43_PORTBDATAOUT_bus;
wire [143:0] ram_block1a44_PORTBDATAOUT_bus;
wire [143:0] ram_block1a45_PORTBDATAOUT_bus;
wire [143:0] ram_block1a46_PORTBDATAOUT_bus;
wire [143:0] ram_block1a47_PORTBDATAOUT_bus;
wire [143:0] ram_block1a56_PORTBDATAOUT_bus;
wire [143:0] ram_block1a57_PORTBDATAOUT_bus;
wire [143:0] ram_block1a58_PORTBDATAOUT_bus;
wire [143:0] ram_block1a59_PORTBDATAOUT_bus;
wire [143:0] ram_block1a60_PORTBDATAOUT_bus;
wire [143:0] ram_block1a61_PORTBDATAOUT_bus;
wire [143:0] ram_block1a62_PORTBDATAOUT_bus;
wire [143:0] ram_block1a63_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];
assign q_b[64] = ram_block1a0_PORTBDATAOUT_bus[1];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];
assign q_b[65] = ram_block1a1_PORTBDATAOUT_bus[1];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];
assign q_b[66] = ram_block1a2_PORTBDATAOUT_bus[1];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];
assign q_b[67] = ram_block1a3_PORTBDATAOUT_bus[1];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];
assign q_b[68] = ram_block1a4_PORTBDATAOUT_bus[1];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];
assign q_b[69] = ram_block1a5_PORTBDATAOUT_bus[1];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];
assign q_b[70] = ram_block1a6_PORTBDATAOUT_bus[1];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];
assign q_b[71] = ram_block1a7_PORTBDATAOUT_bus[1];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];
assign q_b[80] = ram_block1a16_PORTBDATAOUT_bus[1];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];
assign q_b[81] = ram_block1a17_PORTBDATAOUT_bus[1];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];
assign q_b[82] = ram_block1a18_PORTBDATAOUT_bus[1];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];
assign q_b[83] = ram_block1a19_PORTBDATAOUT_bus[1];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];
assign q_b[84] = ram_block1a20_PORTBDATAOUT_bus[1];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];
assign q_b[85] = ram_block1a21_PORTBDATAOUT_bus[1];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];
assign q_b[86] = ram_block1a22_PORTBDATAOUT_bus[1];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];
assign q_b[87] = ram_block1a23_PORTBDATAOUT_bus[1];

assign q_b[32] = ram_block1a32_PORTBDATAOUT_bus[0];
assign q_b[96] = ram_block1a32_PORTBDATAOUT_bus[1];

assign q_b[33] = ram_block1a33_PORTBDATAOUT_bus[0];
assign q_b[97] = ram_block1a33_PORTBDATAOUT_bus[1];

assign q_b[34] = ram_block1a34_PORTBDATAOUT_bus[0];
assign q_b[98] = ram_block1a34_PORTBDATAOUT_bus[1];

assign q_b[35] = ram_block1a35_PORTBDATAOUT_bus[0];
assign q_b[99] = ram_block1a35_PORTBDATAOUT_bus[1];

assign q_b[36] = ram_block1a36_PORTBDATAOUT_bus[0];
assign q_b[100] = ram_block1a36_PORTBDATAOUT_bus[1];

assign q_b[37] = ram_block1a37_PORTBDATAOUT_bus[0];
assign q_b[101] = ram_block1a37_PORTBDATAOUT_bus[1];

assign q_b[38] = ram_block1a38_PORTBDATAOUT_bus[0];
assign q_b[102] = ram_block1a38_PORTBDATAOUT_bus[1];

assign q_b[39] = ram_block1a39_PORTBDATAOUT_bus[0];
assign q_b[103] = ram_block1a39_PORTBDATAOUT_bus[1];

assign q_b[48] = ram_block1a48_PORTBDATAOUT_bus[0];
assign q_b[112] = ram_block1a48_PORTBDATAOUT_bus[1];

assign q_b[49] = ram_block1a49_PORTBDATAOUT_bus[0];
assign q_b[113] = ram_block1a49_PORTBDATAOUT_bus[1];

assign q_b[50] = ram_block1a50_PORTBDATAOUT_bus[0];
assign q_b[114] = ram_block1a50_PORTBDATAOUT_bus[1];

assign q_b[51] = ram_block1a51_PORTBDATAOUT_bus[0];
assign q_b[115] = ram_block1a51_PORTBDATAOUT_bus[1];

assign q_b[52] = ram_block1a52_PORTBDATAOUT_bus[0];
assign q_b[116] = ram_block1a52_PORTBDATAOUT_bus[1];

assign q_b[53] = ram_block1a53_PORTBDATAOUT_bus[0];
assign q_b[117] = ram_block1a53_PORTBDATAOUT_bus[1];

assign q_b[54] = ram_block1a54_PORTBDATAOUT_bus[0];
assign q_b[118] = ram_block1a54_PORTBDATAOUT_bus[1];

assign q_b[55] = ram_block1a55_PORTBDATAOUT_bus[0];
assign q_b[119] = ram_block1a55_PORTBDATAOUT_bus[1];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];
assign q_b[72] = ram_block1a8_PORTBDATAOUT_bus[1];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];
assign q_b[73] = ram_block1a9_PORTBDATAOUT_bus[1];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];
assign q_b[74] = ram_block1a10_PORTBDATAOUT_bus[1];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];
assign q_b[75] = ram_block1a11_PORTBDATAOUT_bus[1];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];
assign q_b[76] = ram_block1a12_PORTBDATAOUT_bus[1];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];
assign q_b[77] = ram_block1a13_PORTBDATAOUT_bus[1];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];
assign q_b[78] = ram_block1a14_PORTBDATAOUT_bus[1];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];
assign q_b[79] = ram_block1a15_PORTBDATAOUT_bus[1];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];
assign q_b[88] = ram_block1a24_PORTBDATAOUT_bus[1];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];
assign q_b[89] = ram_block1a25_PORTBDATAOUT_bus[1];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];
assign q_b[90] = ram_block1a26_PORTBDATAOUT_bus[1];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];
assign q_b[91] = ram_block1a27_PORTBDATAOUT_bus[1];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];
assign q_b[92] = ram_block1a28_PORTBDATAOUT_bus[1];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];
assign q_b[93] = ram_block1a29_PORTBDATAOUT_bus[1];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];
assign q_b[94] = ram_block1a30_PORTBDATAOUT_bus[1];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];
assign q_b[95] = ram_block1a31_PORTBDATAOUT_bus[1];

assign q_b[40] = ram_block1a40_PORTBDATAOUT_bus[0];
assign q_b[104] = ram_block1a40_PORTBDATAOUT_bus[1];

assign q_b[41] = ram_block1a41_PORTBDATAOUT_bus[0];
assign q_b[105] = ram_block1a41_PORTBDATAOUT_bus[1];

assign q_b[42] = ram_block1a42_PORTBDATAOUT_bus[0];
assign q_b[106] = ram_block1a42_PORTBDATAOUT_bus[1];

assign q_b[43] = ram_block1a43_PORTBDATAOUT_bus[0];
assign q_b[107] = ram_block1a43_PORTBDATAOUT_bus[1];

assign q_b[44] = ram_block1a44_PORTBDATAOUT_bus[0];
assign q_b[108] = ram_block1a44_PORTBDATAOUT_bus[1];

assign q_b[45] = ram_block1a45_PORTBDATAOUT_bus[0];
assign q_b[109] = ram_block1a45_PORTBDATAOUT_bus[1];

assign q_b[46] = ram_block1a46_PORTBDATAOUT_bus[0];
assign q_b[110] = ram_block1a46_PORTBDATAOUT_bus[1];

assign q_b[47] = ram_block1a47_PORTBDATAOUT_bus[0];
assign q_b[111] = ram_block1a47_PORTBDATAOUT_bus[1];

assign q_b[56] = ram_block1a56_PORTBDATAOUT_bus[0];
assign q_b[120] = ram_block1a56_PORTBDATAOUT_bus[1];

assign q_b[57] = ram_block1a57_PORTBDATAOUT_bus[0];
assign q_b[121] = ram_block1a57_PORTBDATAOUT_bus[1];

assign q_b[58] = ram_block1a58_PORTBDATAOUT_bus[0];
assign q_b[122] = ram_block1a58_PORTBDATAOUT_bus[1];

assign q_b[59] = ram_block1a59_PORTBDATAOUT_bus[0];
assign q_b[123] = ram_block1a59_PORTBDATAOUT_bus[1];

assign q_b[60] = ram_block1a60_PORTBDATAOUT_bus[0];
assign q_b[124] = ram_block1a60_PORTBDATAOUT_bus[1];

assign q_b[61] = ram_block1a61_PORTBDATAOUT_bus[0];
assign q_b[125] = ram_block1a61_PORTBDATAOUT_bus[1];

assign q_b[62] = ram_block1a62_PORTBDATAOUT_bus[0];
assign q_b[126] = ram_block1a62_PORTBDATAOUT_bus[1];

assign q_b[63] = ram_block1a63_PORTBDATAOUT_bus[0];
assign q_b[127] = ram_block1a63_PORTBDATAOUT_bus[1];

arriaii_ram_block ram_block1a0(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena2";
defparam ram_block1a0.clk1_core_clock_enable = "ena3";
defparam ram_block1a0.clk1_input_clock_enable = "ena3";
defparam ram_block1a0.clock_duty_cycle_dependence = "on";
defparam ram_block1a0.data_interleave_offset_in_bits = 64;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 4;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 15;
defparam ram_block1a0.port_a_logical_ram_depth = 16;
defparam ram_block1a0.port_a_logical_ram_width = 64;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 3;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "clock1";
defparam ram_block1a0.port_b_data_width = 2;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 7;
defparam ram_block1a0.port_b_logical_ram_depth = 8;
defparam ram_block1a0.port_b_logical_ram_width = 128;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

arriaii_ram_block ram_block1a1(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena2";
defparam ram_block1a1.clk1_core_clock_enable = "ena3";
defparam ram_block1a1.clk1_input_clock_enable = "ena3";
defparam ram_block1a1.clock_duty_cycle_dependence = "on";
defparam ram_block1a1.data_interleave_offset_in_bits = 64;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 4;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 15;
defparam ram_block1a1.port_a_logical_ram_depth = 16;
defparam ram_block1a1.port_a_logical_ram_width = 64;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 3;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "clock1";
defparam ram_block1a1.port_b_data_width = 2;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 7;
defparam ram_block1a1.port_b_logical_ram_depth = 8;
defparam ram_block1a1.port_b_logical_ram_width = 128;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

arriaii_ram_block ram_block1a2(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena2";
defparam ram_block1a2.clk1_core_clock_enable = "ena3";
defparam ram_block1a2.clk1_input_clock_enable = "ena3";
defparam ram_block1a2.clock_duty_cycle_dependence = "on";
defparam ram_block1a2.data_interleave_offset_in_bits = 64;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 4;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 15;
defparam ram_block1a2.port_a_logical_ram_depth = 16;
defparam ram_block1a2.port_a_logical_ram_width = 64;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 3;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "clock1";
defparam ram_block1a2.port_b_data_width = 2;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 7;
defparam ram_block1a2.port_b_logical_ram_depth = 8;
defparam ram_block1a2.port_b_logical_ram_width = 128;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

arriaii_ram_block ram_block1a3(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena2";
defparam ram_block1a3.clk1_core_clock_enable = "ena3";
defparam ram_block1a3.clk1_input_clock_enable = "ena3";
defparam ram_block1a3.clock_duty_cycle_dependence = "on";
defparam ram_block1a3.data_interleave_offset_in_bits = 64;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 4;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 15;
defparam ram_block1a3.port_a_logical_ram_depth = 16;
defparam ram_block1a3.port_a_logical_ram_width = 64;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 3;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "clock1";
defparam ram_block1a3.port_b_data_width = 2;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 7;
defparam ram_block1a3.port_b_logical_ram_depth = 8;
defparam ram_block1a3.port_b_logical_ram_width = 128;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

arriaii_ram_block ram_block1a4(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena2";
defparam ram_block1a4.clk1_core_clock_enable = "ena3";
defparam ram_block1a4.clk1_input_clock_enable = "ena3";
defparam ram_block1a4.clock_duty_cycle_dependence = "on";
defparam ram_block1a4.data_interleave_offset_in_bits = 64;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 4;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 15;
defparam ram_block1a4.port_a_logical_ram_depth = 16;
defparam ram_block1a4.port_a_logical_ram_width = 64;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 3;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "clock1";
defparam ram_block1a4.port_b_data_width = 2;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 7;
defparam ram_block1a4.port_b_logical_ram_depth = 8;
defparam ram_block1a4.port_b_logical_ram_width = 128;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

arriaii_ram_block ram_block1a5(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena2";
defparam ram_block1a5.clk1_core_clock_enable = "ena3";
defparam ram_block1a5.clk1_input_clock_enable = "ena3";
defparam ram_block1a5.clock_duty_cycle_dependence = "on";
defparam ram_block1a5.data_interleave_offset_in_bits = 64;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 4;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 15;
defparam ram_block1a5.port_a_logical_ram_depth = 16;
defparam ram_block1a5.port_a_logical_ram_width = 64;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 3;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "clock1";
defparam ram_block1a5.port_b_data_width = 2;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 7;
defparam ram_block1a5.port_b_logical_ram_depth = 8;
defparam ram_block1a5.port_b_logical_ram_width = 128;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

arriaii_ram_block ram_block1a6(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena2";
defparam ram_block1a6.clk1_core_clock_enable = "ena3";
defparam ram_block1a6.clk1_input_clock_enable = "ena3";
defparam ram_block1a6.clock_duty_cycle_dependence = "on";
defparam ram_block1a6.data_interleave_offset_in_bits = 64;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 4;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 15;
defparam ram_block1a6.port_a_logical_ram_depth = 16;
defparam ram_block1a6.port_a_logical_ram_width = 64;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 3;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "clock1";
defparam ram_block1a6.port_b_data_width = 2;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 7;
defparam ram_block1a6.port_b_logical_ram_depth = 8;
defparam ram_block1a6.port_b_logical_ram_width = 128;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

arriaii_ram_block ram_block1a7(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena2";
defparam ram_block1a7.clk1_core_clock_enable = "ena3";
defparam ram_block1a7.clk1_input_clock_enable = "ena3";
defparam ram_block1a7.clock_duty_cycle_dependence = "on";
defparam ram_block1a7.data_interleave_offset_in_bits = 64;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 4;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 15;
defparam ram_block1a7.port_a_logical_ram_depth = 16;
defparam ram_block1a7.port_a_logical_ram_width = 64;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 3;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "clock1";
defparam ram_block1a7.port_b_data_width = 2;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 7;
defparam ram_block1a7.port_b_logical_ram_depth = 8;
defparam ram_block1a7.port_b_logical_ram_width = 128;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

arriaii_ram_block ram_block1a16(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena2";
defparam ram_block1a16.clk1_core_clock_enable = "ena3";
defparam ram_block1a16.clk1_input_clock_enable = "ena3";
defparam ram_block1a16.clock_duty_cycle_dependence = "on";
defparam ram_block1a16.data_interleave_offset_in_bits = 64;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 4;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 15;
defparam ram_block1a16.port_a_logical_ram_depth = 16;
defparam ram_block1a16.port_a_logical_ram_width = 64;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 3;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "clock1";
defparam ram_block1a16.port_b_data_width = 2;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 7;
defparam ram_block1a16.port_b_logical_ram_depth = 8;
defparam ram_block1a16.port_b_logical_ram_width = 128;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

arriaii_ram_block ram_block1a17(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena2";
defparam ram_block1a17.clk1_core_clock_enable = "ena3";
defparam ram_block1a17.clk1_input_clock_enable = "ena3";
defparam ram_block1a17.clock_duty_cycle_dependence = "on";
defparam ram_block1a17.data_interleave_offset_in_bits = 64;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 4;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 15;
defparam ram_block1a17.port_a_logical_ram_depth = 16;
defparam ram_block1a17.port_a_logical_ram_width = 64;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 3;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "clock1";
defparam ram_block1a17.port_b_data_width = 2;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 7;
defparam ram_block1a17.port_b_logical_ram_depth = 8;
defparam ram_block1a17.port_b_logical_ram_width = 128;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

arriaii_ram_block ram_block1a18(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena2";
defparam ram_block1a18.clk1_core_clock_enable = "ena3";
defparam ram_block1a18.clk1_input_clock_enable = "ena3";
defparam ram_block1a18.clock_duty_cycle_dependence = "on";
defparam ram_block1a18.data_interleave_offset_in_bits = 64;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 4;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 15;
defparam ram_block1a18.port_a_logical_ram_depth = 16;
defparam ram_block1a18.port_a_logical_ram_width = 64;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 3;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "clock1";
defparam ram_block1a18.port_b_data_width = 2;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 7;
defparam ram_block1a18.port_b_logical_ram_depth = 8;
defparam ram_block1a18.port_b_logical_ram_width = 128;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

arriaii_ram_block ram_block1a19(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena2";
defparam ram_block1a19.clk1_core_clock_enable = "ena3";
defparam ram_block1a19.clk1_input_clock_enable = "ena3";
defparam ram_block1a19.clock_duty_cycle_dependence = "on";
defparam ram_block1a19.data_interleave_offset_in_bits = 64;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 4;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 15;
defparam ram_block1a19.port_a_logical_ram_depth = 16;
defparam ram_block1a19.port_a_logical_ram_width = 64;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 3;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "clock1";
defparam ram_block1a19.port_b_data_width = 2;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 7;
defparam ram_block1a19.port_b_logical_ram_depth = 8;
defparam ram_block1a19.port_b_logical_ram_width = 128;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

arriaii_ram_block ram_block1a20(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena2";
defparam ram_block1a20.clk1_core_clock_enable = "ena3";
defparam ram_block1a20.clk1_input_clock_enable = "ena3";
defparam ram_block1a20.clock_duty_cycle_dependence = "on";
defparam ram_block1a20.data_interleave_offset_in_bits = 64;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 4;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 15;
defparam ram_block1a20.port_a_logical_ram_depth = 16;
defparam ram_block1a20.port_a_logical_ram_width = 64;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 3;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "clock1";
defparam ram_block1a20.port_b_data_width = 2;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 7;
defparam ram_block1a20.port_b_logical_ram_depth = 8;
defparam ram_block1a20.port_b_logical_ram_width = 128;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

arriaii_ram_block ram_block1a21(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena2";
defparam ram_block1a21.clk1_core_clock_enable = "ena3";
defparam ram_block1a21.clk1_input_clock_enable = "ena3";
defparam ram_block1a21.clock_duty_cycle_dependence = "on";
defparam ram_block1a21.data_interleave_offset_in_bits = 64;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 4;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 15;
defparam ram_block1a21.port_a_logical_ram_depth = 16;
defparam ram_block1a21.port_a_logical_ram_width = 64;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 3;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "clock1";
defparam ram_block1a21.port_b_data_width = 2;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 7;
defparam ram_block1a21.port_b_logical_ram_depth = 8;
defparam ram_block1a21.port_b_logical_ram_width = 128;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

arriaii_ram_block ram_block1a22(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena2";
defparam ram_block1a22.clk1_core_clock_enable = "ena3";
defparam ram_block1a22.clk1_input_clock_enable = "ena3";
defparam ram_block1a22.clock_duty_cycle_dependence = "on";
defparam ram_block1a22.data_interleave_offset_in_bits = 64;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 4;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 15;
defparam ram_block1a22.port_a_logical_ram_depth = 16;
defparam ram_block1a22.port_a_logical_ram_width = 64;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock1";
defparam ram_block1a22.port_b_address_width = 3;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "clock1";
defparam ram_block1a22.port_b_data_width = 2;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 7;
defparam ram_block1a22.port_b_logical_ram_depth = 8;
defparam ram_block1a22.port_b_logical_ram_width = 128;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock1";
defparam ram_block1a22.ram_block_type = "auto";

arriaii_ram_block ram_block1a23(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena2";
defparam ram_block1a23.clk1_core_clock_enable = "ena3";
defparam ram_block1a23.clk1_input_clock_enable = "ena3";
defparam ram_block1a23.clock_duty_cycle_dependence = "on";
defparam ram_block1a23.data_interleave_offset_in_bits = 64;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 4;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 15;
defparam ram_block1a23.port_a_logical_ram_depth = 16;
defparam ram_block1a23.port_a_logical_ram_width = 64;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock1";
defparam ram_block1a23.port_b_address_width = 3;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "clock1";
defparam ram_block1a23.port_b_data_width = 2;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 7;
defparam ram_block1a23.port_b_logical_ram_depth = 8;
defparam ram_block1a23.port_b_logical_ram_width = 128;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock1";
defparam ram_block1a23.ram_block_type = "auto";

arriaii_ram_block ram_block1a32(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[32]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a32_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a32.clk0_core_clock_enable = "ena0";
defparam ram_block1a32.clk0_input_clock_enable = "ena2";
defparam ram_block1a32.clk1_core_clock_enable = "ena3";
defparam ram_block1a32.clk1_input_clock_enable = "ena3";
defparam ram_block1a32.clock_duty_cycle_dependence = "on";
defparam ram_block1a32.data_interleave_offset_in_bits = 64;
defparam ram_block1a32.data_interleave_width_in_bits = 1;
defparam ram_block1a32.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a32.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a32.operation_mode = "dual_port";
defparam ram_block1a32.port_a_address_clear = "none";
defparam ram_block1a32.port_a_address_width = 4;
defparam ram_block1a32.port_a_data_out_clear = "none";
defparam ram_block1a32.port_a_data_out_clock = "none";
defparam ram_block1a32.port_a_data_width = 1;
defparam ram_block1a32.port_a_first_address = 0;
defparam ram_block1a32.port_a_first_bit_number = 32;
defparam ram_block1a32.port_a_last_address = 15;
defparam ram_block1a32.port_a_logical_ram_depth = 16;
defparam ram_block1a32.port_a_logical_ram_width = 64;
defparam ram_block1a32.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a32.port_b_address_clear = "none";
defparam ram_block1a32.port_b_address_clock = "clock1";
defparam ram_block1a32.port_b_address_width = 3;
defparam ram_block1a32.port_b_data_out_clear = "none";
defparam ram_block1a32.port_b_data_out_clock = "clock1";
defparam ram_block1a32.port_b_data_width = 2;
defparam ram_block1a32.port_b_first_address = 0;
defparam ram_block1a32.port_b_first_bit_number = 32;
defparam ram_block1a32.port_b_last_address = 7;
defparam ram_block1a32.port_b_logical_ram_depth = 8;
defparam ram_block1a32.port_b_logical_ram_width = 128;
defparam ram_block1a32.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a32.port_b_read_enable_clock = "clock1";
defparam ram_block1a32.ram_block_type = "auto";

arriaii_ram_block ram_block1a33(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[33]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a33_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a33.clk0_core_clock_enable = "ena0";
defparam ram_block1a33.clk0_input_clock_enable = "ena2";
defparam ram_block1a33.clk1_core_clock_enable = "ena3";
defparam ram_block1a33.clk1_input_clock_enable = "ena3";
defparam ram_block1a33.clock_duty_cycle_dependence = "on";
defparam ram_block1a33.data_interleave_offset_in_bits = 64;
defparam ram_block1a33.data_interleave_width_in_bits = 1;
defparam ram_block1a33.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a33.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a33.operation_mode = "dual_port";
defparam ram_block1a33.port_a_address_clear = "none";
defparam ram_block1a33.port_a_address_width = 4;
defparam ram_block1a33.port_a_data_out_clear = "none";
defparam ram_block1a33.port_a_data_out_clock = "none";
defparam ram_block1a33.port_a_data_width = 1;
defparam ram_block1a33.port_a_first_address = 0;
defparam ram_block1a33.port_a_first_bit_number = 33;
defparam ram_block1a33.port_a_last_address = 15;
defparam ram_block1a33.port_a_logical_ram_depth = 16;
defparam ram_block1a33.port_a_logical_ram_width = 64;
defparam ram_block1a33.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a33.port_b_address_clear = "none";
defparam ram_block1a33.port_b_address_clock = "clock1";
defparam ram_block1a33.port_b_address_width = 3;
defparam ram_block1a33.port_b_data_out_clear = "none";
defparam ram_block1a33.port_b_data_out_clock = "clock1";
defparam ram_block1a33.port_b_data_width = 2;
defparam ram_block1a33.port_b_first_address = 0;
defparam ram_block1a33.port_b_first_bit_number = 33;
defparam ram_block1a33.port_b_last_address = 7;
defparam ram_block1a33.port_b_logical_ram_depth = 8;
defparam ram_block1a33.port_b_logical_ram_width = 128;
defparam ram_block1a33.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a33.port_b_read_enable_clock = "clock1";
defparam ram_block1a33.ram_block_type = "auto";

arriaii_ram_block ram_block1a34(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[34]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a34_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a34.clk0_core_clock_enable = "ena0";
defparam ram_block1a34.clk0_input_clock_enable = "ena2";
defparam ram_block1a34.clk1_core_clock_enable = "ena3";
defparam ram_block1a34.clk1_input_clock_enable = "ena3";
defparam ram_block1a34.clock_duty_cycle_dependence = "on";
defparam ram_block1a34.data_interleave_offset_in_bits = 64;
defparam ram_block1a34.data_interleave_width_in_bits = 1;
defparam ram_block1a34.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a34.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a34.operation_mode = "dual_port";
defparam ram_block1a34.port_a_address_clear = "none";
defparam ram_block1a34.port_a_address_width = 4;
defparam ram_block1a34.port_a_data_out_clear = "none";
defparam ram_block1a34.port_a_data_out_clock = "none";
defparam ram_block1a34.port_a_data_width = 1;
defparam ram_block1a34.port_a_first_address = 0;
defparam ram_block1a34.port_a_first_bit_number = 34;
defparam ram_block1a34.port_a_last_address = 15;
defparam ram_block1a34.port_a_logical_ram_depth = 16;
defparam ram_block1a34.port_a_logical_ram_width = 64;
defparam ram_block1a34.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a34.port_b_address_clear = "none";
defparam ram_block1a34.port_b_address_clock = "clock1";
defparam ram_block1a34.port_b_address_width = 3;
defparam ram_block1a34.port_b_data_out_clear = "none";
defparam ram_block1a34.port_b_data_out_clock = "clock1";
defparam ram_block1a34.port_b_data_width = 2;
defparam ram_block1a34.port_b_first_address = 0;
defparam ram_block1a34.port_b_first_bit_number = 34;
defparam ram_block1a34.port_b_last_address = 7;
defparam ram_block1a34.port_b_logical_ram_depth = 8;
defparam ram_block1a34.port_b_logical_ram_width = 128;
defparam ram_block1a34.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a34.port_b_read_enable_clock = "clock1";
defparam ram_block1a34.ram_block_type = "auto";

arriaii_ram_block ram_block1a35(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[35]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a35_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a35.clk0_core_clock_enable = "ena0";
defparam ram_block1a35.clk0_input_clock_enable = "ena2";
defparam ram_block1a35.clk1_core_clock_enable = "ena3";
defparam ram_block1a35.clk1_input_clock_enable = "ena3";
defparam ram_block1a35.clock_duty_cycle_dependence = "on";
defparam ram_block1a35.data_interleave_offset_in_bits = 64;
defparam ram_block1a35.data_interleave_width_in_bits = 1;
defparam ram_block1a35.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a35.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a35.operation_mode = "dual_port";
defparam ram_block1a35.port_a_address_clear = "none";
defparam ram_block1a35.port_a_address_width = 4;
defparam ram_block1a35.port_a_data_out_clear = "none";
defparam ram_block1a35.port_a_data_out_clock = "none";
defparam ram_block1a35.port_a_data_width = 1;
defparam ram_block1a35.port_a_first_address = 0;
defparam ram_block1a35.port_a_first_bit_number = 35;
defparam ram_block1a35.port_a_last_address = 15;
defparam ram_block1a35.port_a_logical_ram_depth = 16;
defparam ram_block1a35.port_a_logical_ram_width = 64;
defparam ram_block1a35.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a35.port_b_address_clear = "none";
defparam ram_block1a35.port_b_address_clock = "clock1";
defparam ram_block1a35.port_b_address_width = 3;
defparam ram_block1a35.port_b_data_out_clear = "none";
defparam ram_block1a35.port_b_data_out_clock = "clock1";
defparam ram_block1a35.port_b_data_width = 2;
defparam ram_block1a35.port_b_first_address = 0;
defparam ram_block1a35.port_b_first_bit_number = 35;
defparam ram_block1a35.port_b_last_address = 7;
defparam ram_block1a35.port_b_logical_ram_depth = 8;
defparam ram_block1a35.port_b_logical_ram_width = 128;
defparam ram_block1a35.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a35.port_b_read_enable_clock = "clock1";
defparam ram_block1a35.ram_block_type = "auto";

arriaii_ram_block ram_block1a36(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[36]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a36_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a36.clk0_core_clock_enable = "ena0";
defparam ram_block1a36.clk0_input_clock_enable = "ena2";
defparam ram_block1a36.clk1_core_clock_enable = "ena3";
defparam ram_block1a36.clk1_input_clock_enable = "ena3";
defparam ram_block1a36.clock_duty_cycle_dependence = "on";
defparam ram_block1a36.data_interleave_offset_in_bits = 64;
defparam ram_block1a36.data_interleave_width_in_bits = 1;
defparam ram_block1a36.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a36.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a36.operation_mode = "dual_port";
defparam ram_block1a36.port_a_address_clear = "none";
defparam ram_block1a36.port_a_address_width = 4;
defparam ram_block1a36.port_a_data_out_clear = "none";
defparam ram_block1a36.port_a_data_out_clock = "none";
defparam ram_block1a36.port_a_data_width = 1;
defparam ram_block1a36.port_a_first_address = 0;
defparam ram_block1a36.port_a_first_bit_number = 36;
defparam ram_block1a36.port_a_last_address = 15;
defparam ram_block1a36.port_a_logical_ram_depth = 16;
defparam ram_block1a36.port_a_logical_ram_width = 64;
defparam ram_block1a36.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a36.port_b_address_clear = "none";
defparam ram_block1a36.port_b_address_clock = "clock1";
defparam ram_block1a36.port_b_address_width = 3;
defparam ram_block1a36.port_b_data_out_clear = "none";
defparam ram_block1a36.port_b_data_out_clock = "clock1";
defparam ram_block1a36.port_b_data_width = 2;
defparam ram_block1a36.port_b_first_address = 0;
defparam ram_block1a36.port_b_first_bit_number = 36;
defparam ram_block1a36.port_b_last_address = 7;
defparam ram_block1a36.port_b_logical_ram_depth = 8;
defparam ram_block1a36.port_b_logical_ram_width = 128;
defparam ram_block1a36.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a36.port_b_read_enable_clock = "clock1";
defparam ram_block1a36.ram_block_type = "auto";

arriaii_ram_block ram_block1a37(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[37]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a37_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a37.clk0_core_clock_enable = "ena0";
defparam ram_block1a37.clk0_input_clock_enable = "ena2";
defparam ram_block1a37.clk1_core_clock_enable = "ena3";
defparam ram_block1a37.clk1_input_clock_enable = "ena3";
defparam ram_block1a37.clock_duty_cycle_dependence = "on";
defparam ram_block1a37.data_interleave_offset_in_bits = 64;
defparam ram_block1a37.data_interleave_width_in_bits = 1;
defparam ram_block1a37.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a37.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a37.operation_mode = "dual_port";
defparam ram_block1a37.port_a_address_clear = "none";
defparam ram_block1a37.port_a_address_width = 4;
defparam ram_block1a37.port_a_data_out_clear = "none";
defparam ram_block1a37.port_a_data_out_clock = "none";
defparam ram_block1a37.port_a_data_width = 1;
defparam ram_block1a37.port_a_first_address = 0;
defparam ram_block1a37.port_a_first_bit_number = 37;
defparam ram_block1a37.port_a_last_address = 15;
defparam ram_block1a37.port_a_logical_ram_depth = 16;
defparam ram_block1a37.port_a_logical_ram_width = 64;
defparam ram_block1a37.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a37.port_b_address_clear = "none";
defparam ram_block1a37.port_b_address_clock = "clock1";
defparam ram_block1a37.port_b_address_width = 3;
defparam ram_block1a37.port_b_data_out_clear = "none";
defparam ram_block1a37.port_b_data_out_clock = "clock1";
defparam ram_block1a37.port_b_data_width = 2;
defparam ram_block1a37.port_b_first_address = 0;
defparam ram_block1a37.port_b_first_bit_number = 37;
defparam ram_block1a37.port_b_last_address = 7;
defparam ram_block1a37.port_b_logical_ram_depth = 8;
defparam ram_block1a37.port_b_logical_ram_width = 128;
defparam ram_block1a37.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a37.port_b_read_enable_clock = "clock1";
defparam ram_block1a37.ram_block_type = "auto";

arriaii_ram_block ram_block1a38(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[38]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a38_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a38.clk0_core_clock_enable = "ena0";
defparam ram_block1a38.clk0_input_clock_enable = "ena2";
defparam ram_block1a38.clk1_core_clock_enable = "ena3";
defparam ram_block1a38.clk1_input_clock_enable = "ena3";
defparam ram_block1a38.clock_duty_cycle_dependence = "on";
defparam ram_block1a38.data_interleave_offset_in_bits = 64;
defparam ram_block1a38.data_interleave_width_in_bits = 1;
defparam ram_block1a38.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a38.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a38.operation_mode = "dual_port";
defparam ram_block1a38.port_a_address_clear = "none";
defparam ram_block1a38.port_a_address_width = 4;
defparam ram_block1a38.port_a_data_out_clear = "none";
defparam ram_block1a38.port_a_data_out_clock = "none";
defparam ram_block1a38.port_a_data_width = 1;
defparam ram_block1a38.port_a_first_address = 0;
defparam ram_block1a38.port_a_first_bit_number = 38;
defparam ram_block1a38.port_a_last_address = 15;
defparam ram_block1a38.port_a_logical_ram_depth = 16;
defparam ram_block1a38.port_a_logical_ram_width = 64;
defparam ram_block1a38.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a38.port_b_address_clear = "none";
defparam ram_block1a38.port_b_address_clock = "clock1";
defparam ram_block1a38.port_b_address_width = 3;
defparam ram_block1a38.port_b_data_out_clear = "none";
defparam ram_block1a38.port_b_data_out_clock = "clock1";
defparam ram_block1a38.port_b_data_width = 2;
defparam ram_block1a38.port_b_first_address = 0;
defparam ram_block1a38.port_b_first_bit_number = 38;
defparam ram_block1a38.port_b_last_address = 7;
defparam ram_block1a38.port_b_logical_ram_depth = 8;
defparam ram_block1a38.port_b_logical_ram_width = 128;
defparam ram_block1a38.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a38.port_b_read_enable_clock = "clock1";
defparam ram_block1a38.ram_block_type = "auto";

arriaii_ram_block ram_block1a39(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[39]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a39_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a39.clk0_core_clock_enable = "ena0";
defparam ram_block1a39.clk0_input_clock_enable = "ena2";
defparam ram_block1a39.clk1_core_clock_enable = "ena3";
defparam ram_block1a39.clk1_input_clock_enable = "ena3";
defparam ram_block1a39.clock_duty_cycle_dependence = "on";
defparam ram_block1a39.data_interleave_offset_in_bits = 64;
defparam ram_block1a39.data_interleave_width_in_bits = 1;
defparam ram_block1a39.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a39.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a39.operation_mode = "dual_port";
defparam ram_block1a39.port_a_address_clear = "none";
defparam ram_block1a39.port_a_address_width = 4;
defparam ram_block1a39.port_a_data_out_clear = "none";
defparam ram_block1a39.port_a_data_out_clock = "none";
defparam ram_block1a39.port_a_data_width = 1;
defparam ram_block1a39.port_a_first_address = 0;
defparam ram_block1a39.port_a_first_bit_number = 39;
defparam ram_block1a39.port_a_last_address = 15;
defparam ram_block1a39.port_a_logical_ram_depth = 16;
defparam ram_block1a39.port_a_logical_ram_width = 64;
defparam ram_block1a39.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a39.port_b_address_clear = "none";
defparam ram_block1a39.port_b_address_clock = "clock1";
defparam ram_block1a39.port_b_address_width = 3;
defparam ram_block1a39.port_b_data_out_clear = "none";
defparam ram_block1a39.port_b_data_out_clock = "clock1";
defparam ram_block1a39.port_b_data_width = 2;
defparam ram_block1a39.port_b_first_address = 0;
defparam ram_block1a39.port_b_first_bit_number = 39;
defparam ram_block1a39.port_b_last_address = 7;
defparam ram_block1a39.port_b_logical_ram_depth = 8;
defparam ram_block1a39.port_b_logical_ram_width = 128;
defparam ram_block1a39.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a39.port_b_read_enable_clock = "clock1";
defparam ram_block1a39.ram_block_type = "auto";

arriaii_ram_block ram_block1a48(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[48]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a48_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a48.clk0_core_clock_enable = "ena0";
defparam ram_block1a48.clk0_input_clock_enable = "ena2";
defparam ram_block1a48.clk1_core_clock_enable = "ena3";
defparam ram_block1a48.clk1_input_clock_enable = "ena3";
defparam ram_block1a48.clock_duty_cycle_dependence = "on";
defparam ram_block1a48.data_interleave_offset_in_bits = 64;
defparam ram_block1a48.data_interleave_width_in_bits = 1;
defparam ram_block1a48.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a48.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a48.operation_mode = "dual_port";
defparam ram_block1a48.port_a_address_clear = "none";
defparam ram_block1a48.port_a_address_width = 4;
defparam ram_block1a48.port_a_data_out_clear = "none";
defparam ram_block1a48.port_a_data_out_clock = "none";
defparam ram_block1a48.port_a_data_width = 1;
defparam ram_block1a48.port_a_first_address = 0;
defparam ram_block1a48.port_a_first_bit_number = 48;
defparam ram_block1a48.port_a_last_address = 15;
defparam ram_block1a48.port_a_logical_ram_depth = 16;
defparam ram_block1a48.port_a_logical_ram_width = 64;
defparam ram_block1a48.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a48.port_b_address_clear = "none";
defparam ram_block1a48.port_b_address_clock = "clock1";
defparam ram_block1a48.port_b_address_width = 3;
defparam ram_block1a48.port_b_data_out_clear = "none";
defparam ram_block1a48.port_b_data_out_clock = "clock1";
defparam ram_block1a48.port_b_data_width = 2;
defparam ram_block1a48.port_b_first_address = 0;
defparam ram_block1a48.port_b_first_bit_number = 48;
defparam ram_block1a48.port_b_last_address = 7;
defparam ram_block1a48.port_b_logical_ram_depth = 8;
defparam ram_block1a48.port_b_logical_ram_width = 128;
defparam ram_block1a48.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a48.port_b_read_enable_clock = "clock1";
defparam ram_block1a48.ram_block_type = "auto";

arriaii_ram_block ram_block1a49(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[49]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a49_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a49.clk0_core_clock_enable = "ena0";
defparam ram_block1a49.clk0_input_clock_enable = "ena2";
defparam ram_block1a49.clk1_core_clock_enable = "ena3";
defparam ram_block1a49.clk1_input_clock_enable = "ena3";
defparam ram_block1a49.clock_duty_cycle_dependence = "on";
defparam ram_block1a49.data_interleave_offset_in_bits = 64;
defparam ram_block1a49.data_interleave_width_in_bits = 1;
defparam ram_block1a49.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a49.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a49.operation_mode = "dual_port";
defparam ram_block1a49.port_a_address_clear = "none";
defparam ram_block1a49.port_a_address_width = 4;
defparam ram_block1a49.port_a_data_out_clear = "none";
defparam ram_block1a49.port_a_data_out_clock = "none";
defparam ram_block1a49.port_a_data_width = 1;
defparam ram_block1a49.port_a_first_address = 0;
defparam ram_block1a49.port_a_first_bit_number = 49;
defparam ram_block1a49.port_a_last_address = 15;
defparam ram_block1a49.port_a_logical_ram_depth = 16;
defparam ram_block1a49.port_a_logical_ram_width = 64;
defparam ram_block1a49.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a49.port_b_address_clear = "none";
defparam ram_block1a49.port_b_address_clock = "clock1";
defparam ram_block1a49.port_b_address_width = 3;
defparam ram_block1a49.port_b_data_out_clear = "none";
defparam ram_block1a49.port_b_data_out_clock = "clock1";
defparam ram_block1a49.port_b_data_width = 2;
defparam ram_block1a49.port_b_first_address = 0;
defparam ram_block1a49.port_b_first_bit_number = 49;
defparam ram_block1a49.port_b_last_address = 7;
defparam ram_block1a49.port_b_logical_ram_depth = 8;
defparam ram_block1a49.port_b_logical_ram_width = 128;
defparam ram_block1a49.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a49.port_b_read_enable_clock = "clock1";
defparam ram_block1a49.ram_block_type = "auto";

arriaii_ram_block ram_block1a50(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[50]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a50_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a50.clk0_core_clock_enable = "ena0";
defparam ram_block1a50.clk0_input_clock_enable = "ena2";
defparam ram_block1a50.clk1_core_clock_enable = "ena3";
defparam ram_block1a50.clk1_input_clock_enable = "ena3";
defparam ram_block1a50.clock_duty_cycle_dependence = "on";
defparam ram_block1a50.data_interleave_offset_in_bits = 64;
defparam ram_block1a50.data_interleave_width_in_bits = 1;
defparam ram_block1a50.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a50.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a50.operation_mode = "dual_port";
defparam ram_block1a50.port_a_address_clear = "none";
defparam ram_block1a50.port_a_address_width = 4;
defparam ram_block1a50.port_a_data_out_clear = "none";
defparam ram_block1a50.port_a_data_out_clock = "none";
defparam ram_block1a50.port_a_data_width = 1;
defparam ram_block1a50.port_a_first_address = 0;
defparam ram_block1a50.port_a_first_bit_number = 50;
defparam ram_block1a50.port_a_last_address = 15;
defparam ram_block1a50.port_a_logical_ram_depth = 16;
defparam ram_block1a50.port_a_logical_ram_width = 64;
defparam ram_block1a50.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a50.port_b_address_clear = "none";
defparam ram_block1a50.port_b_address_clock = "clock1";
defparam ram_block1a50.port_b_address_width = 3;
defparam ram_block1a50.port_b_data_out_clear = "none";
defparam ram_block1a50.port_b_data_out_clock = "clock1";
defparam ram_block1a50.port_b_data_width = 2;
defparam ram_block1a50.port_b_first_address = 0;
defparam ram_block1a50.port_b_first_bit_number = 50;
defparam ram_block1a50.port_b_last_address = 7;
defparam ram_block1a50.port_b_logical_ram_depth = 8;
defparam ram_block1a50.port_b_logical_ram_width = 128;
defparam ram_block1a50.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a50.port_b_read_enable_clock = "clock1";
defparam ram_block1a50.ram_block_type = "auto";

arriaii_ram_block ram_block1a51(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[51]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a51_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a51.clk0_core_clock_enable = "ena0";
defparam ram_block1a51.clk0_input_clock_enable = "ena2";
defparam ram_block1a51.clk1_core_clock_enable = "ena3";
defparam ram_block1a51.clk1_input_clock_enable = "ena3";
defparam ram_block1a51.clock_duty_cycle_dependence = "on";
defparam ram_block1a51.data_interleave_offset_in_bits = 64;
defparam ram_block1a51.data_interleave_width_in_bits = 1;
defparam ram_block1a51.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a51.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a51.operation_mode = "dual_port";
defparam ram_block1a51.port_a_address_clear = "none";
defparam ram_block1a51.port_a_address_width = 4;
defparam ram_block1a51.port_a_data_out_clear = "none";
defparam ram_block1a51.port_a_data_out_clock = "none";
defparam ram_block1a51.port_a_data_width = 1;
defparam ram_block1a51.port_a_first_address = 0;
defparam ram_block1a51.port_a_first_bit_number = 51;
defparam ram_block1a51.port_a_last_address = 15;
defparam ram_block1a51.port_a_logical_ram_depth = 16;
defparam ram_block1a51.port_a_logical_ram_width = 64;
defparam ram_block1a51.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a51.port_b_address_clear = "none";
defparam ram_block1a51.port_b_address_clock = "clock1";
defparam ram_block1a51.port_b_address_width = 3;
defparam ram_block1a51.port_b_data_out_clear = "none";
defparam ram_block1a51.port_b_data_out_clock = "clock1";
defparam ram_block1a51.port_b_data_width = 2;
defparam ram_block1a51.port_b_first_address = 0;
defparam ram_block1a51.port_b_first_bit_number = 51;
defparam ram_block1a51.port_b_last_address = 7;
defparam ram_block1a51.port_b_logical_ram_depth = 8;
defparam ram_block1a51.port_b_logical_ram_width = 128;
defparam ram_block1a51.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a51.port_b_read_enable_clock = "clock1";
defparam ram_block1a51.ram_block_type = "auto";

arriaii_ram_block ram_block1a52(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[52]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a52_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a52.clk0_core_clock_enable = "ena0";
defparam ram_block1a52.clk0_input_clock_enable = "ena2";
defparam ram_block1a52.clk1_core_clock_enable = "ena3";
defparam ram_block1a52.clk1_input_clock_enable = "ena3";
defparam ram_block1a52.clock_duty_cycle_dependence = "on";
defparam ram_block1a52.data_interleave_offset_in_bits = 64;
defparam ram_block1a52.data_interleave_width_in_bits = 1;
defparam ram_block1a52.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a52.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a52.operation_mode = "dual_port";
defparam ram_block1a52.port_a_address_clear = "none";
defparam ram_block1a52.port_a_address_width = 4;
defparam ram_block1a52.port_a_data_out_clear = "none";
defparam ram_block1a52.port_a_data_out_clock = "none";
defparam ram_block1a52.port_a_data_width = 1;
defparam ram_block1a52.port_a_first_address = 0;
defparam ram_block1a52.port_a_first_bit_number = 52;
defparam ram_block1a52.port_a_last_address = 15;
defparam ram_block1a52.port_a_logical_ram_depth = 16;
defparam ram_block1a52.port_a_logical_ram_width = 64;
defparam ram_block1a52.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a52.port_b_address_clear = "none";
defparam ram_block1a52.port_b_address_clock = "clock1";
defparam ram_block1a52.port_b_address_width = 3;
defparam ram_block1a52.port_b_data_out_clear = "none";
defparam ram_block1a52.port_b_data_out_clock = "clock1";
defparam ram_block1a52.port_b_data_width = 2;
defparam ram_block1a52.port_b_first_address = 0;
defparam ram_block1a52.port_b_first_bit_number = 52;
defparam ram_block1a52.port_b_last_address = 7;
defparam ram_block1a52.port_b_logical_ram_depth = 8;
defparam ram_block1a52.port_b_logical_ram_width = 128;
defparam ram_block1a52.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a52.port_b_read_enable_clock = "clock1";
defparam ram_block1a52.ram_block_type = "auto";

arriaii_ram_block ram_block1a53(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[53]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a53_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a53.clk0_core_clock_enable = "ena0";
defparam ram_block1a53.clk0_input_clock_enable = "ena2";
defparam ram_block1a53.clk1_core_clock_enable = "ena3";
defparam ram_block1a53.clk1_input_clock_enable = "ena3";
defparam ram_block1a53.clock_duty_cycle_dependence = "on";
defparam ram_block1a53.data_interleave_offset_in_bits = 64;
defparam ram_block1a53.data_interleave_width_in_bits = 1;
defparam ram_block1a53.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a53.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a53.operation_mode = "dual_port";
defparam ram_block1a53.port_a_address_clear = "none";
defparam ram_block1a53.port_a_address_width = 4;
defparam ram_block1a53.port_a_data_out_clear = "none";
defparam ram_block1a53.port_a_data_out_clock = "none";
defparam ram_block1a53.port_a_data_width = 1;
defparam ram_block1a53.port_a_first_address = 0;
defparam ram_block1a53.port_a_first_bit_number = 53;
defparam ram_block1a53.port_a_last_address = 15;
defparam ram_block1a53.port_a_logical_ram_depth = 16;
defparam ram_block1a53.port_a_logical_ram_width = 64;
defparam ram_block1a53.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a53.port_b_address_clear = "none";
defparam ram_block1a53.port_b_address_clock = "clock1";
defparam ram_block1a53.port_b_address_width = 3;
defparam ram_block1a53.port_b_data_out_clear = "none";
defparam ram_block1a53.port_b_data_out_clock = "clock1";
defparam ram_block1a53.port_b_data_width = 2;
defparam ram_block1a53.port_b_first_address = 0;
defparam ram_block1a53.port_b_first_bit_number = 53;
defparam ram_block1a53.port_b_last_address = 7;
defparam ram_block1a53.port_b_logical_ram_depth = 8;
defparam ram_block1a53.port_b_logical_ram_width = 128;
defparam ram_block1a53.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a53.port_b_read_enable_clock = "clock1";
defparam ram_block1a53.ram_block_type = "auto";

arriaii_ram_block ram_block1a54(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[54]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a54_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a54.clk0_core_clock_enable = "ena0";
defparam ram_block1a54.clk0_input_clock_enable = "ena2";
defparam ram_block1a54.clk1_core_clock_enable = "ena3";
defparam ram_block1a54.clk1_input_clock_enable = "ena3";
defparam ram_block1a54.clock_duty_cycle_dependence = "on";
defparam ram_block1a54.data_interleave_offset_in_bits = 64;
defparam ram_block1a54.data_interleave_width_in_bits = 1;
defparam ram_block1a54.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a54.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a54.operation_mode = "dual_port";
defparam ram_block1a54.port_a_address_clear = "none";
defparam ram_block1a54.port_a_address_width = 4;
defparam ram_block1a54.port_a_data_out_clear = "none";
defparam ram_block1a54.port_a_data_out_clock = "none";
defparam ram_block1a54.port_a_data_width = 1;
defparam ram_block1a54.port_a_first_address = 0;
defparam ram_block1a54.port_a_first_bit_number = 54;
defparam ram_block1a54.port_a_last_address = 15;
defparam ram_block1a54.port_a_logical_ram_depth = 16;
defparam ram_block1a54.port_a_logical_ram_width = 64;
defparam ram_block1a54.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a54.port_b_address_clear = "none";
defparam ram_block1a54.port_b_address_clock = "clock1";
defparam ram_block1a54.port_b_address_width = 3;
defparam ram_block1a54.port_b_data_out_clear = "none";
defparam ram_block1a54.port_b_data_out_clock = "clock1";
defparam ram_block1a54.port_b_data_width = 2;
defparam ram_block1a54.port_b_first_address = 0;
defparam ram_block1a54.port_b_first_bit_number = 54;
defparam ram_block1a54.port_b_last_address = 7;
defparam ram_block1a54.port_b_logical_ram_depth = 8;
defparam ram_block1a54.port_b_logical_ram_width = 128;
defparam ram_block1a54.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a54.port_b_read_enable_clock = "clock1";
defparam ram_block1a54.ram_block_type = "auto";

arriaii_ram_block ram_block1a55(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[55]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a55_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a55.clk0_core_clock_enable = "ena0";
defparam ram_block1a55.clk0_input_clock_enable = "ena2";
defparam ram_block1a55.clk1_core_clock_enable = "ena3";
defparam ram_block1a55.clk1_input_clock_enable = "ena3";
defparam ram_block1a55.clock_duty_cycle_dependence = "on";
defparam ram_block1a55.data_interleave_offset_in_bits = 64;
defparam ram_block1a55.data_interleave_width_in_bits = 1;
defparam ram_block1a55.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a55.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a55.operation_mode = "dual_port";
defparam ram_block1a55.port_a_address_clear = "none";
defparam ram_block1a55.port_a_address_width = 4;
defparam ram_block1a55.port_a_data_out_clear = "none";
defparam ram_block1a55.port_a_data_out_clock = "none";
defparam ram_block1a55.port_a_data_width = 1;
defparam ram_block1a55.port_a_first_address = 0;
defparam ram_block1a55.port_a_first_bit_number = 55;
defparam ram_block1a55.port_a_last_address = 15;
defparam ram_block1a55.port_a_logical_ram_depth = 16;
defparam ram_block1a55.port_a_logical_ram_width = 64;
defparam ram_block1a55.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a55.port_b_address_clear = "none";
defparam ram_block1a55.port_b_address_clock = "clock1";
defparam ram_block1a55.port_b_address_width = 3;
defparam ram_block1a55.port_b_data_out_clear = "none";
defparam ram_block1a55.port_b_data_out_clock = "clock1";
defparam ram_block1a55.port_b_data_width = 2;
defparam ram_block1a55.port_b_first_address = 0;
defparam ram_block1a55.port_b_first_bit_number = 55;
defparam ram_block1a55.port_b_last_address = 7;
defparam ram_block1a55.port_b_logical_ram_depth = 8;
defparam ram_block1a55.port_b_logical_ram_width = 128;
defparam ram_block1a55.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a55.port_b_read_enable_clock = "clock1";
defparam ram_block1a55.ram_block_type = "auto";

arriaii_ram_block ram_block1a8(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena2";
defparam ram_block1a8.clk1_core_clock_enable = "ena3";
defparam ram_block1a8.clk1_input_clock_enable = "ena3";
defparam ram_block1a8.clock_duty_cycle_dependence = "on";
defparam ram_block1a8.data_interleave_offset_in_bits = 64;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 4;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 15;
defparam ram_block1a8.port_a_logical_ram_depth = 16;
defparam ram_block1a8.port_a_logical_ram_width = 64;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 3;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "clock1";
defparam ram_block1a8.port_b_data_width = 2;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 7;
defparam ram_block1a8.port_b_logical_ram_depth = 8;
defparam ram_block1a8.port_b_logical_ram_width = 128;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

arriaii_ram_block ram_block1a9(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena2";
defparam ram_block1a9.clk1_core_clock_enable = "ena3";
defparam ram_block1a9.clk1_input_clock_enable = "ena3";
defparam ram_block1a9.clock_duty_cycle_dependence = "on";
defparam ram_block1a9.data_interleave_offset_in_bits = 64;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 4;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 15;
defparam ram_block1a9.port_a_logical_ram_depth = 16;
defparam ram_block1a9.port_a_logical_ram_width = 64;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 3;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "clock1";
defparam ram_block1a9.port_b_data_width = 2;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 7;
defparam ram_block1a9.port_b_logical_ram_depth = 8;
defparam ram_block1a9.port_b_logical_ram_width = 128;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

arriaii_ram_block ram_block1a10(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena2";
defparam ram_block1a10.clk1_core_clock_enable = "ena3";
defparam ram_block1a10.clk1_input_clock_enable = "ena3";
defparam ram_block1a10.clock_duty_cycle_dependence = "on";
defparam ram_block1a10.data_interleave_offset_in_bits = 64;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 4;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 15;
defparam ram_block1a10.port_a_logical_ram_depth = 16;
defparam ram_block1a10.port_a_logical_ram_width = 64;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 3;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "clock1";
defparam ram_block1a10.port_b_data_width = 2;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 7;
defparam ram_block1a10.port_b_logical_ram_depth = 8;
defparam ram_block1a10.port_b_logical_ram_width = 128;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

arriaii_ram_block ram_block1a11(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena2";
defparam ram_block1a11.clk1_core_clock_enable = "ena3";
defparam ram_block1a11.clk1_input_clock_enable = "ena3";
defparam ram_block1a11.clock_duty_cycle_dependence = "on";
defparam ram_block1a11.data_interleave_offset_in_bits = 64;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 4;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 15;
defparam ram_block1a11.port_a_logical_ram_depth = 16;
defparam ram_block1a11.port_a_logical_ram_width = 64;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 3;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "clock1";
defparam ram_block1a11.port_b_data_width = 2;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 7;
defparam ram_block1a11.port_b_logical_ram_depth = 8;
defparam ram_block1a11.port_b_logical_ram_width = 128;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

arriaii_ram_block ram_block1a12(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena2";
defparam ram_block1a12.clk1_core_clock_enable = "ena3";
defparam ram_block1a12.clk1_input_clock_enable = "ena3";
defparam ram_block1a12.clock_duty_cycle_dependence = "on";
defparam ram_block1a12.data_interleave_offset_in_bits = 64;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 4;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 15;
defparam ram_block1a12.port_a_logical_ram_depth = 16;
defparam ram_block1a12.port_a_logical_ram_width = 64;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 3;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "clock1";
defparam ram_block1a12.port_b_data_width = 2;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 7;
defparam ram_block1a12.port_b_logical_ram_depth = 8;
defparam ram_block1a12.port_b_logical_ram_width = 128;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

arriaii_ram_block ram_block1a13(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena2";
defparam ram_block1a13.clk1_core_clock_enable = "ena3";
defparam ram_block1a13.clk1_input_clock_enable = "ena3";
defparam ram_block1a13.clock_duty_cycle_dependence = "on";
defparam ram_block1a13.data_interleave_offset_in_bits = 64;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 4;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 15;
defparam ram_block1a13.port_a_logical_ram_depth = 16;
defparam ram_block1a13.port_a_logical_ram_width = 64;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 3;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "clock1";
defparam ram_block1a13.port_b_data_width = 2;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 7;
defparam ram_block1a13.port_b_logical_ram_depth = 8;
defparam ram_block1a13.port_b_logical_ram_width = 128;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

arriaii_ram_block ram_block1a14(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena2";
defparam ram_block1a14.clk1_core_clock_enable = "ena3";
defparam ram_block1a14.clk1_input_clock_enable = "ena3";
defparam ram_block1a14.clock_duty_cycle_dependence = "on";
defparam ram_block1a14.data_interleave_offset_in_bits = 64;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 4;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 15;
defparam ram_block1a14.port_a_logical_ram_depth = 16;
defparam ram_block1a14.port_a_logical_ram_width = 64;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 3;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "clock1";
defparam ram_block1a14.port_b_data_width = 2;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 7;
defparam ram_block1a14.port_b_logical_ram_depth = 8;
defparam ram_block1a14.port_b_logical_ram_width = 128;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

arriaii_ram_block ram_block1a15(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena2";
defparam ram_block1a15.clk1_core_clock_enable = "ena3";
defparam ram_block1a15.clk1_input_clock_enable = "ena3";
defparam ram_block1a15.clock_duty_cycle_dependence = "on";
defparam ram_block1a15.data_interleave_offset_in_bits = 64;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 4;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 15;
defparam ram_block1a15.port_a_logical_ram_depth = 16;
defparam ram_block1a15.port_a_logical_ram_width = 64;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 3;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "clock1";
defparam ram_block1a15.port_b_data_width = 2;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 7;
defparam ram_block1a15.port_b_logical_ram_depth = 8;
defparam ram_block1a15.port_b_logical_ram_width = 128;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

arriaii_ram_block ram_block1a24(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk0_input_clock_enable = "ena2";
defparam ram_block1a24.clk1_core_clock_enable = "ena3";
defparam ram_block1a24.clk1_input_clock_enable = "ena3";
defparam ram_block1a24.clock_duty_cycle_dependence = "on";
defparam ram_block1a24.data_interleave_offset_in_bits = 64;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 4;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 15;
defparam ram_block1a24.port_a_logical_ram_depth = 16;
defparam ram_block1a24.port_a_logical_ram_width = 64;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock1";
defparam ram_block1a24.port_b_address_width = 3;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "clock1";
defparam ram_block1a24.port_b_data_width = 2;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 7;
defparam ram_block1a24.port_b_logical_ram_depth = 8;
defparam ram_block1a24.port_b_logical_ram_width = 128;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock1";
defparam ram_block1a24.ram_block_type = "auto";

arriaii_ram_block ram_block1a25(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk0_input_clock_enable = "ena2";
defparam ram_block1a25.clk1_core_clock_enable = "ena3";
defparam ram_block1a25.clk1_input_clock_enable = "ena3";
defparam ram_block1a25.clock_duty_cycle_dependence = "on";
defparam ram_block1a25.data_interleave_offset_in_bits = 64;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 4;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 15;
defparam ram_block1a25.port_a_logical_ram_depth = 16;
defparam ram_block1a25.port_a_logical_ram_width = 64;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock1";
defparam ram_block1a25.port_b_address_width = 3;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "clock1";
defparam ram_block1a25.port_b_data_width = 2;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 7;
defparam ram_block1a25.port_b_logical_ram_depth = 8;
defparam ram_block1a25.port_b_logical_ram_width = 128;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock1";
defparam ram_block1a25.ram_block_type = "auto";

arriaii_ram_block ram_block1a26(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk0_input_clock_enable = "ena2";
defparam ram_block1a26.clk1_core_clock_enable = "ena3";
defparam ram_block1a26.clk1_input_clock_enable = "ena3";
defparam ram_block1a26.clock_duty_cycle_dependence = "on";
defparam ram_block1a26.data_interleave_offset_in_bits = 64;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 4;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 15;
defparam ram_block1a26.port_a_logical_ram_depth = 16;
defparam ram_block1a26.port_a_logical_ram_width = 64;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock1";
defparam ram_block1a26.port_b_address_width = 3;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "clock1";
defparam ram_block1a26.port_b_data_width = 2;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 7;
defparam ram_block1a26.port_b_logical_ram_depth = 8;
defparam ram_block1a26.port_b_logical_ram_width = 128;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock1";
defparam ram_block1a26.ram_block_type = "auto";

arriaii_ram_block ram_block1a27(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk0_input_clock_enable = "ena2";
defparam ram_block1a27.clk1_core_clock_enable = "ena3";
defparam ram_block1a27.clk1_input_clock_enable = "ena3";
defparam ram_block1a27.clock_duty_cycle_dependence = "on";
defparam ram_block1a27.data_interleave_offset_in_bits = 64;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 4;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 15;
defparam ram_block1a27.port_a_logical_ram_depth = 16;
defparam ram_block1a27.port_a_logical_ram_width = 64;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock1";
defparam ram_block1a27.port_b_address_width = 3;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "clock1";
defparam ram_block1a27.port_b_data_width = 2;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 7;
defparam ram_block1a27.port_b_logical_ram_depth = 8;
defparam ram_block1a27.port_b_logical_ram_width = 128;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock1";
defparam ram_block1a27.ram_block_type = "auto";

arriaii_ram_block ram_block1a28(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk0_input_clock_enable = "ena2";
defparam ram_block1a28.clk1_core_clock_enable = "ena3";
defparam ram_block1a28.clk1_input_clock_enable = "ena3";
defparam ram_block1a28.clock_duty_cycle_dependence = "on";
defparam ram_block1a28.data_interleave_offset_in_bits = 64;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 4;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 15;
defparam ram_block1a28.port_a_logical_ram_depth = 16;
defparam ram_block1a28.port_a_logical_ram_width = 64;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock1";
defparam ram_block1a28.port_b_address_width = 3;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "clock1";
defparam ram_block1a28.port_b_data_width = 2;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 7;
defparam ram_block1a28.port_b_logical_ram_depth = 8;
defparam ram_block1a28.port_b_logical_ram_width = 128;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock1";
defparam ram_block1a28.ram_block_type = "auto";

arriaii_ram_block ram_block1a29(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk0_input_clock_enable = "ena2";
defparam ram_block1a29.clk1_core_clock_enable = "ena3";
defparam ram_block1a29.clk1_input_clock_enable = "ena3";
defparam ram_block1a29.clock_duty_cycle_dependence = "on";
defparam ram_block1a29.data_interleave_offset_in_bits = 64;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 4;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 15;
defparam ram_block1a29.port_a_logical_ram_depth = 16;
defparam ram_block1a29.port_a_logical_ram_width = 64;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock1";
defparam ram_block1a29.port_b_address_width = 3;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "clock1";
defparam ram_block1a29.port_b_data_width = 2;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 7;
defparam ram_block1a29.port_b_logical_ram_depth = 8;
defparam ram_block1a29.port_b_logical_ram_width = 128;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock1";
defparam ram_block1a29.ram_block_type = "auto";

arriaii_ram_block ram_block1a30(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk0_input_clock_enable = "ena2";
defparam ram_block1a30.clk1_core_clock_enable = "ena3";
defparam ram_block1a30.clk1_input_clock_enable = "ena3";
defparam ram_block1a30.clock_duty_cycle_dependence = "on";
defparam ram_block1a30.data_interleave_offset_in_bits = 64;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 4;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 15;
defparam ram_block1a30.port_a_logical_ram_depth = 16;
defparam ram_block1a30.port_a_logical_ram_width = 64;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock1";
defparam ram_block1a30.port_b_address_width = 3;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "clock1";
defparam ram_block1a30.port_b_data_width = 2;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 7;
defparam ram_block1a30.port_b_logical_ram_depth = 8;
defparam ram_block1a30.port_b_logical_ram_width = 128;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock1";
defparam ram_block1a30.ram_block_type = "auto";

arriaii_ram_block ram_block1a31(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk0_input_clock_enable = "ena2";
defparam ram_block1a31.clk1_core_clock_enable = "ena3";
defparam ram_block1a31.clk1_input_clock_enable = "ena3";
defparam ram_block1a31.clock_duty_cycle_dependence = "on";
defparam ram_block1a31.data_interleave_offset_in_bits = 64;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 4;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 15;
defparam ram_block1a31.port_a_logical_ram_depth = 16;
defparam ram_block1a31.port_a_logical_ram_width = 64;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock1";
defparam ram_block1a31.port_b_address_width = 3;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "clock1";
defparam ram_block1a31.port_b_data_width = 2;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 7;
defparam ram_block1a31.port_b_logical_ram_depth = 8;
defparam ram_block1a31.port_b_logical_ram_width = 128;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock1";
defparam ram_block1a31.ram_block_type = "auto";

arriaii_ram_block ram_block1a40(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[40]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a40_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a40.clk0_core_clock_enable = "ena0";
defparam ram_block1a40.clk0_input_clock_enable = "ena2";
defparam ram_block1a40.clk1_core_clock_enable = "ena3";
defparam ram_block1a40.clk1_input_clock_enable = "ena3";
defparam ram_block1a40.clock_duty_cycle_dependence = "on";
defparam ram_block1a40.data_interleave_offset_in_bits = 64;
defparam ram_block1a40.data_interleave_width_in_bits = 1;
defparam ram_block1a40.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a40.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a40.operation_mode = "dual_port";
defparam ram_block1a40.port_a_address_clear = "none";
defparam ram_block1a40.port_a_address_width = 4;
defparam ram_block1a40.port_a_data_out_clear = "none";
defparam ram_block1a40.port_a_data_out_clock = "none";
defparam ram_block1a40.port_a_data_width = 1;
defparam ram_block1a40.port_a_first_address = 0;
defparam ram_block1a40.port_a_first_bit_number = 40;
defparam ram_block1a40.port_a_last_address = 15;
defparam ram_block1a40.port_a_logical_ram_depth = 16;
defparam ram_block1a40.port_a_logical_ram_width = 64;
defparam ram_block1a40.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a40.port_b_address_clear = "none";
defparam ram_block1a40.port_b_address_clock = "clock1";
defparam ram_block1a40.port_b_address_width = 3;
defparam ram_block1a40.port_b_data_out_clear = "none";
defparam ram_block1a40.port_b_data_out_clock = "clock1";
defparam ram_block1a40.port_b_data_width = 2;
defparam ram_block1a40.port_b_first_address = 0;
defparam ram_block1a40.port_b_first_bit_number = 40;
defparam ram_block1a40.port_b_last_address = 7;
defparam ram_block1a40.port_b_logical_ram_depth = 8;
defparam ram_block1a40.port_b_logical_ram_width = 128;
defparam ram_block1a40.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a40.port_b_read_enable_clock = "clock1";
defparam ram_block1a40.ram_block_type = "auto";

arriaii_ram_block ram_block1a41(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[41]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a41_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a41.clk0_core_clock_enable = "ena0";
defparam ram_block1a41.clk0_input_clock_enable = "ena2";
defparam ram_block1a41.clk1_core_clock_enable = "ena3";
defparam ram_block1a41.clk1_input_clock_enable = "ena3";
defparam ram_block1a41.clock_duty_cycle_dependence = "on";
defparam ram_block1a41.data_interleave_offset_in_bits = 64;
defparam ram_block1a41.data_interleave_width_in_bits = 1;
defparam ram_block1a41.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a41.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a41.operation_mode = "dual_port";
defparam ram_block1a41.port_a_address_clear = "none";
defparam ram_block1a41.port_a_address_width = 4;
defparam ram_block1a41.port_a_data_out_clear = "none";
defparam ram_block1a41.port_a_data_out_clock = "none";
defparam ram_block1a41.port_a_data_width = 1;
defparam ram_block1a41.port_a_first_address = 0;
defparam ram_block1a41.port_a_first_bit_number = 41;
defparam ram_block1a41.port_a_last_address = 15;
defparam ram_block1a41.port_a_logical_ram_depth = 16;
defparam ram_block1a41.port_a_logical_ram_width = 64;
defparam ram_block1a41.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a41.port_b_address_clear = "none";
defparam ram_block1a41.port_b_address_clock = "clock1";
defparam ram_block1a41.port_b_address_width = 3;
defparam ram_block1a41.port_b_data_out_clear = "none";
defparam ram_block1a41.port_b_data_out_clock = "clock1";
defparam ram_block1a41.port_b_data_width = 2;
defparam ram_block1a41.port_b_first_address = 0;
defparam ram_block1a41.port_b_first_bit_number = 41;
defparam ram_block1a41.port_b_last_address = 7;
defparam ram_block1a41.port_b_logical_ram_depth = 8;
defparam ram_block1a41.port_b_logical_ram_width = 128;
defparam ram_block1a41.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a41.port_b_read_enable_clock = "clock1";
defparam ram_block1a41.ram_block_type = "auto";

arriaii_ram_block ram_block1a42(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[42]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a42_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a42.clk0_core_clock_enable = "ena0";
defparam ram_block1a42.clk0_input_clock_enable = "ena2";
defparam ram_block1a42.clk1_core_clock_enable = "ena3";
defparam ram_block1a42.clk1_input_clock_enable = "ena3";
defparam ram_block1a42.clock_duty_cycle_dependence = "on";
defparam ram_block1a42.data_interleave_offset_in_bits = 64;
defparam ram_block1a42.data_interleave_width_in_bits = 1;
defparam ram_block1a42.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a42.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a42.operation_mode = "dual_port";
defparam ram_block1a42.port_a_address_clear = "none";
defparam ram_block1a42.port_a_address_width = 4;
defparam ram_block1a42.port_a_data_out_clear = "none";
defparam ram_block1a42.port_a_data_out_clock = "none";
defparam ram_block1a42.port_a_data_width = 1;
defparam ram_block1a42.port_a_first_address = 0;
defparam ram_block1a42.port_a_first_bit_number = 42;
defparam ram_block1a42.port_a_last_address = 15;
defparam ram_block1a42.port_a_logical_ram_depth = 16;
defparam ram_block1a42.port_a_logical_ram_width = 64;
defparam ram_block1a42.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a42.port_b_address_clear = "none";
defparam ram_block1a42.port_b_address_clock = "clock1";
defparam ram_block1a42.port_b_address_width = 3;
defparam ram_block1a42.port_b_data_out_clear = "none";
defparam ram_block1a42.port_b_data_out_clock = "clock1";
defparam ram_block1a42.port_b_data_width = 2;
defparam ram_block1a42.port_b_first_address = 0;
defparam ram_block1a42.port_b_first_bit_number = 42;
defparam ram_block1a42.port_b_last_address = 7;
defparam ram_block1a42.port_b_logical_ram_depth = 8;
defparam ram_block1a42.port_b_logical_ram_width = 128;
defparam ram_block1a42.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a42.port_b_read_enable_clock = "clock1";
defparam ram_block1a42.ram_block_type = "auto";

arriaii_ram_block ram_block1a43(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[43]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a43_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a43.clk0_core_clock_enable = "ena0";
defparam ram_block1a43.clk0_input_clock_enable = "ena2";
defparam ram_block1a43.clk1_core_clock_enable = "ena3";
defparam ram_block1a43.clk1_input_clock_enable = "ena3";
defparam ram_block1a43.clock_duty_cycle_dependence = "on";
defparam ram_block1a43.data_interleave_offset_in_bits = 64;
defparam ram_block1a43.data_interleave_width_in_bits = 1;
defparam ram_block1a43.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a43.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a43.operation_mode = "dual_port";
defparam ram_block1a43.port_a_address_clear = "none";
defparam ram_block1a43.port_a_address_width = 4;
defparam ram_block1a43.port_a_data_out_clear = "none";
defparam ram_block1a43.port_a_data_out_clock = "none";
defparam ram_block1a43.port_a_data_width = 1;
defparam ram_block1a43.port_a_first_address = 0;
defparam ram_block1a43.port_a_first_bit_number = 43;
defparam ram_block1a43.port_a_last_address = 15;
defparam ram_block1a43.port_a_logical_ram_depth = 16;
defparam ram_block1a43.port_a_logical_ram_width = 64;
defparam ram_block1a43.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a43.port_b_address_clear = "none";
defparam ram_block1a43.port_b_address_clock = "clock1";
defparam ram_block1a43.port_b_address_width = 3;
defparam ram_block1a43.port_b_data_out_clear = "none";
defparam ram_block1a43.port_b_data_out_clock = "clock1";
defparam ram_block1a43.port_b_data_width = 2;
defparam ram_block1a43.port_b_first_address = 0;
defparam ram_block1a43.port_b_first_bit_number = 43;
defparam ram_block1a43.port_b_last_address = 7;
defparam ram_block1a43.port_b_logical_ram_depth = 8;
defparam ram_block1a43.port_b_logical_ram_width = 128;
defparam ram_block1a43.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a43.port_b_read_enable_clock = "clock1";
defparam ram_block1a43.ram_block_type = "auto";

arriaii_ram_block ram_block1a44(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[44]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a44_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a44.clk0_core_clock_enable = "ena0";
defparam ram_block1a44.clk0_input_clock_enable = "ena2";
defparam ram_block1a44.clk1_core_clock_enable = "ena3";
defparam ram_block1a44.clk1_input_clock_enable = "ena3";
defparam ram_block1a44.clock_duty_cycle_dependence = "on";
defparam ram_block1a44.data_interleave_offset_in_bits = 64;
defparam ram_block1a44.data_interleave_width_in_bits = 1;
defparam ram_block1a44.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a44.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a44.operation_mode = "dual_port";
defparam ram_block1a44.port_a_address_clear = "none";
defparam ram_block1a44.port_a_address_width = 4;
defparam ram_block1a44.port_a_data_out_clear = "none";
defparam ram_block1a44.port_a_data_out_clock = "none";
defparam ram_block1a44.port_a_data_width = 1;
defparam ram_block1a44.port_a_first_address = 0;
defparam ram_block1a44.port_a_first_bit_number = 44;
defparam ram_block1a44.port_a_last_address = 15;
defparam ram_block1a44.port_a_logical_ram_depth = 16;
defparam ram_block1a44.port_a_logical_ram_width = 64;
defparam ram_block1a44.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a44.port_b_address_clear = "none";
defparam ram_block1a44.port_b_address_clock = "clock1";
defparam ram_block1a44.port_b_address_width = 3;
defparam ram_block1a44.port_b_data_out_clear = "none";
defparam ram_block1a44.port_b_data_out_clock = "clock1";
defparam ram_block1a44.port_b_data_width = 2;
defparam ram_block1a44.port_b_first_address = 0;
defparam ram_block1a44.port_b_first_bit_number = 44;
defparam ram_block1a44.port_b_last_address = 7;
defparam ram_block1a44.port_b_logical_ram_depth = 8;
defparam ram_block1a44.port_b_logical_ram_width = 128;
defparam ram_block1a44.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a44.port_b_read_enable_clock = "clock1";
defparam ram_block1a44.ram_block_type = "auto";

arriaii_ram_block ram_block1a45(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[45]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a45_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a45.clk0_core_clock_enable = "ena0";
defparam ram_block1a45.clk0_input_clock_enable = "ena2";
defparam ram_block1a45.clk1_core_clock_enable = "ena3";
defparam ram_block1a45.clk1_input_clock_enable = "ena3";
defparam ram_block1a45.clock_duty_cycle_dependence = "on";
defparam ram_block1a45.data_interleave_offset_in_bits = 64;
defparam ram_block1a45.data_interleave_width_in_bits = 1;
defparam ram_block1a45.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a45.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a45.operation_mode = "dual_port";
defparam ram_block1a45.port_a_address_clear = "none";
defparam ram_block1a45.port_a_address_width = 4;
defparam ram_block1a45.port_a_data_out_clear = "none";
defparam ram_block1a45.port_a_data_out_clock = "none";
defparam ram_block1a45.port_a_data_width = 1;
defparam ram_block1a45.port_a_first_address = 0;
defparam ram_block1a45.port_a_first_bit_number = 45;
defparam ram_block1a45.port_a_last_address = 15;
defparam ram_block1a45.port_a_logical_ram_depth = 16;
defparam ram_block1a45.port_a_logical_ram_width = 64;
defparam ram_block1a45.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a45.port_b_address_clear = "none";
defparam ram_block1a45.port_b_address_clock = "clock1";
defparam ram_block1a45.port_b_address_width = 3;
defparam ram_block1a45.port_b_data_out_clear = "none";
defparam ram_block1a45.port_b_data_out_clock = "clock1";
defparam ram_block1a45.port_b_data_width = 2;
defparam ram_block1a45.port_b_first_address = 0;
defparam ram_block1a45.port_b_first_bit_number = 45;
defparam ram_block1a45.port_b_last_address = 7;
defparam ram_block1a45.port_b_logical_ram_depth = 8;
defparam ram_block1a45.port_b_logical_ram_width = 128;
defparam ram_block1a45.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a45.port_b_read_enable_clock = "clock1";
defparam ram_block1a45.ram_block_type = "auto";

arriaii_ram_block ram_block1a46(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[46]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a46_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a46.clk0_core_clock_enable = "ena0";
defparam ram_block1a46.clk0_input_clock_enable = "ena2";
defparam ram_block1a46.clk1_core_clock_enable = "ena3";
defparam ram_block1a46.clk1_input_clock_enable = "ena3";
defparam ram_block1a46.clock_duty_cycle_dependence = "on";
defparam ram_block1a46.data_interleave_offset_in_bits = 64;
defparam ram_block1a46.data_interleave_width_in_bits = 1;
defparam ram_block1a46.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a46.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a46.operation_mode = "dual_port";
defparam ram_block1a46.port_a_address_clear = "none";
defparam ram_block1a46.port_a_address_width = 4;
defparam ram_block1a46.port_a_data_out_clear = "none";
defparam ram_block1a46.port_a_data_out_clock = "none";
defparam ram_block1a46.port_a_data_width = 1;
defparam ram_block1a46.port_a_first_address = 0;
defparam ram_block1a46.port_a_first_bit_number = 46;
defparam ram_block1a46.port_a_last_address = 15;
defparam ram_block1a46.port_a_logical_ram_depth = 16;
defparam ram_block1a46.port_a_logical_ram_width = 64;
defparam ram_block1a46.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a46.port_b_address_clear = "none";
defparam ram_block1a46.port_b_address_clock = "clock1";
defparam ram_block1a46.port_b_address_width = 3;
defparam ram_block1a46.port_b_data_out_clear = "none";
defparam ram_block1a46.port_b_data_out_clock = "clock1";
defparam ram_block1a46.port_b_data_width = 2;
defparam ram_block1a46.port_b_first_address = 0;
defparam ram_block1a46.port_b_first_bit_number = 46;
defparam ram_block1a46.port_b_last_address = 7;
defparam ram_block1a46.port_b_logical_ram_depth = 8;
defparam ram_block1a46.port_b_logical_ram_width = 128;
defparam ram_block1a46.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a46.port_b_read_enable_clock = "clock1";
defparam ram_block1a46.ram_block_type = "auto";

arriaii_ram_block ram_block1a47(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[47]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a47_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a47.clk0_core_clock_enable = "ena0";
defparam ram_block1a47.clk0_input_clock_enable = "ena2";
defparam ram_block1a47.clk1_core_clock_enable = "ena3";
defparam ram_block1a47.clk1_input_clock_enable = "ena3";
defparam ram_block1a47.clock_duty_cycle_dependence = "on";
defparam ram_block1a47.data_interleave_offset_in_bits = 64;
defparam ram_block1a47.data_interleave_width_in_bits = 1;
defparam ram_block1a47.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a47.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a47.operation_mode = "dual_port";
defparam ram_block1a47.port_a_address_clear = "none";
defparam ram_block1a47.port_a_address_width = 4;
defparam ram_block1a47.port_a_data_out_clear = "none";
defparam ram_block1a47.port_a_data_out_clock = "none";
defparam ram_block1a47.port_a_data_width = 1;
defparam ram_block1a47.port_a_first_address = 0;
defparam ram_block1a47.port_a_first_bit_number = 47;
defparam ram_block1a47.port_a_last_address = 15;
defparam ram_block1a47.port_a_logical_ram_depth = 16;
defparam ram_block1a47.port_a_logical_ram_width = 64;
defparam ram_block1a47.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a47.port_b_address_clear = "none";
defparam ram_block1a47.port_b_address_clock = "clock1";
defparam ram_block1a47.port_b_address_width = 3;
defparam ram_block1a47.port_b_data_out_clear = "none";
defparam ram_block1a47.port_b_data_out_clock = "clock1";
defparam ram_block1a47.port_b_data_width = 2;
defparam ram_block1a47.port_b_first_address = 0;
defparam ram_block1a47.port_b_first_bit_number = 47;
defparam ram_block1a47.port_b_last_address = 7;
defparam ram_block1a47.port_b_logical_ram_depth = 8;
defparam ram_block1a47.port_b_logical_ram_width = 128;
defparam ram_block1a47.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a47.port_b_read_enable_clock = "clock1";
defparam ram_block1a47.ram_block_type = "auto";

arriaii_ram_block ram_block1a56(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[56]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a56_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a56.clk0_core_clock_enable = "ena0";
defparam ram_block1a56.clk0_input_clock_enable = "ena2";
defparam ram_block1a56.clk1_core_clock_enable = "ena3";
defparam ram_block1a56.clk1_input_clock_enable = "ena3";
defparam ram_block1a56.clock_duty_cycle_dependence = "on";
defparam ram_block1a56.data_interleave_offset_in_bits = 64;
defparam ram_block1a56.data_interleave_width_in_bits = 1;
defparam ram_block1a56.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a56.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a56.operation_mode = "dual_port";
defparam ram_block1a56.port_a_address_clear = "none";
defparam ram_block1a56.port_a_address_width = 4;
defparam ram_block1a56.port_a_data_out_clear = "none";
defparam ram_block1a56.port_a_data_out_clock = "none";
defparam ram_block1a56.port_a_data_width = 1;
defparam ram_block1a56.port_a_first_address = 0;
defparam ram_block1a56.port_a_first_bit_number = 56;
defparam ram_block1a56.port_a_last_address = 15;
defparam ram_block1a56.port_a_logical_ram_depth = 16;
defparam ram_block1a56.port_a_logical_ram_width = 64;
defparam ram_block1a56.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a56.port_b_address_clear = "none";
defparam ram_block1a56.port_b_address_clock = "clock1";
defparam ram_block1a56.port_b_address_width = 3;
defparam ram_block1a56.port_b_data_out_clear = "none";
defparam ram_block1a56.port_b_data_out_clock = "clock1";
defparam ram_block1a56.port_b_data_width = 2;
defparam ram_block1a56.port_b_first_address = 0;
defparam ram_block1a56.port_b_first_bit_number = 56;
defparam ram_block1a56.port_b_last_address = 7;
defparam ram_block1a56.port_b_logical_ram_depth = 8;
defparam ram_block1a56.port_b_logical_ram_width = 128;
defparam ram_block1a56.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a56.port_b_read_enable_clock = "clock1";
defparam ram_block1a56.ram_block_type = "auto";

arriaii_ram_block ram_block1a57(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[57]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a57_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a57.clk0_core_clock_enable = "ena0";
defparam ram_block1a57.clk0_input_clock_enable = "ena2";
defparam ram_block1a57.clk1_core_clock_enable = "ena3";
defparam ram_block1a57.clk1_input_clock_enable = "ena3";
defparam ram_block1a57.clock_duty_cycle_dependence = "on";
defparam ram_block1a57.data_interleave_offset_in_bits = 64;
defparam ram_block1a57.data_interleave_width_in_bits = 1;
defparam ram_block1a57.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a57.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a57.operation_mode = "dual_port";
defparam ram_block1a57.port_a_address_clear = "none";
defparam ram_block1a57.port_a_address_width = 4;
defparam ram_block1a57.port_a_data_out_clear = "none";
defparam ram_block1a57.port_a_data_out_clock = "none";
defparam ram_block1a57.port_a_data_width = 1;
defparam ram_block1a57.port_a_first_address = 0;
defparam ram_block1a57.port_a_first_bit_number = 57;
defparam ram_block1a57.port_a_last_address = 15;
defparam ram_block1a57.port_a_logical_ram_depth = 16;
defparam ram_block1a57.port_a_logical_ram_width = 64;
defparam ram_block1a57.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a57.port_b_address_clear = "none";
defparam ram_block1a57.port_b_address_clock = "clock1";
defparam ram_block1a57.port_b_address_width = 3;
defparam ram_block1a57.port_b_data_out_clear = "none";
defparam ram_block1a57.port_b_data_out_clock = "clock1";
defparam ram_block1a57.port_b_data_width = 2;
defparam ram_block1a57.port_b_first_address = 0;
defparam ram_block1a57.port_b_first_bit_number = 57;
defparam ram_block1a57.port_b_last_address = 7;
defparam ram_block1a57.port_b_logical_ram_depth = 8;
defparam ram_block1a57.port_b_logical_ram_width = 128;
defparam ram_block1a57.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a57.port_b_read_enable_clock = "clock1";
defparam ram_block1a57.ram_block_type = "auto";

arriaii_ram_block ram_block1a58(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[58]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a58_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a58.clk0_core_clock_enable = "ena0";
defparam ram_block1a58.clk0_input_clock_enable = "ena2";
defparam ram_block1a58.clk1_core_clock_enable = "ena3";
defparam ram_block1a58.clk1_input_clock_enable = "ena3";
defparam ram_block1a58.clock_duty_cycle_dependence = "on";
defparam ram_block1a58.data_interleave_offset_in_bits = 64;
defparam ram_block1a58.data_interleave_width_in_bits = 1;
defparam ram_block1a58.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a58.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a58.operation_mode = "dual_port";
defparam ram_block1a58.port_a_address_clear = "none";
defparam ram_block1a58.port_a_address_width = 4;
defparam ram_block1a58.port_a_data_out_clear = "none";
defparam ram_block1a58.port_a_data_out_clock = "none";
defparam ram_block1a58.port_a_data_width = 1;
defparam ram_block1a58.port_a_first_address = 0;
defparam ram_block1a58.port_a_first_bit_number = 58;
defparam ram_block1a58.port_a_last_address = 15;
defparam ram_block1a58.port_a_logical_ram_depth = 16;
defparam ram_block1a58.port_a_logical_ram_width = 64;
defparam ram_block1a58.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a58.port_b_address_clear = "none";
defparam ram_block1a58.port_b_address_clock = "clock1";
defparam ram_block1a58.port_b_address_width = 3;
defparam ram_block1a58.port_b_data_out_clear = "none";
defparam ram_block1a58.port_b_data_out_clock = "clock1";
defparam ram_block1a58.port_b_data_width = 2;
defparam ram_block1a58.port_b_first_address = 0;
defparam ram_block1a58.port_b_first_bit_number = 58;
defparam ram_block1a58.port_b_last_address = 7;
defparam ram_block1a58.port_b_logical_ram_depth = 8;
defparam ram_block1a58.port_b_logical_ram_width = 128;
defparam ram_block1a58.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a58.port_b_read_enable_clock = "clock1";
defparam ram_block1a58.ram_block_type = "auto";

arriaii_ram_block ram_block1a59(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[59]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a59_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a59.clk0_core_clock_enable = "ena0";
defparam ram_block1a59.clk0_input_clock_enable = "ena2";
defparam ram_block1a59.clk1_core_clock_enable = "ena3";
defparam ram_block1a59.clk1_input_clock_enable = "ena3";
defparam ram_block1a59.clock_duty_cycle_dependence = "on";
defparam ram_block1a59.data_interleave_offset_in_bits = 64;
defparam ram_block1a59.data_interleave_width_in_bits = 1;
defparam ram_block1a59.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a59.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a59.operation_mode = "dual_port";
defparam ram_block1a59.port_a_address_clear = "none";
defparam ram_block1a59.port_a_address_width = 4;
defparam ram_block1a59.port_a_data_out_clear = "none";
defparam ram_block1a59.port_a_data_out_clock = "none";
defparam ram_block1a59.port_a_data_width = 1;
defparam ram_block1a59.port_a_first_address = 0;
defparam ram_block1a59.port_a_first_bit_number = 59;
defparam ram_block1a59.port_a_last_address = 15;
defparam ram_block1a59.port_a_logical_ram_depth = 16;
defparam ram_block1a59.port_a_logical_ram_width = 64;
defparam ram_block1a59.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a59.port_b_address_clear = "none";
defparam ram_block1a59.port_b_address_clock = "clock1";
defparam ram_block1a59.port_b_address_width = 3;
defparam ram_block1a59.port_b_data_out_clear = "none";
defparam ram_block1a59.port_b_data_out_clock = "clock1";
defparam ram_block1a59.port_b_data_width = 2;
defparam ram_block1a59.port_b_first_address = 0;
defparam ram_block1a59.port_b_first_bit_number = 59;
defparam ram_block1a59.port_b_last_address = 7;
defparam ram_block1a59.port_b_logical_ram_depth = 8;
defparam ram_block1a59.port_b_logical_ram_width = 128;
defparam ram_block1a59.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a59.port_b_read_enable_clock = "clock1";
defparam ram_block1a59.ram_block_type = "auto";

arriaii_ram_block ram_block1a60(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[60]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a60_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a60.clk0_core_clock_enable = "ena0";
defparam ram_block1a60.clk0_input_clock_enable = "ena2";
defparam ram_block1a60.clk1_core_clock_enable = "ena3";
defparam ram_block1a60.clk1_input_clock_enable = "ena3";
defparam ram_block1a60.clock_duty_cycle_dependence = "on";
defparam ram_block1a60.data_interleave_offset_in_bits = 64;
defparam ram_block1a60.data_interleave_width_in_bits = 1;
defparam ram_block1a60.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a60.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a60.operation_mode = "dual_port";
defparam ram_block1a60.port_a_address_clear = "none";
defparam ram_block1a60.port_a_address_width = 4;
defparam ram_block1a60.port_a_data_out_clear = "none";
defparam ram_block1a60.port_a_data_out_clock = "none";
defparam ram_block1a60.port_a_data_width = 1;
defparam ram_block1a60.port_a_first_address = 0;
defparam ram_block1a60.port_a_first_bit_number = 60;
defparam ram_block1a60.port_a_last_address = 15;
defparam ram_block1a60.port_a_logical_ram_depth = 16;
defparam ram_block1a60.port_a_logical_ram_width = 64;
defparam ram_block1a60.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a60.port_b_address_clear = "none";
defparam ram_block1a60.port_b_address_clock = "clock1";
defparam ram_block1a60.port_b_address_width = 3;
defparam ram_block1a60.port_b_data_out_clear = "none";
defparam ram_block1a60.port_b_data_out_clock = "clock1";
defparam ram_block1a60.port_b_data_width = 2;
defparam ram_block1a60.port_b_first_address = 0;
defparam ram_block1a60.port_b_first_bit_number = 60;
defparam ram_block1a60.port_b_last_address = 7;
defparam ram_block1a60.port_b_logical_ram_depth = 8;
defparam ram_block1a60.port_b_logical_ram_width = 128;
defparam ram_block1a60.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a60.port_b_read_enable_clock = "clock1";
defparam ram_block1a60.ram_block_type = "auto";

arriaii_ram_block ram_block1a61(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[61]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a61_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a61.clk0_core_clock_enable = "ena0";
defparam ram_block1a61.clk0_input_clock_enable = "ena2";
defparam ram_block1a61.clk1_core_clock_enable = "ena3";
defparam ram_block1a61.clk1_input_clock_enable = "ena3";
defparam ram_block1a61.clock_duty_cycle_dependence = "on";
defparam ram_block1a61.data_interleave_offset_in_bits = 64;
defparam ram_block1a61.data_interleave_width_in_bits = 1;
defparam ram_block1a61.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a61.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a61.operation_mode = "dual_port";
defparam ram_block1a61.port_a_address_clear = "none";
defparam ram_block1a61.port_a_address_width = 4;
defparam ram_block1a61.port_a_data_out_clear = "none";
defparam ram_block1a61.port_a_data_out_clock = "none";
defparam ram_block1a61.port_a_data_width = 1;
defparam ram_block1a61.port_a_first_address = 0;
defparam ram_block1a61.port_a_first_bit_number = 61;
defparam ram_block1a61.port_a_last_address = 15;
defparam ram_block1a61.port_a_logical_ram_depth = 16;
defparam ram_block1a61.port_a_logical_ram_width = 64;
defparam ram_block1a61.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a61.port_b_address_clear = "none";
defparam ram_block1a61.port_b_address_clock = "clock1";
defparam ram_block1a61.port_b_address_width = 3;
defparam ram_block1a61.port_b_data_out_clear = "none";
defparam ram_block1a61.port_b_data_out_clock = "clock1";
defparam ram_block1a61.port_b_data_width = 2;
defparam ram_block1a61.port_b_first_address = 0;
defparam ram_block1a61.port_b_first_bit_number = 61;
defparam ram_block1a61.port_b_last_address = 7;
defparam ram_block1a61.port_b_logical_ram_depth = 8;
defparam ram_block1a61.port_b_logical_ram_width = 128;
defparam ram_block1a61.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a61.port_b_read_enable_clock = "clock1";
defparam ram_block1a61.ram_block_type = "auto";

arriaii_ram_block ram_block1a62(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[62]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a62_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a62.clk0_core_clock_enable = "ena0";
defparam ram_block1a62.clk0_input_clock_enable = "ena2";
defparam ram_block1a62.clk1_core_clock_enable = "ena3";
defparam ram_block1a62.clk1_input_clock_enable = "ena3";
defparam ram_block1a62.clock_duty_cycle_dependence = "on";
defparam ram_block1a62.data_interleave_offset_in_bits = 64;
defparam ram_block1a62.data_interleave_width_in_bits = 1;
defparam ram_block1a62.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a62.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a62.operation_mode = "dual_port";
defparam ram_block1a62.port_a_address_clear = "none";
defparam ram_block1a62.port_a_address_width = 4;
defparam ram_block1a62.port_a_data_out_clear = "none";
defparam ram_block1a62.port_a_data_out_clock = "none";
defparam ram_block1a62.port_a_data_width = 1;
defparam ram_block1a62.port_a_first_address = 0;
defparam ram_block1a62.port_a_first_bit_number = 62;
defparam ram_block1a62.port_a_last_address = 15;
defparam ram_block1a62.port_a_logical_ram_depth = 16;
defparam ram_block1a62.port_a_logical_ram_width = 64;
defparam ram_block1a62.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a62.port_b_address_clear = "none";
defparam ram_block1a62.port_b_address_clock = "clock1";
defparam ram_block1a62.port_b_address_width = 3;
defparam ram_block1a62.port_b_data_out_clear = "none";
defparam ram_block1a62.port_b_data_out_clock = "clock1";
defparam ram_block1a62.port_b_data_width = 2;
defparam ram_block1a62.port_b_first_address = 0;
defparam ram_block1a62.port_b_first_bit_number = 62;
defparam ram_block1a62.port_b_last_address = 7;
defparam ram_block1a62.port_b_logical_ram_depth = 8;
defparam ram_block1a62.port_b_logical_ram_width = 128;
defparam ram_block1a62.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a62.port_b_read_enable_clock = "clock1";
defparam ram_block1a62.ram_block_type = "auto";

arriaii_ram_block ram_block1a63(
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[63]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(2'b00),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a63_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a63.clk0_core_clock_enable = "ena0";
defparam ram_block1a63.clk0_input_clock_enable = "ena2";
defparam ram_block1a63.clk1_core_clock_enable = "ena3";
defparam ram_block1a63.clk1_input_clock_enable = "ena3";
defparam ram_block1a63.clock_duty_cycle_dependence = "on";
defparam ram_block1a63.data_interleave_offset_in_bits = 64;
defparam ram_block1a63.data_interleave_width_in_bits = 1;
defparam ram_block1a63.logical_ram_name = "ddr3_int_controller_phy:ddr3_int_controller_phy_inst|ddr3_int_phy:ddr3_int_phy_inst|ddr3_int_phy_alt_mem_phy:ddr3_int_phy_alt_mem_phy_inst|ddr3_int_phy_alt_mem_phy_read_dp:rdp|altsyncram:half_rate_ram_gen.altsyncram_component|altsyncram_lbh1:auto_generated|ALTSYNCRAM";
defparam ram_block1a63.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a63.operation_mode = "dual_port";
defparam ram_block1a63.port_a_address_clear = "none";
defparam ram_block1a63.port_a_address_width = 4;
defparam ram_block1a63.port_a_data_out_clear = "none";
defparam ram_block1a63.port_a_data_out_clock = "none";
defparam ram_block1a63.port_a_data_width = 1;
defparam ram_block1a63.port_a_first_address = 0;
defparam ram_block1a63.port_a_first_bit_number = 63;
defparam ram_block1a63.port_a_last_address = 15;
defparam ram_block1a63.port_a_logical_ram_depth = 16;
defparam ram_block1a63.port_a_logical_ram_width = 64;
defparam ram_block1a63.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a63.port_b_address_clear = "none";
defparam ram_block1a63.port_b_address_clock = "clock1";
defparam ram_block1a63.port_b_address_width = 3;
defparam ram_block1a63.port_b_data_out_clear = "none";
defparam ram_block1a63.port_b_data_out_clock = "clock1";
defparam ram_block1a63.port_b_data_width = 2;
defparam ram_block1a63.port_b_first_address = 0;
defparam ram_block1a63.port_b_first_bit_number = 63;
defparam ram_block1a63.port_b_last_address = 7;
defparam ram_block1a63.port_b_logical_ram_depth = 8;
defparam ram_block1a63.port_b_logical_ram_width = 128;
defparam ram_block1a63.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a63.port_b_read_enable_clock = "clock1";
defparam ram_block1a63.ram_block_type = "auto";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_seq_wrapper (
	q_b_0,
	q_b_64,
	q_b_1,
	q_b_65,
	q_b_2,
	q_b_66,
	q_b_3,
	q_b_67,
	q_b_4,
	q_b_68,
	q_b_5,
	q_b_69,
	q_b_6,
	q_b_70,
	q_b_7,
	q_b_71,
	q_b_16,
	q_b_80,
	q_b_17,
	q_b_81,
	q_b_18,
	q_b_82,
	q_b_19,
	q_b_83,
	q_b_20,
	q_b_84,
	q_b_21,
	q_b_85,
	q_b_22,
	q_b_86,
	q_b_23,
	q_b_87,
	q_b_32,
	q_b_96,
	q_b_33,
	q_b_97,
	q_b_34,
	q_b_98,
	q_b_35,
	q_b_99,
	q_b_36,
	q_b_100,
	q_b_37,
	q_b_101,
	q_b_38,
	q_b_102,
	q_b_39,
	q_b_103,
	q_b_48,
	q_b_112,
	q_b_49,
	q_b_113,
	q_b_50,
	q_b_114,
	q_b_51,
	q_b_115,
	q_b_52,
	q_b_116,
	q_b_53,
	q_b_117,
	q_b_54,
	q_b_118,
	q_b_55,
	q_b_119,
	q_b_8,
	q_b_72,
	q_b_9,
	q_b_73,
	q_b_10,
	q_b_74,
	q_b_11,
	q_b_75,
	q_b_12,
	q_b_76,
	q_b_13,
	q_b_77,
	q_b_14,
	q_b_78,
	q_b_15,
	q_b_79,
	q_b_24,
	q_b_88,
	q_b_25,
	q_b_89,
	q_b_26,
	q_b_90,
	q_b_27,
	q_b_91,
	q_b_28,
	q_b_92,
	q_b_29,
	q_b_93,
	q_b_30,
	q_b_94,
	q_b_31,
	q_b_95,
	q_b_40,
	q_b_104,
	q_b_41,
	q_b_105,
	q_b_42,
	q_b_106,
	q_b_43,
	q_b_107,
	q_b_44,
	q_b_108,
	q_b_45,
	q_b_109,
	q_b_46,
	q_b_110,
	q_b_47,
	q_b_111,
	q_b_56,
	q_b_120,
	q_b_57,
	q_b_121,
	q_b_58,
	q_b_122,
	q_b_59,
	q_b_123,
	q_b_60,
	q_b_124,
	q_b_61,
	q_b_125,
	q_b_62,
	q_b_126,
	q_b_63,
	q_b_127,
	clk_0,
	seq_ac_cke_1,
	seq_ac_addr_0,
	seq_ac_addr_14,
	seq_ac_addr_1,
	seq_ac_addr_15,
	seq_ac_addr_16,
	seq_ac_addr_17,
	seq_ac_addr_18,
	seq_ac_addr_5,
	seq_ac_addr_19,
	seq_ac_addr_8,
	seq_ac_addr_22,
	seq_ac_addr_10,
	seq_ac_addr_24,
	seq_ac_addr_12,
	seq_ac_addr_26,
	seq_ac_ba_0,
	seq_ac_ba_3,
	seq_ac_ba_1,
	seq_ac_ba_4,
	seq_ac_rst_n_0,
	ctl_init_fail,
	ctl_init_success,
	reset_phy_clk_1x_n,
	ctl_init_fail1,
	ctl_init_success1,
	seq_rdv_doing_rd_7,
	seq_rdp_reset_req_n,
	seq_ac_add_1t_ac_lat_internal,
	wd_lat_2,
	wd_lat_1,
	wd_lat_0,
	wd_lat_3,
	wd_lat_4,
	seq_rdata_valid_lat_dec,
	seq_rdv_doing_rd_4,
	seq_pll_inc_dec_n,
	seq_pll_start_reconfig,
	seq_pll_select_2,
	seq_pll_select_1,
	seq_mem_clk_disable,
	seq_rdata_valid_0,
	seq_rdata_valid_1,
	seq_ac_cs_n_0,
	seq_ac_sel,
	dgwb_wdp_ovride,
	seq_wdp_ovride,
	dgwb_wdata_120,
	dgwb_wdata_56,
	dgwb_wdata_88,
	dgwb_wdata_24,
	dgwb_wdata_121,
	dgwb_wdata_57,
	dgwb_wdata_89,
	dgwb_wdata_25,
	dgwb_wdata_122,
	dgwb_wdata_58,
	dgwb_wdata_90,
	dgwb_wdata_26,
	dgwb_wdata_123,
	dgwb_wdata_59,
	dgwb_wdata_91,
	dgwb_wdata_27,
	dgwb_wdata_124,
	dgwb_wdata_60,
	dgwb_wdata_92,
	dgwb_wdata_28,
	dgwb_wdata_125,
	dgwb_wdata_61,
	dgwb_wdata_93,
	dgwb_wdata_29,
	dgwb_wdata_126,
	dgwb_wdata_62,
	dgwb_wdata_94,
	dgwb_wdata_30,
	dgwb_wdata_127,
	dgwb_wdata_63,
	dgwb_wdata_95,
	dgwb_wdata_31,
	seq_poa_protection_override_1x,
	seq_poa_lat_dec_1x_0,
	mimic_done_out,
	phs_shft_busy_siii,
	seq_mmc_start,
	mimic_value_captured,
	GND_port,
	dgwb_wdp_ovride1,
	seq_ac_cas_n_0,
	seq_ac_cas_n_1,
	seq_ac_cs_n_1,
	seq_ac_ras_n_0,
	seq_ac_ras_n_1,
	seq_ac_we_n_0,
	seq_ac_we_n_1)/* synthesis synthesis_greybox=0 */;
input 	q_b_0;
input 	q_b_64;
input 	q_b_1;
input 	q_b_65;
input 	q_b_2;
input 	q_b_66;
input 	q_b_3;
input 	q_b_67;
input 	q_b_4;
input 	q_b_68;
input 	q_b_5;
input 	q_b_69;
input 	q_b_6;
input 	q_b_70;
input 	q_b_7;
input 	q_b_71;
input 	q_b_16;
input 	q_b_80;
input 	q_b_17;
input 	q_b_81;
input 	q_b_18;
input 	q_b_82;
input 	q_b_19;
input 	q_b_83;
input 	q_b_20;
input 	q_b_84;
input 	q_b_21;
input 	q_b_85;
input 	q_b_22;
input 	q_b_86;
input 	q_b_23;
input 	q_b_87;
input 	q_b_32;
input 	q_b_96;
input 	q_b_33;
input 	q_b_97;
input 	q_b_34;
input 	q_b_98;
input 	q_b_35;
input 	q_b_99;
input 	q_b_36;
input 	q_b_100;
input 	q_b_37;
input 	q_b_101;
input 	q_b_38;
input 	q_b_102;
input 	q_b_39;
input 	q_b_103;
input 	q_b_48;
input 	q_b_112;
input 	q_b_49;
input 	q_b_113;
input 	q_b_50;
input 	q_b_114;
input 	q_b_51;
input 	q_b_115;
input 	q_b_52;
input 	q_b_116;
input 	q_b_53;
input 	q_b_117;
input 	q_b_54;
input 	q_b_118;
input 	q_b_55;
input 	q_b_119;
input 	q_b_8;
input 	q_b_72;
input 	q_b_9;
input 	q_b_73;
input 	q_b_10;
input 	q_b_74;
input 	q_b_11;
input 	q_b_75;
input 	q_b_12;
input 	q_b_76;
input 	q_b_13;
input 	q_b_77;
input 	q_b_14;
input 	q_b_78;
input 	q_b_15;
input 	q_b_79;
input 	q_b_24;
input 	q_b_88;
input 	q_b_25;
input 	q_b_89;
input 	q_b_26;
input 	q_b_90;
input 	q_b_27;
input 	q_b_91;
input 	q_b_28;
input 	q_b_92;
input 	q_b_29;
input 	q_b_93;
input 	q_b_30;
input 	q_b_94;
input 	q_b_31;
input 	q_b_95;
input 	q_b_40;
input 	q_b_104;
input 	q_b_41;
input 	q_b_105;
input 	q_b_42;
input 	q_b_106;
input 	q_b_43;
input 	q_b_107;
input 	q_b_44;
input 	q_b_108;
input 	q_b_45;
input 	q_b_109;
input 	q_b_46;
input 	q_b_110;
input 	q_b_47;
input 	q_b_111;
input 	q_b_56;
input 	q_b_120;
input 	q_b_57;
input 	q_b_121;
input 	q_b_58;
input 	q_b_122;
input 	q_b_59;
input 	q_b_123;
input 	q_b_60;
input 	q_b_124;
input 	q_b_61;
input 	q_b_125;
input 	q_b_62;
input 	q_b_126;
input 	q_b_63;
input 	q_b_127;
input 	clk_0;
output 	seq_ac_cke_1;
output 	seq_ac_addr_0;
output 	seq_ac_addr_14;
output 	seq_ac_addr_1;
output 	seq_ac_addr_15;
output 	seq_ac_addr_16;
output 	seq_ac_addr_17;
output 	seq_ac_addr_18;
output 	seq_ac_addr_5;
output 	seq_ac_addr_19;
output 	seq_ac_addr_8;
output 	seq_ac_addr_22;
output 	seq_ac_addr_10;
output 	seq_ac_addr_24;
output 	seq_ac_addr_12;
output 	seq_ac_addr_26;
output 	seq_ac_ba_0;
output 	seq_ac_ba_3;
output 	seq_ac_ba_1;
output 	seq_ac_ba_4;
output 	seq_ac_rst_n_0;
output 	ctl_init_fail;
output 	ctl_init_success;
input 	reset_phy_clk_1x_n;
output 	ctl_init_fail1;
output 	ctl_init_success1;
output 	seq_rdv_doing_rd_7;
output 	seq_rdp_reset_req_n;
output 	seq_ac_add_1t_ac_lat_internal;
output 	wd_lat_2;
output 	wd_lat_1;
output 	wd_lat_0;
output 	wd_lat_3;
output 	wd_lat_4;
output 	seq_rdata_valid_lat_dec;
output 	seq_rdv_doing_rd_4;
output 	seq_pll_inc_dec_n;
output 	seq_pll_start_reconfig;
output 	seq_pll_select_2;
output 	seq_pll_select_1;
output 	seq_mem_clk_disable;
input 	seq_rdata_valid_0;
input 	seq_rdata_valid_1;
output 	seq_ac_cs_n_0;
output 	seq_ac_sel;
output 	dgwb_wdp_ovride;
output 	seq_wdp_ovride;
output 	dgwb_wdata_120;
output 	dgwb_wdata_56;
output 	dgwb_wdata_88;
output 	dgwb_wdata_24;
output 	dgwb_wdata_121;
output 	dgwb_wdata_57;
output 	dgwb_wdata_89;
output 	dgwb_wdata_25;
output 	dgwb_wdata_122;
output 	dgwb_wdata_58;
output 	dgwb_wdata_90;
output 	dgwb_wdata_26;
output 	dgwb_wdata_123;
output 	dgwb_wdata_59;
output 	dgwb_wdata_91;
output 	dgwb_wdata_27;
output 	dgwb_wdata_124;
output 	dgwb_wdata_60;
output 	dgwb_wdata_92;
output 	dgwb_wdata_28;
output 	dgwb_wdata_125;
output 	dgwb_wdata_61;
output 	dgwb_wdata_93;
output 	dgwb_wdata_29;
output 	dgwb_wdata_126;
output 	dgwb_wdata_62;
output 	dgwb_wdata_94;
output 	dgwb_wdata_30;
output 	dgwb_wdata_127;
output 	dgwb_wdata_63;
output 	dgwb_wdata_95;
output 	dgwb_wdata_31;
output 	seq_poa_protection_override_1x;
output 	seq_poa_lat_dec_1x_0;
input 	mimic_done_out;
input 	phs_shft_busy_siii;
output 	seq_mmc_start;
input 	mimic_value_captured;
input 	GND_port;
output 	dgwb_wdp_ovride1;
output 	seq_ac_cas_n_0;
output 	seq_ac_cas_n_1;
output 	seq_ac_cs_n_1;
output 	seq_ac_ras_n_0;
output 	seq_ac_ras_n_1;
output 	seq_ac_we_n_0;
output 	seq_ac_we_n_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ddr3_int_ddr3_int_phy_alt_mem_phy_seq seq_inst(
	.q_b_0(q_b_0),
	.q_b_64(q_b_64),
	.q_b_1(q_b_1),
	.q_b_65(q_b_65),
	.q_b_2(q_b_2),
	.q_b_66(q_b_66),
	.q_b_3(q_b_3),
	.q_b_67(q_b_67),
	.q_b_4(q_b_4),
	.q_b_68(q_b_68),
	.q_b_5(q_b_5),
	.q_b_69(q_b_69),
	.q_b_6(q_b_6),
	.q_b_70(q_b_70),
	.q_b_7(q_b_7),
	.q_b_71(q_b_71),
	.q_b_16(q_b_16),
	.q_b_80(q_b_80),
	.q_b_17(q_b_17),
	.q_b_81(q_b_81),
	.q_b_18(q_b_18),
	.q_b_82(q_b_82),
	.q_b_19(q_b_19),
	.q_b_83(q_b_83),
	.q_b_20(q_b_20),
	.q_b_84(q_b_84),
	.q_b_21(q_b_21),
	.q_b_85(q_b_85),
	.q_b_22(q_b_22),
	.q_b_86(q_b_86),
	.q_b_23(q_b_23),
	.q_b_87(q_b_87),
	.q_b_32(q_b_32),
	.q_b_96(q_b_96),
	.q_b_33(q_b_33),
	.q_b_97(q_b_97),
	.q_b_34(q_b_34),
	.q_b_98(q_b_98),
	.q_b_35(q_b_35),
	.q_b_99(q_b_99),
	.q_b_36(q_b_36),
	.q_b_100(q_b_100),
	.q_b_37(q_b_37),
	.q_b_101(q_b_101),
	.q_b_38(q_b_38),
	.q_b_102(q_b_102),
	.q_b_39(q_b_39),
	.q_b_103(q_b_103),
	.q_b_48(q_b_48),
	.q_b_112(q_b_112),
	.q_b_49(q_b_49),
	.q_b_113(q_b_113),
	.q_b_50(q_b_50),
	.q_b_114(q_b_114),
	.q_b_51(q_b_51),
	.q_b_115(q_b_115),
	.q_b_52(q_b_52),
	.q_b_116(q_b_116),
	.q_b_53(q_b_53),
	.q_b_117(q_b_117),
	.q_b_54(q_b_54),
	.q_b_118(q_b_118),
	.q_b_55(q_b_55),
	.q_b_119(q_b_119),
	.q_b_8(q_b_8),
	.q_b_72(q_b_72),
	.q_b_9(q_b_9),
	.q_b_73(q_b_73),
	.q_b_10(q_b_10),
	.q_b_74(q_b_74),
	.q_b_11(q_b_11),
	.q_b_75(q_b_75),
	.q_b_12(q_b_12),
	.q_b_76(q_b_76),
	.q_b_13(q_b_13),
	.q_b_77(q_b_77),
	.q_b_14(q_b_14),
	.q_b_78(q_b_78),
	.q_b_15(q_b_15),
	.q_b_79(q_b_79),
	.q_b_24(q_b_24),
	.q_b_88(q_b_88),
	.q_b_25(q_b_25),
	.q_b_89(q_b_89),
	.q_b_26(q_b_26),
	.q_b_90(q_b_90),
	.q_b_27(q_b_27),
	.q_b_91(q_b_91),
	.q_b_28(q_b_28),
	.q_b_92(q_b_92),
	.q_b_29(q_b_29),
	.q_b_93(q_b_93),
	.q_b_30(q_b_30),
	.q_b_94(q_b_94),
	.q_b_31(q_b_31),
	.q_b_95(q_b_95),
	.q_b_40(q_b_40),
	.q_b_104(q_b_104),
	.q_b_41(q_b_41),
	.q_b_105(q_b_105),
	.q_b_42(q_b_42),
	.q_b_106(q_b_106),
	.q_b_43(q_b_43),
	.q_b_107(q_b_107),
	.q_b_44(q_b_44),
	.q_b_108(q_b_108),
	.q_b_45(q_b_45),
	.q_b_109(q_b_109),
	.q_b_46(q_b_46),
	.q_b_110(q_b_110),
	.q_b_47(q_b_47),
	.q_b_111(q_b_111),
	.q_b_56(q_b_56),
	.q_b_120(q_b_120),
	.q_b_57(q_b_57),
	.q_b_121(q_b_121),
	.q_b_58(q_b_58),
	.q_b_122(q_b_122),
	.q_b_59(q_b_59),
	.q_b_123(q_b_123),
	.q_b_60(q_b_60),
	.q_b_124(q_b_124),
	.q_b_61(q_b_61),
	.q_b_125(q_b_125),
	.q_b_62(q_b_62),
	.q_b_126(q_b_126),
	.q_b_63(q_b_63),
	.q_b_127(q_b_127),
	.clk(clk_0),
	.seq_ac_cke_1(seq_ac_cke_1),
	.seq_ac_addr_0(seq_ac_addr_0),
	.seq_ac_addr_14(seq_ac_addr_14),
	.seq_ac_addr_1(seq_ac_addr_1),
	.seq_ac_addr_15(seq_ac_addr_15),
	.seq_ac_addr_16(seq_ac_addr_16),
	.seq_ac_addr_17(seq_ac_addr_17),
	.seq_ac_addr_18(seq_ac_addr_18),
	.seq_ac_addr_5(seq_ac_addr_5),
	.seq_ac_addr_19(seq_ac_addr_19),
	.seq_ac_addr_8(seq_ac_addr_8),
	.seq_ac_addr_22(seq_ac_addr_22),
	.seq_ac_addr_10(seq_ac_addr_10),
	.seq_ac_addr_24(seq_ac_addr_24),
	.seq_ac_addr_12(seq_ac_addr_12),
	.seq_ac_addr_26(seq_ac_addr_26),
	.seq_ac_ba_0(seq_ac_ba_0),
	.seq_ac_ba_3(seq_ac_ba_3),
	.seq_ac_ba_1(seq_ac_ba_1),
	.seq_ac_ba_4(seq_ac_ba_4),
	.seq_ac_rst_n_0(seq_ac_rst_n_0),
	.ctl_init_fail1(ctl_init_fail),
	.ctl_init_success1(ctl_init_success),
	.rst_n(reset_phy_clk_1x_n),
	.ctl_init_fail2(ctl_init_fail1),
	.ctl_init_success2(ctl_init_success1),
	.seq_rdv_doing_rd_7(seq_rdv_doing_rd_7),
	.seq_rdp_reset_req_n1(seq_rdp_reset_req_n),
	.seq_ac_add_1t_ac_lat_internal1(seq_ac_add_1t_ac_lat_internal),
	.wd_lat_2(wd_lat_2),
	.wd_lat_1(wd_lat_1),
	.wd_lat_0(wd_lat_0),
	.wd_lat_3(wd_lat_3),
	.wd_lat_4(wd_lat_4),
	.seq_rdata_valid_lat_dec1(seq_rdata_valid_lat_dec),
	.seq_rdv_doing_rd_4(seq_rdv_doing_rd_4),
	.seq_pll_inc_dec_n1(seq_pll_inc_dec_n),
	.seq_pll_start_reconfig1(seq_pll_start_reconfig),
	.seq_pll_select_2(seq_pll_select_2),
	.seq_pll_select_1(seq_pll_select_1),
	.seq_mem_clk_disable1(seq_mem_clk_disable),
	.rdata_valid({gnd,seq_rdata_valid_0}),
	.seq_rdata_valid_1(seq_rdata_valid_1),
	.seq_ac_cs_n_0(seq_ac_cs_n_0),
	.seq_ac_sel(seq_ac_sel),
	.dgwb_wdp_ovride(dgwb_wdp_ovride),
	.seq_wdp_ovride(seq_wdp_ovride),
	.dgwb_wdata_120(dgwb_wdata_120),
	.dgwb_wdata_56(dgwb_wdata_56),
	.dgwb_wdata_88(dgwb_wdata_88),
	.dgwb_wdata_24(dgwb_wdata_24),
	.dgwb_wdata_121(dgwb_wdata_121),
	.dgwb_wdata_57(dgwb_wdata_57),
	.dgwb_wdata_89(dgwb_wdata_89),
	.dgwb_wdata_25(dgwb_wdata_25),
	.dgwb_wdata_122(dgwb_wdata_122),
	.dgwb_wdata_58(dgwb_wdata_58),
	.dgwb_wdata_90(dgwb_wdata_90),
	.dgwb_wdata_26(dgwb_wdata_26),
	.dgwb_wdata_123(dgwb_wdata_123),
	.dgwb_wdata_59(dgwb_wdata_59),
	.dgwb_wdata_91(dgwb_wdata_91),
	.dgwb_wdata_27(dgwb_wdata_27),
	.dgwb_wdata_124(dgwb_wdata_124),
	.dgwb_wdata_60(dgwb_wdata_60),
	.dgwb_wdata_92(dgwb_wdata_92),
	.dgwb_wdata_28(dgwb_wdata_28),
	.dgwb_wdata_125(dgwb_wdata_125),
	.dgwb_wdata_61(dgwb_wdata_61),
	.dgwb_wdata_93(dgwb_wdata_93),
	.dgwb_wdata_29(dgwb_wdata_29),
	.dgwb_wdata_126(dgwb_wdata_126),
	.dgwb_wdata_62(dgwb_wdata_62),
	.dgwb_wdata_94(dgwb_wdata_94),
	.dgwb_wdata_30(dgwb_wdata_30),
	.dgwb_wdata_127(dgwb_wdata_127),
	.dgwb_wdata_63(dgwb_wdata_63),
	.dgwb_wdata_95(dgwb_wdata_95),
	.dgwb_wdata_31(dgwb_wdata_31),
	.seq_poa_protection_override_1x1(seq_poa_protection_override_1x),
	.seq_poa_lat_dec_1x_0(seq_poa_lat_dec_1x_0),
	.mmc_seq_done(mimic_done_out),
	.seq_pll_phs_shift_busy(phs_shft_busy_siii),
	.seq_mmc_start(seq_mmc_start),
	.mmc_seq_value(mimic_value_captured),
	.GND_port(GND_port),
	.dgwb_wdp_ovride1(dgwb_wdp_ovride1),
	.seq_ac_cas_n_0(seq_ac_cas_n_0),
	.seq_ac_cas_n_1(seq_ac_cas_n_1),
	.seq_ac_cs_n_1(seq_ac_cs_n_1),
	.seq_ac_ras_n_0(seq_ac_ras_n_0),
	.seq_ac_ras_n_1(seq_ac_ras_n_1),
	.seq_ac_we_n_0(seq_ac_we_n_0),
	.seq_ac_we_n_1(seq_ac_we_n_1));

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_seq (
	q_b_0,
	q_b_64,
	q_b_1,
	q_b_65,
	q_b_2,
	q_b_66,
	q_b_3,
	q_b_67,
	q_b_4,
	q_b_68,
	q_b_5,
	q_b_69,
	q_b_6,
	q_b_70,
	q_b_7,
	q_b_71,
	q_b_16,
	q_b_80,
	q_b_17,
	q_b_81,
	q_b_18,
	q_b_82,
	q_b_19,
	q_b_83,
	q_b_20,
	q_b_84,
	q_b_21,
	q_b_85,
	q_b_22,
	q_b_86,
	q_b_23,
	q_b_87,
	q_b_32,
	q_b_96,
	q_b_33,
	q_b_97,
	q_b_34,
	q_b_98,
	q_b_35,
	q_b_99,
	q_b_36,
	q_b_100,
	q_b_37,
	q_b_101,
	q_b_38,
	q_b_102,
	q_b_39,
	q_b_103,
	q_b_48,
	q_b_112,
	q_b_49,
	q_b_113,
	q_b_50,
	q_b_114,
	q_b_51,
	q_b_115,
	q_b_52,
	q_b_116,
	q_b_53,
	q_b_117,
	q_b_54,
	q_b_118,
	q_b_55,
	q_b_119,
	q_b_8,
	q_b_72,
	q_b_9,
	q_b_73,
	q_b_10,
	q_b_74,
	q_b_11,
	q_b_75,
	q_b_12,
	q_b_76,
	q_b_13,
	q_b_77,
	q_b_14,
	q_b_78,
	q_b_15,
	q_b_79,
	q_b_24,
	q_b_88,
	q_b_25,
	q_b_89,
	q_b_26,
	q_b_90,
	q_b_27,
	q_b_91,
	q_b_28,
	q_b_92,
	q_b_29,
	q_b_93,
	q_b_30,
	q_b_94,
	q_b_31,
	q_b_95,
	q_b_40,
	q_b_104,
	q_b_41,
	q_b_105,
	q_b_42,
	q_b_106,
	q_b_43,
	q_b_107,
	q_b_44,
	q_b_108,
	q_b_45,
	q_b_109,
	q_b_46,
	q_b_110,
	q_b_47,
	q_b_111,
	q_b_56,
	q_b_120,
	q_b_57,
	q_b_121,
	q_b_58,
	q_b_122,
	q_b_59,
	q_b_123,
	q_b_60,
	q_b_124,
	q_b_61,
	q_b_125,
	q_b_62,
	q_b_126,
	q_b_63,
	q_b_127,
	clk,
	seq_ac_cke_1,
	seq_ac_addr_0,
	seq_ac_addr_14,
	seq_ac_addr_1,
	seq_ac_addr_15,
	seq_ac_addr_16,
	seq_ac_addr_17,
	seq_ac_addr_18,
	seq_ac_addr_5,
	seq_ac_addr_19,
	seq_ac_addr_8,
	seq_ac_addr_22,
	seq_ac_addr_10,
	seq_ac_addr_24,
	seq_ac_addr_12,
	seq_ac_addr_26,
	seq_ac_ba_0,
	seq_ac_ba_3,
	seq_ac_ba_1,
	seq_ac_ba_4,
	seq_ac_rst_n_0,
	ctl_init_fail1,
	ctl_init_success1,
	rst_n,
	ctl_init_fail2,
	ctl_init_success2,
	seq_rdv_doing_rd_7,
	seq_rdp_reset_req_n1,
	seq_ac_add_1t_ac_lat_internal1,
	wd_lat_2,
	wd_lat_1,
	wd_lat_0,
	wd_lat_3,
	wd_lat_4,
	seq_rdata_valid_lat_dec1,
	seq_rdv_doing_rd_4,
	seq_pll_inc_dec_n1,
	seq_pll_start_reconfig1,
	seq_pll_select_2,
	seq_pll_select_1,
	seq_mem_clk_disable1,
	rdata_valid,
	seq_rdata_valid_1,
	seq_ac_cs_n_0,
	seq_ac_sel,
	dgwb_wdp_ovride,
	seq_wdp_ovride,
	dgwb_wdata_120,
	dgwb_wdata_56,
	dgwb_wdata_88,
	dgwb_wdata_24,
	dgwb_wdata_121,
	dgwb_wdata_57,
	dgwb_wdata_89,
	dgwb_wdata_25,
	dgwb_wdata_122,
	dgwb_wdata_58,
	dgwb_wdata_90,
	dgwb_wdata_26,
	dgwb_wdata_123,
	dgwb_wdata_59,
	dgwb_wdata_91,
	dgwb_wdata_27,
	dgwb_wdata_124,
	dgwb_wdata_60,
	dgwb_wdata_92,
	dgwb_wdata_28,
	dgwb_wdata_125,
	dgwb_wdata_61,
	dgwb_wdata_93,
	dgwb_wdata_29,
	dgwb_wdata_126,
	dgwb_wdata_62,
	dgwb_wdata_94,
	dgwb_wdata_30,
	dgwb_wdata_127,
	dgwb_wdata_63,
	dgwb_wdata_95,
	dgwb_wdata_31,
	seq_poa_protection_override_1x1,
	seq_poa_lat_dec_1x_0,
	mmc_seq_done,
	seq_pll_phs_shift_busy,
	seq_mmc_start,
	mmc_seq_value,
	GND_port,
	dgwb_wdp_ovride1,
	seq_ac_cas_n_0,
	seq_ac_cas_n_1,
	seq_ac_cs_n_1,
	seq_ac_ras_n_0,
	seq_ac_ras_n_1,
	seq_ac_we_n_0,
	seq_ac_we_n_1)/* synthesis synthesis_greybox=0 */;
input 	q_b_0;
input 	q_b_64;
input 	q_b_1;
input 	q_b_65;
input 	q_b_2;
input 	q_b_66;
input 	q_b_3;
input 	q_b_67;
input 	q_b_4;
input 	q_b_68;
input 	q_b_5;
input 	q_b_69;
input 	q_b_6;
input 	q_b_70;
input 	q_b_7;
input 	q_b_71;
input 	q_b_16;
input 	q_b_80;
input 	q_b_17;
input 	q_b_81;
input 	q_b_18;
input 	q_b_82;
input 	q_b_19;
input 	q_b_83;
input 	q_b_20;
input 	q_b_84;
input 	q_b_21;
input 	q_b_85;
input 	q_b_22;
input 	q_b_86;
input 	q_b_23;
input 	q_b_87;
input 	q_b_32;
input 	q_b_96;
input 	q_b_33;
input 	q_b_97;
input 	q_b_34;
input 	q_b_98;
input 	q_b_35;
input 	q_b_99;
input 	q_b_36;
input 	q_b_100;
input 	q_b_37;
input 	q_b_101;
input 	q_b_38;
input 	q_b_102;
input 	q_b_39;
input 	q_b_103;
input 	q_b_48;
input 	q_b_112;
input 	q_b_49;
input 	q_b_113;
input 	q_b_50;
input 	q_b_114;
input 	q_b_51;
input 	q_b_115;
input 	q_b_52;
input 	q_b_116;
input 	q_b_53;
input 	q_b_117;
input 	q_b_54;
input 	q_b_118;
input 	q_b_55;
input 	q_b_119;
input 	q_b_8;
input 	q_b_72;
input 	q_b_9;
input 	q_b_73;
input 	q_b_10;
input 	q_b_74;
input 	q_b_11;
input 	q_b_75;
input 	q_b_12;
input 	q_b_76;
input 	q_b_13;
input 	q_b_77;
input 	q_b_14;
input 	q_b_78;
input 	q_b_15;
input 	q_b_79;
input 	q_b_24;
input 	q_b_88;
input 	q_b_25;
input 	q_b_89;
input 	q_b_26;
input 	q_b_90;
input 	q_b_27;
input 	q_b_91;
input 	q_b_28;
input 	q_b_92;
input 	q_b_29;
input 	q_b_93;
input 	q_b_30;
input 	q_b_94;
input 	q_b_31;
input 	q_b_95;
input 	q_b_40;
input 	q_b_104;
input 	q_b_41;
input 	q_b_105;
input 	q_b_42;
input 	q_b_106;
input 	q_b_43;
input 	q_b_107;
input 	q_b_44;
input 	q_b_108;
input 	q_b_45;
input 	q_b_109;
input 	q_b_46;
input 	q_b_110;
input 	q_b_47;
input 	q_b_111;
input 	q_b_56;
input 	q_b_120;
input 	q_b_57;
input 	q_b_121;
input 	q_b_58;
input 	q_b_122;
input 	q_b_59;
input 	q_b_123;
input 	q_b_60;
input 	q_b_124;
input 	q_b_61;
input 	q_b_125;
input 	q_b_62;
input 	q_b_126;
input 	q_b_63;
input 	q_b_127;
input 	clk;
output 	seq_ac_cke_1;
output 	seq_ac_addr_0;
output 	seq_ac_addr_14;
output 	seq_ac_addr_1;
output 	seq_ac_addr_15;
output 	seq_ac_addr_16;
output 	seq_ac_addr_17;
output 	seq_ac_addr_18;
output 	seq_ac_addr_5;
output 	seq_ac_addr_19;
output 	seq_ac_addr_8;
output 	seq_ac_addr_22;
output 	seq_ac_addr_10;
output 	seq_ac_addr_24;
output 	seq_ac_addr_12;
output 	seq_ac_addr_26;
output 	seq_ac_ba_0;
output 	seq_ac_ba_3;
output 	seq_ac_ba_1;
output 	seq_ac_ba_4;
output 	seq_ac_rst_n_0;
output 	ctl_init_fail1;
output 	ctl_init_success1;
input 	rst_n;
output 	ctl_init_fail2;
output 	ctl_init_success2;
output 	seq_rdv_doing_rd_7;
output 	seq_rdp_reset_req_n1;
output 	seq_ac_add_1t_ac_lat_internal1;
output 	wd_lat_2;
output 	wd_lat_1;
output 	wd_lat_0;
output 	wd_lat_3;
output 	wd_lat_4;
output 	seq_rdata_valid_lat_dec1;
output 	seq_rdv_doing_rd_4;
output 	seq_pll_inc_dec_n1;
output 	seq_pll_start_reconfig1;
output 	seq_pll_select_2;
output 	seq_pll_select_1;
output 	seq_mem_clk_disable1;
input 	[1:0] rdata_valid;
input 	seq_rdata_valid_1;
output 	seq_ac_cs_n_0;
output 	seq_ac_sel;
output 	dgwb_wdp_ovride;
output 	seq_wdp_ovride;
output 	dgwb_wdata_120;
output 	dgwb_wdata_56;
output 	dgwb_wdata_88;
output 	dgwb_wdata_24;
output 	dgwb_wdata_121;
output 	dgwb_wdata_57;
output 	dgwb_wdata_89;
output 	dgwb_wdata_25;
output 	dgwb_wdata_122;
output 	dgwb_wdata_58;
output 	dgwb_wdata_90;
output 	dgwb_wdata_26;
output 	dgwb_wdata_123;
output 	dgwb_wdata_59;
output 	dgwb_wdata_91;
output 	dgwb_wdata_27;
output 	dgwb_wdata_124;
output 	dgwb_wdata_60;
output 	dgwb_wdata_92;
output 	dgwb_wdata_28;
output 	dgwb_wdata_125;
output 	dgwb_wdata_61;
output 	dgwb_wdata_93;
output 	dgwb_wdata_29;
output 	dgwb_wdata_126;
output 	dgwb_wdata_62;
output 	dgwb_wdata_94;
output 	dgwb_wdata_30;
output 	dgwb_wdata_127;
output 	dgwb_wdata_63;
output 	dgwb_wdata_95;
output 	dgwb_wdata_31;
output 	seq_poa_protection_override_1x1;
output 	seq_poa_lat_dec_1x_0;
input 	mmc_seq_done;
input 	seq_pll_phs_shift_busy;
output 	seq_mmc_start;
input 	mmc_seq_value;
input 	GND_port;
output 	dgwb_wdp_ovride1;
output 	seq_ac_cas_n_0;
output 	seq_ac_cas_n_1;
output 	seq_ac_cs_n_1;
output 	seq_ac_ras_n_0;
output 	seq_ac_ras_n_1;
output 	seq_ac_we_n_0;
output 	seq_ac_we_n_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \dgwb|sig_addr_cmd[0].addr[2]~q ;
wire \dgwb|sig_addr_cmd[0].addr[3]~q ;
wire \dgwb|sig_addr_cmd[0].addr[4]~q ;
wire \dgwb|sig_addr_cmd[0].addr[5]~q ;
wire \dgwb|sig_addr_cmd[0].cas_n~q ;
wire \dgrb|sig_doing_rd[0]~q ;
wire \ctrl|state.s_rrp_sweep~q ;
wire \ctrl|state.s_rdv~q ;
wire \ctrl|state.s_rrp_seek~q ;
wire \ctrl|state.s_was~q ;
wire \ctrl|state.s_adv_wr_lat~q ;
wire \ctrl|state.s_adv_rd_lat~q ;
wire \ctrl|state.s_prep_customer_mr_setup~q ;
wire \ctrl|master_ctrl_op_rec~0_combout ;
wire \ctrl|ac_nt[0]~q ;
wire \dgrb|seq_rdata_valid_lat_dec~q ;
wire \dgrb|sig_doing_rd[4]~q ;
wire \dgb_ac_access_gnt_r~q ;
wire \dgrb|dgrb_ctrl_ac_nt_good~q ;
wire \dgrb|seq_pll_inc_dec_n~q ;
wire \ctrl|Selector61~0_combout ;
wire \ctrl|WideOr35~0_combout ;
wire \dgrb|seq_pll_start_reconfig~q ;
wire \dgrb|dgrb_ctrl.command_done~q ;
wire \ctrl|curr_cmd.cmd_was~q ;
wire \ctrl|curr_cmd.cmd_write_btp~q ;
wire \ctrl|curr_cmd.cmd_write_mtp~q ;
wire \ctrl|curr_ctrl.command_ack~0_combout ;
wire \ctrl|curr_cmd.cmd_idle~q ;
wire \ctrl|curr_cmd.cmd_prep_customer_mr_setup~q ;
wire \ctrl|curr_cmd.cmd_init_dram~q ;
wire \ctrl|curr_cmd.cmd_prog_cal_mr~q ;
wire \ctrl|WideOr0~0_combout ;
wire \dgwb|dgwb_ctrl.command_done~q ;
wire \admin|admin_ctrl.command_done~q ;
wire \admin|ac_access_gnt~q ;
wire \dgrb|dgrb_ctrl.command_err~q ;
wire \dgrb|seq_pll_select[0]~q ;
wire \dgrb|seq_pll_select[1]~q ;
wire \ctrl|WideOr2~combout ;
wire \ctrl|Selector61~1_combout ;
wire \dgwb|sig_addr_cmd[0].cke[0]~q ;
wire \dgrb|dgrb_ac_access_req~q ;
wire \dgwb|dgwb_ac_access_req~q ;
wire \admin|addr_cmd[0].cs_n[0]~q ;
wire \seq_ac_ras_n[1]~0_combout ;
wire \dgwb|sig_addr_cmd[1].cs_n[0]~q ;
wire \dgrb|sig_addr_cmd[1].cs_n[0]~q ;
wire \admin|addr_cmd[1].cs_n[0]~q ;
wire \admin|addr_cmd[0].cke[0]~q ;
wire \admin|addr_cmd[0].addr[0]~q ;
wire \admin|addr_cmd[1].addr[0]~q ;
wire \admin|addr_cmd[0].addr[1]~q ;
wire \admin|addr_cmd[1].addr[1]~q ;
wire \dgrb|sig_addr_cmd[0].addr[3]~q ;
wire \dgrb|sig_addr_cmd[0].addr[4]~q ;
wire \dgrb|sig_addr_cmd[0].addr[5]~q ;
wire \admin|addr_cmd[0].addr[8]~q ;
wire \admin|addr_cmd[1].addr[8]~q ;
wire \admin|addr_cmd[0].addr[10]~q ;
wire \admin|addr_cmd[1].addr[10]~q ;
wire \dgwb|sig_addr_cmd[0].addr[12]~q ;
wire \dgrb|sig_addr_cmd[0].addr[12]~q ;
wire \admin|addr_cmd[0].ba[0]~q ;
wire \admin|addr_cmd[1].ba[0]~q ;
wire \admin|addr_cmd[0].ba[1]~q ;
wire \admin|addr_cmd[1].ba[1]~q ;
wire \admin|addr_cmd[0].ras_n~q ;
wire \admin|addr_cmd[1].ras_n~q ;
wire \admin|addr_cmd[0].cas_n~q ;
wire \admin|addr_cmd[1].cas_n~q ;
wire \admin|addr_cmd[0].we_n~q ;
wire \admin|addr_cmd[1].we_n~q ;
wire \dgwb|sig_addr_cmd[0].rst_n~q ;
wire \admin|addr_cmd[0].rst_n~q ;
wire \ctrl|master_ctrl_op_rec~7_combout ;
wire \ctrl|master_ctrl_op_rec~8_combout ;
wire \dgb_ac_access_req~0_combout ;
wire \ctrl|master_ctrl_op_rec~9_combout ;
wire \dgrb|dgrb_ctrl.command_ack~q ;
wire \dgwb|dgwb_ctrl.command_ack~q ;
wire \admin|admin_ctrl.command_ack~q ;
wire \ctrl|master_ctrl_op_rec~10_combout ;
wire \ctrl|master_ctrl_op_rec~11_combout ;
wire \ctrl|master_ctrl_op_rec~12_combout ;
wire \ctrl|Selector60~0_combout ;
wire \ctrl|master_ctrl_op_rec~13_combout ;
wire \ctrl|master_ctrl_op_rec~14_combout ;
wire \dgrb_phs_shft_busy~q ;
wire \ctrl|ctrl_op_rec.command_op.mtp_almt~0_combout ;
wire \seq_pll_phs_shift_busy_ccd~q ;
wire \dgrb_phs_shft_busy~0_combout ;
wire \dgrb|seq_poa_lat_dec_1x[0]~q ;
wire \ctrl|ctrl_op_rec.command_op.single_bit~0_combout ;
wire \seq_pll_phs_shift_busy_r~q ;
wire \dgrb|dgrb_ctrl.command_result[5]~q ;
wire \dgrb|dgrb_ctrl.command_result[2]~q ;
wire \dgrb|dgrb_ctrl.command_result[1]~q ;
wire \dgrb|dgrb_ctrl.command_result[0]~q ;
wire \dgrb|dgrb_ctrl.command_result[3]~q ;
wire \dgrb|dgrb_ctrl.command_result[4]~q ;
wire \seq_ac_cke~0_combout ;
wire \ac_mux:ctrl_broadcast_r.command_req~q ;
wire \ac_mux:mem_clk_disable[0]~0_combout ;
wire \ac_mux:mem_clk_disable[0]~q ;
wire \seq_ac_addr~0_combout ;
wire \seq_ac_addr~1_combout ;
wire \seq_ac_addr~2_combout ;
wire \seq_ac_addr~3_combout ;
wire \seq_ac_addr~4_combout ;
wire \seq_ac_addr~5_combout ;
wire \seq_ac_addr~6_combout ;
wire \process_4~1_combout ;
wire \process_4~2_combout ;
wire \seq_ac_addr~7_combout ;
wire \seq_ac_addr~8_combout ;
wire \seq_ac_addr~9_combout ;
wire \seq_ac_addr~10_combout ;
wire \seq_ac_addr~11_combout ;
wire \seq_ac_addr~12_combout ;
wire \seq_ac_addr~13_combout ;
wire \seq_ac_addr~14_combout ;
wire \seq_ac_ba~0_combout ;
wire \seq_ac_ba~1_combout ;
wire \seq_ac_ba~2_combout ;
wire \seq_ac_ba~3_combout ;
wire \seq_ac_rst_n~0_combout ;
wire \seq_rdp_reset_req_n~0_combout ;
wire \seq_ac_add_1t_ac_lat_internal~0_combout ;
wire \seq_pll_inc_dec_n~0_combout ;
wire \seq_pll_start_reconfig~0_combout ;
wire \seq_pll_select~0_combout ;
wire \seq_pll_select~1_combout ;
wire \ac_mux:mem_clk_disable[1]~q ;
wire \ac_mux:mem_clk_disable[2]~q ;
wire \seq_ac_cs_n~0_combout ;
wire \WideNor0~combout ;
wire \seq_ac_ras_n[1]~1_combout ;
wire \seq_ac_cas_n~0_combout ;
wire \seq_ac_cas_n[0]~q ;
wire \seq_ac_cas_n~1_combout ;
wire \seq_ac_cas_n[1]~q ;
wire \seq_ac_cs_n~1_combout ;
wire \seq_ac_cs_n[1]~q ;
wire \seq_ac_ras_n~2_combout ;
wire \seq_ac_ras_n[0]~q ;
wire \seq_ac_ras_n~3_combout ;
wire \seq_ac_ras_n[1]~q ;
wire \seq_ac_we_n~0_combout ;
wire \seq_ac_we_n[0]~q ;
wire \seq_ac_we_n~1_combout ;
wire \seq_ac_we_n[1]~q ;


ddr3_int_ddr3_int_phy_alt_mem_phy_ctrl ctrl(
	.clk(clk),
	.rst_n(rst_n),
	.ctl_init_fail1(ctl_init_fail2),
	.ctl_init_success1(ctl_init_success2),
	.states_rrp_sweep(\ctrl|state.s_rrp_sweep~q ),
	.states_rdv(\ctrl|state.s_rdv~q ),
	.states_rrp_seek(\ctrl|state.s_rrp_seek~q ),
	.states_was(\ctrl|state.s_was~q ),
	.states_adv_wr_lat(\ctrl|state.s_adv_wr_lat~q ),
	.states_adv_rd_lat(\ctrl|state.s_adv_rd_lat~q ),
	.states_prep_customer_mr_setup(\ctrl|state.s_prep_customer_mr_setup~q ),
	.master_ctrl_op_rec(\ctrl|master_ctrl_op_rec~0_combout ),
	.ac_nt_0(\ctrl|ac_nt[0]~q ),
	.dgrb_ctrl_ac_nt_good(\dgrb|dgrb_ctrl_ac_nt_good~q ),
	.Selector61(\ctrl|Selector61~0_combout ),
	.WideOr35(\ctrl|WideOr35~0_combout ),
	.dgrb_ctrlcommand_done(\dgrb|dgrb_ctrl.command_done~q ),
	.curr_cmdcmd_was(\ctrl|curr_cmd.cmd_was~q ),
	.curr_cmdcmd_write_btp(\ctrl|curr_cmd.cmd_write_btp~q ),
	.curr_cmdcmd_write_mtp(\ctrl|curr_cmd.cmd_write_mtp~q ),
	.curr_ctrlcommand_ack(\ctrl|curr_ctrl.command_ack~0_combout ),
	.curr_cmdcmd_idle(\ctrl|curr_cmd.cmd_idle~q ),
	.curr_cmdcmd_prep_customer_mr_setup(\ctrl|curr_cmd.cmd_prep_customer_mr_setup~q ),
	.curr_cmdcmd_init_dram(\ctrl|curr_cmd.cmd_init_dram~q ),
	.curr_cmdcmd_prog_cal_mr(\ctrl|curr_cmd.cmd_prog_cal_mr~q ),
	.WideOr0(\ctrl|WideOr0~0_combout ),
	.dgwb_ctrlcommand_done(\dgwb|dgwb_ctrl.command_done~q ),
	.admin_ctrlcommand_done(\admin|admin_ctrl.command_done~q ),
	.dgrb_ctrlcommand_err(\dgrb|dgrb_ctrl.command_err~q ),
	.WideOr21(\ctrl|WideOr2~combout ),
	.Selector611(\ctrl|Selector61~1_combout ),
	.master_ctrl_op_rec1(\ctrl|master_ctrl_op_rec~7_combout ),
	.master_ctrl_op_rec2(\ctrl|master_ctrl_op_rec~8_combout ),
	.master_ctrl_op_rec3(\ctrl|master_ctrl_op_rec~9_combout ),
	.dgrb_ctrlcommand_ack(\dgrb|dgrb_ctrl.command_ack~q ),
	.dgwb_ctrlcommand_ack(\dgwb|dgwb_ctrl.command_ack~q ),
	.admin_ctrlcommand_ack(\admin|admin_ctrl.command_ack~q ),
	.master_ctrl_op_rec4(\ctrl|master_ctrl_op_rec~10_combout ),
	.master_ctrl_op_rec5(\ctrl|master_ctrl_op_rec~11_combout ),
	.master_ctrl_op_rec6(\ctrl|master_ctrl_op_rec~12_combout ),
	.Selector60(\ctrl|Selector60~0_combout ),
	.master_ctrl_op_rec7(\ctrl|master_ctrl_op_rec~13_combout ),
	.master_ctrl_op_rec8(\ctrl|master_ctrl_op_rec~14_combout ),
	.ctrl_op_reccommand_opmtp_almt(\ctrl|ctrl_op_rec.command_op.mtp_almt~0_combout ),
	.ctrl_op_reccommand_opsingle_bit(\ctrl|ctrl_op_rec.command_op.single_bit~0_combout ),
	.dgrb_ctrlcommand_result_5(\dgrb|dgrb_ctrl.command_result[5]~q ),
	.dgrb_ctrlcommand_result_2(\dgrb|dgrb_ctrl.command_result[2]~q ),
	.dgrb_ctrlcommand_result_1(\dgrb|dgrb_ctrl.command_result[1]~q ),
	.dgrb_ctrlcommand_result_0(\dgrb|dgrb_ctrl.command_result[0]~q ),
	.dgrb_ctrlcommand_result_3(\dgrb|dgrb_ctrl.command_result[3]~q ),
	.dgrb_ctrlcommand_result_4(\dgrb|dgrb_ctrl.command_result[4]~q ),
	.GND_port(GND_port));

ddr3_int_ddr3_int_phy_alt_mem_phy_dgrb dgrb(
	.q_b_0(q_b_0),
	.q_b_64(q_b_64),
	.q_b_1(q_b_1),
	.q_b_65(q_b_65),
	.q_b_2(q_b_2),
	.q_b_66(q_b_66),
	.q_b_3(q_b_3),
	.q_b_67(q_b_67),
	.q_b_4(q_b_4),
	.q_b_68(q_b_68),
	.q_b_5(q_b_5),
	.q_b_69(q_b_69),
	.q_b_6(q_b_6),
	.q_b_70(q_b_70),
	.q_b_7(q_b_7),
	.q_b_71(q_b_71),
	.q_b_16(q_b_16),
	.q_b_80(q_b_80),
	.q_b_17(q_b_17),
	.q_b_81(q_b_81),
	.q_b_18(q_b_18),
	.q_b_82(q_b_82),
	.q_b_19(q_b_19),
	.q_b_83(q_b_83),
	.q_b_20(q_b_20),
	.q_b_84(q_b_84),
	.q_b_21(q_b_21),
	.q_b_85(q_b_85),
	.q_b_22(q_b_22),
	.q_b_86(q_b_86),
	.q_b_23(q_b_23),
	.q_b_87(q_b_87),
	.q_b_32(q_b_32),
	.q_b_96(q_b_96),
	.q_b_33(q_b_33),
	.q_b_97(q_b_97),
	.q_b_34(q_b_34),
	.q_b_98(q_b_98),
	.q_b_35(q_b_35),
	.q_b_99(q_b_99),
	.q_b_36(q_b_36),
	.q_b_100(q_b_100),
	.q_b_37(q_b_37),
	.q_b_101(q_b_101),
	.q_b_38(q_b_38),
	.q_b_102(q_b_102),
	.q_b_39(q_b_39),
	.q_b_103(q_b_103),
	.q_b_48(q_b_48),
	.q_b_112(q_b_112),
	.q_b_49(q_b_49),
	.q_b_113(q_b_113),
	.q_b_50(q_b_50),
	.q_b_114(q_b_114),
	.q_b_51(q_b_51),
	.q_b_115(q_b_115),
	.q_b_52(q_b_52),
	.q_b_116(q_b_116),
	.q_b_53(q_b_53),
	.q_b_117(q_b_117),
	.q_b_54(q_b_54),
	.q_b_118(q_b_118),
	.q_b_55(q_b_55),
	.q_b_119(q_b_119),
	.q_b_8(q_b_8),
	.q_b_72(q_b_72),
	.q_b_9(q_b_9),
	.q_b_73(q_b_73),
	.q_b_10(q_b_10),
	.q_b_74(q_b_74),
	.q_b_11(q_b_11),
	.q_b_75(q_b_75),
	.q_b_12(q_b_12),
	.q_b_76(q_b_76),
	.q_b_13(q_b_13),
	.q_b_77(q_b_77),
	.q_b_14(q_b_14),
	.q_b_78(q_b_78),
	.q_b_15(q_b_15),
	.q_b_79(q_b_79),
	.q_b_24(q_b_24),
	.q_b_88(q_b_88),
	.q_b_25(q_b_25),
	.q_b_89(q_b_89),
	.q_b_26(q_b_26),
	.q_b_90(q_b_90),
	.q_b_27(q_b_27),
	.q_b_91(q_b_91),
	.q_b_28(q_b_28),
	.q_b_92(q_b_92),
	.q_b_29(q_b_29),
	.q_b_93(q_b_93),
	.q_b_30(q_b_30),
	.q_b_94(q_b_94),
	.q_b_31(q_b_31),
	.q_b_95(q_b_95),
	.q_b_40(q_b_40),
	.q_b_104(q_b_104),
	.q_b_41(q_b_41),
	.q_b_105(q_b_105),
	.q_b_42(q_b_42),
	.q_b_106(q_b_106),
	.q_b_43(q_b_43),
	.q_b_107(q_b_107),
	.q_b_44(q_b_44),
	.q_b_108(q_b_108),
	.q_b_45(q_b_45),
	.q_b_109(q_b_109),
	.q_b_46(q_b_46),
	.q_b_110(q_b_110),
	.q_b_47(q_b_47),
	.q_b_111(q_b_111),
	.q_b_56(q_b_56),
	.q_b_120(q_b_120),
	.q_b_57(q_b_57),
	.q_b_121(q_b_121),
	.q_b_58(q_b_58),
	.q_b_122(q_b_122),
	.q_b_59(q_b_59),
	.q_b_123(q_b_123),
	.q_b_60(q_b_60),
	.q_b_124(q_b_124),
	.q_b_61(q_b_61),
	.q_b_125(q_b_125),
	.q_b_62(q_b_62),
	.q_b_126(q_b_126),
	.q_b_63(q_b_63),
	.q_b_127(q_b_127),
	.clk(clk),
	.rst_n(rst_n),
	.wd_lat_2(wd_lat_2),
	.wd_lat_1(wd_lat_1),
	.wd_lat_0(wd_lat_0),
	.wd_lat_3(wd_lat_3),
	.wd_lat_4(wd_lat_4),
	.sig_doing_rd_0(\dgrb|sig_doing_rd[0]~q ),
	.seq_rdata_valid_lat_dec1(\dgrb|seq_rdata_valid_lat_dec~q ),
	.sig_doing_rd_4(\dgrb|sig_doing_rd[4]~q ),
	.dgb_ac_access_gnt_r(\dgb_ac_access_gnt_r~q ),
	.dgrb_ctrl_ac_nt_good1(\dgrb|dgrb_ctrl_ac_nt_good~q ),
	.seq_pll_inc_dec_n1(\dgrb|seq_pll_inc_dec_n~q ),
	.seq_pll_start_reconfig1(\dgrb|seq_pll_start_reconfig~q ),
	.dgrb_ctrlcommand_done(\dgrb|dgrb_ctrl.command_done~q ),
	.curr_ctrlcommand_ack(\ctrl|curr_ctrl.command_ack~0_combout ),
	.curr_cmdcmd_idle(\ctrl|curr_cmd.cmd_idle~q ),
	.WideOr0(\ctrl|WideOr0~0_combout ),
	.rdata_valid({gnd,rdata_valid[0]}),
	.seq_rdata_valid_1(seq_rdata_valid_1),
	.dgrb_ctrlcommand_err(\dgrb|dgrb_ctrl.command_err~q ),
	.seq_pll_select_0(\dgrb|seq_pll_select[0]~q ),
	.seq_pll_select_1(\dgrb|seq_pll_select[1]~q ),
	.WideOr2(\ctrl|WideOr2~combout ),
	.ac_muxctrl_broadcast_rcommand_req(\ac_mux:ctrl_broadcast_r.command_req~q ),
	.sig_addr_cmd0cke0(\dgwb|sig_addr_cmd[0].cke[0]~q ),
	.dgrb_ac_access_req1(\dgrb|dgrb_ac_access_req~q ),
	.sig_addr_cmd1cs_n0(\dgrb|sig_addr_cmd[1].cs_n[0]~q ),
	.sig_addr_cmd0addr3(\dgrb|sig_addr_cmd[0].addr[3]~q ),
	.sig_addr_cmd0addr4(\dgrb|sig_addr_cmd[0].addr[4]~q ),
	.sig_addr_cmd0addr5(\dgrb|sig_addr_cmd[0].addr[5]~q ),
	.sig_addr_cmd0addr12(\dgrb|sig_addr_cmd[0].addr[12]~q ),
	.\ctrl_dgrb.command.cmd_prep_adv_wr_lat (\ctrl|master_ctrl_op_rec~7_combout ),
	.\ctrl_dgrb.command.cmd_rdv (\ctrl|master_ctrl_op_rec~8_combout ),
	.\ctrl_dgrb.command.cmd_read_mtp (\ctrl|master_ctrl_op_rec~9_combout ),
	.dgrb_ctrlcommand_ack(\dgrb|dgrb_ctrl.command_ack~q ),
	.\ctrl_dgrb.command.cmd_rrp_seek (\ctrl|master_ctrl_op_rec~10_combout ),
	.\ctrl_dgrb.command.cmd_rrp_reset (\ctrl|master_ctrl_op_rec~11_combout ),
	.\ctrl_dgrb.command.cmd_rrp_sweep (\ctrl|master_ctrl_op_rec~12_combout ),
	.\ctrl_dgrb.command.cmd_tr_due (\ctrl|Selector60~0_combout ),
	.\ctrl_dgrb.command.cmd_poa (\ctrl|master_ctrl_op_rec~13_combout ),
	.\ctrl_dgrb.command.cmd_prep_adv_rd_lat (\ctrl|master_ctrl_op_rec~14_combout ),
	.phs_shft_busy(\dgrb_phs_shft_busy~q ),
	.\ctrl_dgrb.command_op.mtp_almt (\ctrl|ctrl_op_rec.command_op.mtp_almt~0_combout ),
	.mmc_seq_done(mmc_seq_done),
	.seq_poa_lat_dec_1x_0(\dgrb|seq_poa_lat_dec_1x[0]~q ),
	.\ctrl_dgrb.command_op.single_bit (\ctrl|ctrl_op_rec.command_op.single_bit~0_combout ),
	.dgrb_ctrlcommand_result_5(\dgrb|dgrb_ctrl.command_result[5]~q ),
	.dgrb_ctrlcommand_result_2(\dgrb|dgrb_ctrl.command_result[2]~q ),
	.dgrb_ctrlcommand_result_1(\dgrb|dgrb_ctrl.command_result[1]~q ),
	.dgrb_ctrlcommand_result_0(\dgrb|dgrb_ctrl.command_result[0]~q ),
	.dgrb_ctrlcommand_result_3(\dgrb|dgrb_ctrl.command_result[3]~q ),
	.dgrb_ctrlcommand_result_4(\dgrb|dgrb_ctrl.command_result[4]~q ),
	.seq_mmc_start1(seq_mmc_start),
	.mmc_seq_value(mmc_seq_value),
	.GND_port(GND_port));

ddr3_int_ddr3_int_phy_alt_mem_phy_dgwb dgwb(
	.clk(clk),
	.sig_addr_cmd0addr2(\dgwb|sig_addr_cmd[0].addr[2]~q ),
	.sig_addr_cmd0addr3(\dgwb|sig_addr_cmd[0].addr[3]~q ),
	.sig_addr_cmd0addr4(\dgwb|sig_addr_cmd[0].addr[4]~q ),
	.sig_addr_cmd0addr5(\dgwb|sig_addr_cmd[0].addr[5]~q ),
	.sig_addr_cmd0cas_n(\dgwb|sig_addr_cmd[0].cas_n~q ),
	.rst_n(rst_n),
	.dgb_ac_access_gnt_r(\dgb_ac_access_gnt_r~q ),
	.curr_cmdcmd_was(\ctrl|curr_cmd.cmd_was~q ),
	.curr_cmdcmd_write_btp(\ctrl|curr_cmd.cmd_write_btp~q ),
	.curr_cmdcmd_write_mtp(\ctrl|curr_cmd.cmd_write_mtp~q ),
	.curr_ctrlcommand_ack(\ctrl|curr_ctrl.command_ack~0_combout ),
	.dgwb_ctrlcommand_done(\dgwb|dgwb_ctrl.command_done~q ),
	.dgwb_wdp_ovride1(dgwb_wdp_ovride),
	.ac_muxctrl_broadcast_rcommand_req(\ac_mux:ctrl_broadcast_r.command_req~q ),
	.sig_addr_cmd0cke0(\dgwb|sig_addr_cmd[0].cke[0]~q ),
	.dgwb_ac_access_req1(\dgwb|dgwb_ac_access_req~q ),
	.sig_addr_cmd1cs_n0(\dgwb|sig_addr_cmd[1].cs_n[0]~q ),
	.sig_addr_cmd0addr12(\dgwb|sig_addr_cmd[0].addr[12]~q ),
	.sig_addr_cmd0rst_n(\dgwb|sig_addr_cmd[0].rst_n~q ),
	.dgwb_wdata_120(dgwb_wdata_120),
	.dgwb_wdata_56(dgwb_wdata_56),
	.dgwb_wdata_88(dgwb_wdata_88),
	.dgwb_wdata_24(dgwb_wdata_24),
	.dgwb_wdata_121(dgwb_wdata_121),
	.dgwb_wdata_57(dgwb_wdata_57),
	.dgwb_wdata_89(dgwb_wdata_89),
	.dgwb_wdata_25(dgwb_wdata_25),
	.dgwb_wdata_122(dgwb_wdata_122),
	.dgwb_wdata_58(dgwb_wdata_58),
	.dgwb_wdata_90(dgwb_wdata_90),
	.dgwb_wdata_26(dgwb_wdata_26),
	.dgwb_wdata_123(dgwb_wdata_123),
	.dgwb_wdata_59(dgwb_wdata_59),
	.dgwb_wdata_91(dgwb_wdata_91),
	.dgwb_wdata_27(dgwb_wdata_27),
	.dgwb_wdata_124(dgwb_wdata_124),
	.dgwb_wdata_60(dgwb_wdata_60),
	.dgwb_wdata_92(dgwb_wdata_92),
	.dgwb_wdata_28(dgwb_wdata_28),
	.dgwb_wdata_125(dgwb_wdata_125),
	.dgwb_wdata_61(dgwb_wdata_61),
	.dgwb_wdata_93(dgwb_wdata_93),
	.dgwb_wdata_29(dgwb_wdata_29),
	.dgwb_wdata_126(dgwb_wdata_126),
	.dgwb_wdata_62(dgwb_wdata_62),
	.dgwb_wdata_94(dgwb_wdata_94),
	.dgwb_wdata_30(dgwb_wdata_30),
	.dgwb_wdata_127(dgwb_wdata_127),
	.dgwb_wdata_63(dgwb_wdata_63),
	.dgwb_wdata_95(dgwb_wdata_95),
	.dgwb_wdata_31(dgwb_wdata_31),
	.dgwb_ctrlcommand_ack(\dgwb|dgwb_ctrl.command_ack~q ),
	.dgwb_wdp_ovride2(dgwb_wdp_ovride1));

ddr3_int_ddr3_int_phy_alt_mem_phy_admin admin(
	.clk(clk),
	.rst_n(rst_n),
	.ctl_init_fail(ctl_init_fail2),
	.ctl_init_success(ctl_init_success2),
	.curr_cmdcmd_prep_customer_mr_setup(\ctrl|curr_cmd.cmd_prep_customer_mr_setup~q ),
	.curr_cmdcmd_init_dram(\ctrl|curr_cmd.cmd_init_dram~q ),
	.curr_cmdcmd_prog_cal_mr(\ctrl|curr_cmd.cmd_prog_cal_mr~q ),
	.WideOr0(\ctrl|WideOr0~0_combout ),
	.admin_ctrlcommand_done(\admin|admin_ctrl.command_done~q ),
	.ac_access_gnt1(\admin|ac_access_gnt~q ),
	.seq_ac_sel1(seq_ac_sel),
	.ac_muxctrl_broadcast_rcommand_req(\ac_mux:ctrl_broadcast_r.command_req~q ),
	.dgrb_ac_access_req(\dgrb|dgrb_ac_access_req~q ),
	.dgwb_ac_access_req(\dgwb|dgwb_ac_access_req~q ),
	.addr_cmd0cs_n0(\admin|addr_cmd[0].cs_n[0]~q ),
	.addr_cmd1cs_n0(\admin|addr_cmd[1].cs_n[0]~q ),
	.addr_cmd0cke0(\admin|addr_cmd[0].cke[0]~q ),
	.addr_cmd0addr0(\admin|addr_cmd[0].addr[0]~q ),
	.addr_cmd1addr0(\admin|addr_cmd[1].addr[0]~q ),
	.addr_cmd0addr1(\admin|addr_cmd[0].addr[1]~q ),
	.addr_cmd1addr1(\admin|addr_cmd[1].addr[1]~q ),
	.addr_cmd0addr8(\admin|addr_cmd[0].addr[8]~q ),
	.addr_cmd1addr8(\admin|addr_cmd[1].addr[8]~q ),
	.addr_cmd0addr10(\admin|addr_cmd[0].addr[10]~q ),
	.addr_cmd1addr10(\admin|addr_cmd[1].addr[10]~q ),
	.addr_cmd0ba0(\admin|addr_cmd[0].ba[0]~q ),
	.addr_cmd1ba0(\admin|addr_cmd[1].ba[0]~q ),
	.addr_cmd0ba1(\admin|addr_cmd[0].ba[1]~q ),
	.addr_cmd1ba1(\admin|addr_cmd[1].ba[1]~q ),
	.addr_cmd0ras_n(\admin|addr_cmd[0].ras_n~q ),
	.addr_cmd1ras_n(\admin|addr_cmd[1].ras_n~q ),
	.addr_cmd0cas_n(\admin|addr_cmd[0].cas_n~q ),
	.addr_cmd1cas_n(\admin|addr_cmd[1].cas_n~q ),
	.addr_cmd0we_n(\admin|addr_cmd[0].we_n~q ),
	.addr_cmd1we_n(\admin|addr_cmd[1].we_n~q ),
	.addr_cmd0rst_n(\admin|addr_cmd[0].rst_n~q ),
	.dgb_ac_access_req(\dgb_ac_access_req~0_combout ),
	.admin_ctrlcommand_ack(\admin|admin_ctrl.command_ack~q ));

dffeas dgb_ac_access_gnt_r(
	.clk(clk),
	.d(\admin|ac_access_gnt~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dgb_ac_access_gnt_r~q ),
	.prn(vcc));
defparam dgb_ac_access_gnt_r.is_wysiwyg = "true";
defparam dgb_ac_access_gnt_r.power_up = "low";

arriaii_lcell_comb \seq_ac_ras_n[1]~0 (
	.dataa(!\admin|ac_access_gnt~q ),
	.datab(!\dgrb|dgrb_ac_access_req~q ),
	.datac(!\dgwb|dgwb_ac_access_req~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_ac_ras_n[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_ras_n[1]~0 .extended_lut = "off";
defparam \seq_ac_ras_n[1]~0 .lut_mask = 64'h1515151515151515;
defparam \seq_ac_ras_n[1]~0 .shared_arith = "off";

arriaii_lcell_comb \dgb_ac_access_req~0 (
	.dataa(!\dgrb|dgrb_ac_access_req~q ),
	.datab(!\dgwb|dgwb_ac_access_req~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dgb_ac_access_req~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dgb_ac_access_req~0 .extended_lut = "off";
defparam \dgb_ac_access_req~0 .lut_mask = 64'h6666666666666666;
defparam \dgb_ac_access_req~0 .shared_arith = "off";

dffeas dgrb_phs_shft_busy(
	.clk(clk),
	.d(\dgrb_phs_shft_busy~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dgrb_phs_shft_busy~q ),
	.prn(vcc));
defparam dgrb_phs_shft_busy.is_wysiwyg = "true";
defparam dgrb_phs_shft_busy.power_up = "low";

dffeas seq_pll_phs_shift_busy_ccd(
	.clk(clk),
	.d(\seq_pll_phs_shift_busy_r~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_pll_phs_shift_busy_ccd~q ),
	.prn(vcc));
defparam seq_pll_phs_shift_busy_ccd.is_wysiwyg = "true";
defparam seq_pll_phs_shift_busy_ccd.power_up = "low";

arriaii_lcell_comb \dgrb_phs_shft_busy~0 (
	.dataa(!\ctrl|state.s_was~q ),
	.datab(!\ctrl|state.s_prep_customer_mr_setup~q ),
	.datac(!\ctrl|Selector61~0_combout ),
	.datad(!\ctrl|WideOr35~0_combout ),
	.datae(!\seq_pll_phs_shift_busy_ccd~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dgrb_phs_shft_busy~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dgrb_phs_shft_busy~0 .extended_lut = "off";
defparam \dgrb_phs_shft_busy~0 .lut_mask = 64'h0000000800000008;
defparam \dgrb_phs_shft_busy~0 .shared_arith = "off";

dffeas seq_pll_phs_shift_busy_r(
	.clk(clk),
	.d(seq_pll_phs_shift_busy),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_pll_phs_shift_busy_r~q ),
	.prn(vcc));
defparam seq_pll_phs_shift_busy_r.is_wysiwyg = "true";
defparam seq_pll_phs_shift_busy_r.power_up = "low";

dffeas \seq_ac_cke[1] (
	.clk(clk),
	.d(\seq_ac_cke~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\ac_mux:mem_clk_disable[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_cke_1),
	.prn(vcc));
defparam \seq_ac_cke[1] .is_wysiwyg = "true";
defparam \seq_ac_cke[1] .power_up = "low";

dffeas \seq_ac_addr[0] (
	.clk(clk),
	.d(\seq_ac_addr~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\ac_mux:mem_clk_disable[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_addr_0),
	.prn(vcc));
defparam \seq_ac_addr[0] .is_wysiwyg = "true";
defparam \seq_ac_addr[0] .power_up = "low";

dffeas \seq_ac_addr[14] (
	.clk(clk),
	.d(\seq_ac_addr~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\ac_mux:mem_clk_disable[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_addr_14),
	.prn(vcc));
defparam \seq_ac_addr[14] .is_wysiwyg = "true";
defparam \seq_ac_addr[14] .power_up = "low";

dffeas \seq_ac_addr[1] (
	.clk(clk),
	.d(\seq_ac_addr~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\ac_mux:mem_clk_disable[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_addr_1),
	.prn(vcc));
defparam \seq_ac_addr[1] .is_wysiwyg = "true";
defparam \seq_ac_addr[1] .power_up = "low";

dffeas \seq_ac_addr[15] (
	.clk(clk),
	.d(\seq_ac_addr~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\ac_mux:mem_clk_disable[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_addr_15),
	.prn(vcc));
defparam \seq_ac_addr[15] .is_wysiwyg = "true";
defparam \seq_ac_addr[15] .power_up = "low";

dffeas \seq_ac_addr[16] (
	.clk(clk),
	.d(\seq_ac_addr~4_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\ac_mux:mem_clk_disable[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_addr_16),
	.prn(vcc));
defparam \seq_ac_addr[16] .is_wysiwyg = "true";
defparam \seq_ac_addr[16] .power_up = "low";

dffeas \seq_ac_addr[17] (
	.clk(clk),
	.d(\seq_ac_addr~5_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\ac_mux:mem_clk_disable[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_addr_17),
	.prn(vcc));
defparam \seq_ac_addr[17] .is_wysiwyg = "true";
defparam \seq_ac_addr[17] .power_up = "low";

dffeas \seq_ac_addr[18] (
	.clk(clk),
	.d(\seq_ac_addr~6_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\ac_mux:mem_clk_disable[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_addr_18),
	.prn(vcc));
defparam \seq_ac_addr[18] .is_wysiwyg = "true";
defparam \seq_ac_addr[18] .power_up = "low";

dffeas \seq_ac_addr[5] (
	.clk(clk),
	.d(\seq_ac_addr~7_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\ac_mux:mem_clk_disable[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_addr_5),
	.prn(vcc));
defparam \seq_ac_addr[5] .is_wysiwyg = "true";
defparam \seq_ac_addr[5] .power_up = "low";

dffeas \seq_ac_addr[19] (
	.clk(clk),
	.d(\seq_ac_addr~8_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\ac_mux:mem_clk_disable[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_addr_19),
	.prn(vcc));
defparam \seq_ac_addr[19] .is_wysiwyg = "true";
defparam \seq_ac_addr[19] .power_up = "low";

dffeas \seq_ac_addr[8] (
	.clk(clk),
	.d(\seq_ac_addr~9_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\ac_mux:mem_clk_disable[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_addr_8),
	.prn(vcc));
defparam \seq_ac_addr[8] .is_wysiwyg = "true";
defparam \seq_ac_addr[8] .power_up = "low";

dffeas \seq_ac_addr[22] (
	.clk(clk),
	.d(\seq_ac_addr~10_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\ac_mux:mem_clk_disable[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_addr_22),
	.prn(vcc));
defparam \seq_ac_addr[22] .is_wysiwyg = "true";
defparam \seq_ac_addr[22] .power_up = "low";

dffeas \seq_ac_addr[10] (
	.clk(clk),
	.d(\seq_ac_addr~11_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\ac_mux:mem_clk_disable[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_addr_10),
	.prn(vcc));
defparam \seq_ac_addr[10] .is_wysiwyg = "true";
defparam \seq_ac_addr[10] .power_up = "low";

dffeas \seq_ac_addr[24] (
	.clk(clk),
	.d(\seq_ac_addr~12_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\ac_mux:mem_clk_disable[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_addr_24),
	.prn(vcc));
defparam \seq_ac_addr[24] .is_wysiwyg = "true";
defparam \seq_ac_addr[24] .power_up = "low";

dffeas \seq_ac_addr[12] (
	.clk(clk),
	.d(\seq_ac_addr~13_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\ac_mux:mem_clk_disable[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_addr_12),
	.prn(vcc));
defparam \seq_ac_addr[12] .is_wysiwyg = "true";
defparam \seq_ac_addr[12] .power_up = "low";

dffeas \seq_ac_addr[26] (
	.clk(clk),
	.d(\seq_ac_addr~14_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\ac_mux:mem_clk_disable[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_addr_26),
	.prn(vcc));
defparam \seq_ac_addr[26] .is_wysiwyg = "true";
defparam \seq_ac_addr[26] .power_up = "low";

dffeas \seq_ac_ba[0] (
	.clk(clk),
	.d(\seq_ac_ba~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\ac_mux:mem_clk_disable[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_ba_0),
	.prn(vcc));
defparam \seq_ac_ba[0] .is_wysiwyg = "true";
defparam \seq_ac_ba[0] .power_up = "low";

dffeas \seq_ac_ba[3] (
	.clk(clk),
	.d(\seq_ac_ba~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\ac_mux:mem_clk_disable[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_ba_3),
	.prn(vcc));
defparam \seq_ac_ba[3] .is_wysiwyg = "true";
defparam \seq_ac_ba[3] .power_up = "low";

dffeas \seq_ac_ba[1] (
	.clk(clk),
	.d(\seq_ac_ba~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\ac_mux:mem_clk_disable[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_ba_1),
	.prn(vcc));
defparam \seq_ac_ba[1] .is_wysiwyg = "true";
defparam \seq_ac_ba[1] .power_up = "low";

dffeas \seq_ac_ba[4] (
	.clk(clk),
	.d(\seq_ac_ba~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\ac_mux:mem_clk_disable[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_ba_4),
	.prn(vcc));
defparam \seq_ac_ba[4] .is_wysiwyg = "true";
defparam \seq_ac_ba[4] .power_up = "low";

dffeas \seq_ac_rst_n[0] (
	.clk(clk),
	.d(\seq_ac_rst_n~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\ac_mux:mem_clk_disable[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_rst_n_0),
	.prn(vcc));
defparam \seq_ac_rst_n[0] .is_wysiwyg = "true";
defparam \seq_ac_rst_n[0] .power_up = "low";

dffeas ctl_init_fail(
	.clk(clk),
	.d(ctl_init_fail2),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ctl_init_fail1),
	.prn(vcc));
defparam ctl_init_fail.is_wysiwyg = "true";
defparam ctl_init_fail.power_up = "low";

dffeas ctl_init_success(
	.clk(clk),
	.d(ctl_init_success2),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ctl_init_success1),
	.prn(vcc));
defparam ctl_init_success.is_wysiwyg = "true";
defparam ctl_init_success.power_up = "low";

dffeas \seq_rdv_doing_rd[7] (
	.clk(clk),
	.d(\dgrb|sig_doing_rd[0]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_rdv_doing_rd_7),
	.prn(vcc));
defparam \seq_rdv_doing_rd[7] .is_wysiwyg = "true";
defparam \seq_rdv_doing_rd[7] .power_up = "low";

dffeas seq_rdp_reset_req_n(
	.clk(clk),
	.d(\seq_rdp_reset_req_n~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_rdp_reset_req_n1),
	.prn(vcc));
defparam seq_rdp_reset_req_n.is_wysiwyg = "true";
defparam seq_rdp_reset_req_n.power_up = "low";

dffeas seq_ac_add_1t_ac_lat_internal(
	.clk(clk),
	.d(\seq_ac_add_1t_ac_lat_internal~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_add_1t_ac_lat_internal1),
	.prn(vcc));
defparam seq_ac_add_1t_ac_lat_internal.is_wysiwyg = "true";
defparam seq_ac_add_1t_ac_lat_internal.power_up = "low";

dffeas seq_rdata_valid_lat_dec(
	.clk(clk),
	.d(\dgrb|seq_rdata_valid_lat_dec~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_rdata_valid_lat_dec1),
	.prn(vcc));
defparam seq_rdata_valid_lat_dec.is_wysiwyg = "true";
defparam seq_rdata_valid_lat_dec.power_up = "low";

dffeas \seq_rdv_doing_rd[4] (
	.clk(clk),
	.d(\dgrb|sig_doing_rd[4]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_rdv_doing_rd_4),
	.prn(vcc));
defparam \seq_rdv_doing_rd[4] .is_wysiwyg = "true";
defparam \seq_rdv_doing_rd[4] .power_up = "low";

dffeas seq_pll_inc_dec_n(
	.clk(clk),
	.d(\seq_pll_inc_dec_n~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_pll_inc_dec_n1),
	.prn(vcc));
defparam seq_pll_inc_dec_n.is_wysiwyg = "true";
defparam seq_pll_inc_dec_n.power_up = "low";

dffeas seq_pll_start_reconfig(
	.clk(clk),
	.d(\seq_pll_start_reconfig~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_pll_start_reconfig1),
	.prn(vcc));
defparam seq_pll_start_reconfig.is_wysiwyg = "true";
defparam seq_pll_start_reconfig.power_up = "low";

dffeas \seq_pll_select[2] (
	.clk(clk),
	.d(\seq_pll_select~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_pll_select_2),
	.prn(vcc));
defparam \seq_pll_select[2] .is_wysiwyg = "true";
defparam \seq_pll_select[2] .power_up = "low";

dffeas \seq_pll_select[1] (
	.clk(clk),
	.d(\seq_pll_select~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_pll_select_1),
	.prn(vcc));
defparam \seq_pll_select[1] .is_wysiwyg = "true";
defparam \seq_pll_select[1] .power_up = "low";

dffeas seq_mem_clk_disable(
	.clk(clk),
	.d(\ac_mux:mem_clk_disable[2]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_mem_clk_disable1),
	.prn(vcc));
defparam seq_mem_clk_disable.is_wysiwyg = "true";
defparam seq_mem_clk_disable.power_up = "low";

dffeas \seq_ac_cs_n[0] (
	.clk(clk),
	.d(\seq_ac_cs_n~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_cs_n_0),
	.prn(vcc));
defparam \seq_ac_cs_n[0] .is_wysiwyg = "true";
defparam \seq_ac_cs_n[0] .power_up = "low";

arriaii_lcell_comb \seq_wdp_ovride~0 (
	.dataa(!ctl_init_fail2),
	.datab(!ctl_init_success2),
	.datac(!dgwb_wdp_ovride),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(seq_wdp_ovride),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_wdp_ovride~0 .extended_lut = "off";
defparam \seq_wdp_ovride~0 .lut_mask = 64'h0808080808080808;
defparam \seq_wdp_ovride~0 .shared_arith = "off";

dffeas seq_poa_protection_override_1x(
	.clk(clk),
	.d(\WideNor0~combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_poa_protection_override_1x1),
	.prn(vcc));
defparam seq_poa_protection_override_1x.is_wysiwyg = "true";
defparam seq_poa_protection_override_1x.power_up = "low";

dffeas \seq_poa_lat_dec_1x[0] (
	.clk(clk),
	.d(\dgrb|seq_poa_lat_dec_1x[0]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_poa_lat_dec_1x_0),
	.prn(vcc));
defparam \seq_poa_lat_dec_1x[0] .is_wysiwyg = "true";
defparam \seq_poa_lat_dec_1x[0] .power_up = "low";

arriaii_lcell_comb \seq_ac_cas_n[0]~_wirecell (
	.dataa(!\seq_ac_cas_n[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(seq_ac_cas_n_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_cas_n[0]~_wirecell .extended_lut = "off";
defparam \seq_ac_cas_n[0]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \seq_ac_cas_n[0]~_wirecell .shared_arith = "off";

arriaii_lcell_comb \seq_ac_cas_n[1]~_wirecell (
	.dataa(!\seq_ac_cas_n[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(seq_ac_cas_n_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_cas_n[1]~_wirecell .extended_lut = "off";
defparam \seq_ac_cas_n[1]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \seq_ac_cas_n[1]~_wirecell .shared_arith = "off";

arriaii_lcell_comb \seq_ac_cs_n[1]~_wirecell (
	.dataa(!\seq_ac_cs_n[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(seq_ac_cs_n_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_cs_n[1]~_wirecell .extended_lut = "off";
defparam \seq_ac_cs_n[1]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \seq_ac_cs_n[1]~_wirecell .shared_arith = "off";

arriaii_lcell_comb \seq_ac_ras_n[0]~_wirecell (
	.dataa(!\seq_ac_ras_n[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(seq_ac_ras_n_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_ras_n[0]~_wirecell .extended_lut = "off";
defparam \seq_ac_ras_n[0]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \seq_ac_ras_n[0]~_wirecell .shared_arith = "off";

arriaii_lcell_comb \seq_ac_ras_n[1]~_wirecell (
	.dataa(!\seq_ac_ras_n[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(seq_ac_ras_n_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_ras_n[1]~_wirecell .extended_lut = "off";
defparam \seq_ac_ras_n[1]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \seq_ac_ras_n[1]~_wirecell .shared_arith = "off";

arriaii_lcell_comb \seq_ac_we_n[0]~_wirecell (
	.dataa(!\seq_ac_we_n[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(seq_ac_we_n_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_we_n[0]~_wirecell .extended_lut = "off";
defparam \seq_ac_we_n[0]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \seq_ac_we_n[0]~_wirecell .shared_arith = "off";

arriaii_lcell_comb \seq_ac_we_n[1]~_wirecell (
	.dataa(!\seq_ac_we_n[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(seq_ac_we_n_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_we_n[1]~_wirecell .extended_lut = "off";
defparam \seq_ac_we_n[1]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \seq_ac_we_n[1]~_wirecell .shared_arith = "off";

arriaii_lcell_comb \seq_ac_cke~0 (
	.dataa(!\admin|ac_access_gnt~q ),
	.datab(!\dgwb|sig_addr_cmd[0].cke[0]~q ),
	.datac(!\dgrb|dgrb_ac_access_req~q ),
	.datad(!\dgwb|dgwb_ac_access_req~q ),
	.datae(!\admin|addr_cmd[0].cke[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_ac_cke~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_cke~0 .extended_lut = "off";
defparam \seq_ac_cke~0 .lut_mask = 64'h0111FBBB0111FBBB;
defparam \seq_ac_cke~0 .shared_arith = "off";

dffeas \ac_mux:ctrl_broadcast_r.command_req (
	.clk(clk),
	.d(\ctrl|Selector61~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_mux:ctrl_broadcast_r.command_req~q ),
	.prn(vcc));
defparam \ac_mux:ctrl_broadcast_r.command_req .is_wysiwyg = "true";
defparam \ac_mux:ctrl_broadcast_r.command_req .power_up = "low";

arriaii_lcell_comb \ac_mux:mem_clk_disable[0]~0 (
	.dataa(!\ctrl|curr_cmd.cmd_init_dram~q ),
	.datab(!\ac_mux:ctrl_broadcast_r.command_req~q ),
	.datac(!\ac_mux:mem_clk_disable[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_mux:mem_clk_disable[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_mux:mem_clk_disable[0]~0 .extended_lut = "off";
defparam \ac_mux:mem_clk_disable[0]~0 .lut_mask = 64'h1F1F1F1F1F1F1F1F;
defparam \ac_mux:mem_clk_disable[0]~0 .shared_arith = "off";

dffeas \ac_mux:mem_clk_disable[0] (
	.clk(clk),
	.d(\ac_mux:mem_clk_disable[0]~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_mux:mem_clk_disable[0]~q ),
	.prn(vcc));
defparam \ac_mux:mem_clk_disable[0] .is_wysiwyg = "true";
defparam \ac_mux:mem_clk_disable[0] .power_up = "low";

arriaii_lcell_comb \seq_ac_addr~0 (
	.dataa(!\admin|ac_access_gnt~q ),
	.datab(!\dgrb|dgrb_ac_access_req~q ),
	.datac(!\dgwb|dgwb_ac_access_req~q ),
	.datad(!\admin|addr_cmd[0].addr[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_ac_addr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_addr~0 .extended_lut = "off";
defparam \seq_ac_addr~0 .lut_mask = 64'h00EA00EA00EA00EA;
defparam \seq_ac_addr~0 .shared_arith = "off";

arriaii_lcell_comb \seq_ac_addr~1 (
	.dataa(!\admin|ac_access_gnt~q ),
	.datab(!\dgrb|dgrb_ac_access_req~q ),
	.datac(!\dgwb|dgwb_ac_access_req~q ),
	.datad(!\admin|addr_cmd[1].addr[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_ac_addr~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_addr~1 .extended_lut = "off";
defparam \seq_ac_addr~1 .lut_mask = 64'h00EA00EA00EA00EA;
defparam \seq_ac_addr~1 .shared_arith = "off";

arriaii_lcell_comb \seq_ac_addr~2 (
	.dataa(!\admin|ac_access_gnt~q ),
	.datab(!\dgrb|dgrb_ac_access_req~q ),
	.datac(!\dgwb|dgwb_ac_access_req~q ),
	.datad(!\admin|addr_cmd[0].addr[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_ac_addr~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_addr~2 .extended_lut = "off";
defparam \seq_ac_addr~2 .lut_mask = 64'h00EA00EA00EA00EA;
defparam \seq_ac_addr~2 .shared_arith = "off";

arriaii_lcell_comb \seq_ac_addr~3 (
	.dataa(!\admin|ac_access_gnt~q ),
	.datab(!\dgrb|dgrb_ac_access_req~q ),
	.datac(!\dgwb|dgwb_ac_access_req~q ),
	.datad(!\admin|addr_cmd[1].addr[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_ac_addr~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_addr~3 .extended_lut = "off";
defparam \seq_ac_addr~3 .lut_mask = 64'h00EA00EA00EA00EA;
defparam \seq_ac_addr~3 .shared_arith = "off";

arriaii_lcell_comb \seq_ac_addr~4 (
	.dataa(!\admin|ac_access_gnt~q ),
	.datab(!\dgwb|dgwb_ac_access_req~q ),
	.datac(!\dgwb|sig_addr_cmd[0].addr[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_ac_addr~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_addr~4 .extended_lut = "off";
defparam \seq_ac_addr~4 .lut_mask = 64'h0101010101010101;
defparam \seq_ac_addr~4 .shared_arith = "off";

arriaii_lcell_comb \seq_ac_addr~5 (
	.dataa(!\admin|ac_access_gnt~q ),
	.datab(!\dgrb|dgrb_ac_access_req~q ),
	.datac(!\dgwb|dgwb_ac_access_req~q ),
	.datad(!\dgwb|sig_addr_cmd[0].addr[3]~q ),
	.datae(!\dgrb|sig_addr_cmd[0].addr[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_ac_addr~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_addr~5 .extended_lut = "off";
defparam \seq_ac_addr~5 .lut_mask = 64'h0005101500051015;
defparam \seq_ac_addr~5 .shared_arith = "off";

arriaii_lcell_comb \seq_ac_addr~6 (
	.dataa(!\admin|ac_access_gnt~q ),
	.datab(!\dgrb|dgrb_ac_access_req~q ),
	.datac(!\dgwb|dgwb_ac_access_req~q ),
	.datad(!\dgwb|sig_addr_cmd[0].addr[4]~q ),
	.datae(!\dgrb|sig_addr_cmd[0].addr[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_ac_addr~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_addr~6 .extended_lut = "off";
defparam \seq_ac_addr~6 .lut_mask = 64'h0005101500051015;
defparam \seq_ac_addr~6 .shared_arith = "off";

arriaii_lcell_comb \process_4~1 (
	.dataa(!\admin|ac_access_gnt~q ),
	.datab(!\dgwb|dgwb_ac_access_req~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\process_4~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \process_4~1 .extended_lut = "off";
defparam \process_4~1 .lut_mask = 64'h1111111111111111;
defparam \process_4~1 .shared_arith = "off";

arriaii_lcell_comb \process_4~2 (
	.dataa(!\admin|ac_access_gnt~q ),
	.datab(!\dgrb|dgrb_ac_access_req~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\process_4~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \process_4~2 .extended_lut = "off";
defparam \process_4~2 .lut_mask = 64'h1111111111111111;
defparam \process_4~2 .shared_arith = "off";

arriaii_lcell_comb \seq_ac_addr~7 (
	.dataa(!\process_4~1_combout ),
	.datab(!\process_4~2_combout ),
	.datac(!\admin|addr_cmd[0].addr[0]~q ),
	.datad(!\dgwb|sig_addr_cmd[0].addr[5]~q ),
	.datae(!\dgrb|sig_addr_cmd[0].addr[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_ac_addr~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_addr~7 .extended_lut = "off";
defparam \seq_ac_addr~7 .lut_mask = 64'h085D2A7F085D2A7F;
defparam \seq_ac_addr~7 .shared_arith = "off";

arriaii_lcell_comb \seq_ac_addr~8 (
	.dataa(!\process_4~1_combout ),
	.datab(!\process_4~2_combout ),
	.datac(!\admin|addr_cmd[1].addr[0]~q ),
	.datad(!\dgwb|sig_addr_cmd[0].addr[5]~q ),
	.datae(!\dgrb|sig_addr_cmd[0].addr[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_ac_addr~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_addr~8 .extended_lut = "off";
defparam \seq_ac_addr~8 .lut_mask = 64'h085D2A7F085D2A7F;
defparam \seq_ac_addr~8 .shared_arith = "off";

arriaii_lcell_comb \seq_ac_addr~9 (
	.dataa(!\admin|ac_access_gnt~q ),
	.datab(!\dgrb|dgrb_ac_access_req~q ),
	.datac(!\dgwb|dgwb_ac_access_req~q ),
	.datad(!\admin|addr_cmd[0].addr[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_ac_addr~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_addr~9 .extended_lut = "off";
defparam \seq_ac_addr~9 .lut_mask = 64'h00EA00EA00EA00EA;
defparam \seq_ac_addr~9 .shared_arith = "off";

arriaii_lcell_comb \seq_ac_addr~10 (
	.dataa(!\admin|ac_access_gnt~q ),
	.datab(!\dgrb|dgrb_ac_access_req~q ),
	.datac(!\dgwb|dgwb_ac_access_req~q ),
	.datad(!\admin|addr_cmd[1].addr[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_ac_addr~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_addr~10 .extended_lut = "off";
defparam \seq_ac_addr~10 .lut_mask = 64'h00EA00EA00EA00EA;
defparam \seq_ac_addr~10 .shared_arith = "off";

arriaii_lcell_comb \seq_ac_addr~11 (
	.dataa(!\admin|ac_access_gnt~q ),
	.datab(!\dgrb|dgrb_ac_access_req~q ),
	.datac(!\dgwb|dgwb_ac_access_req~q ),
	.datad(!\admin|addr_cmd[0].addr[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_ac_addr~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_addr~11 .extended_lut = "off";
defparam \seq_ac_addr~11 .lut_mask = 64'h00EA00EA00EA00EA;
defparam \seq_ac_addr~11 .shared_arith = "off";

arriaii_lcell_comb \seq_ac_addr~12 (
	.dataa(!\admin|ac_access_gnt~q ),
	.datab(!\dgrb|dgrb_ac_access_req~q ),
	.datac(!\dgwb|dgwb_ac_access_req~q ),
	.datad(!\admin|addr_cmd[1].addr[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_ac_addr~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_addr~12 .extended_lut = "off";
defparam \seq_ac_addr~12 .lut_mask = 64'h00EA00EA00EA00EA;
defparam \seq_ac_addr~12 .shared_arith = "off";

arriaii_lcell_comb \seq_ac_addr~13 (
	.dataa(!\process_4~1_combout ),
	.datab(!\process_4~2_combout ),
	.datac(!\admin|addr_cmd[0].addr[0]~q ),
	.datad(!\dgwb|sig_addr_cmd[0].addr[12]~q ),
	.datae(!\dgrb|sig_addr_cmd[0].addr[12]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_ac_addr~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_addr~13 .extended_lut = "off";
defparam \seq_ac_addr~13 .lut_mask = 64'h085D2A7F085D2A7F;
defparam \seq_ac_addr~13 .shared_arith = "off";

arriaii_lcell_comb \seq_ac_addr~14 (
	.dataa(!\process_4~1_combout ),
	.datab(!\process_4~2_combout ),
	.datac(!\admin|addr_cmd[1].addr[0]~q ),
	.datad(!\dgwb|sig_addr_cmd[0].addr[12]~q ),
	.datae(!\dgrb|sig_addr_cmd[0].addr[12]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_ac_addr~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_addr~14 .extended_lut = "off";
defparam \seq_ac_addr~14 .lut_mask = 64'h085D2A7F085D2A7F;
defparam \seq_ac_addr~14 .shared_arith = "off";

arriaii_lcell_comb \seq_ac_ba~0 (
	.dataa(!\admin|ac_access_gnt~q ),
	.datab(!\dgrb|dgrb_ac_access_req~q ),
	.datac(!\dgwb|dgwb_ac_access_req~q ),
	.datad(!\admin|addr_cmd[0].ba[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_ac_ba~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_ba~0 .extended_lut = "off";
defparam \seq_ac_ba~0 .lut_mask = 64'h00EA00EA00EA00EA;
defparam \seq_ac_ba~0 .shared_arith = "off";

arriaii_lcell_comb \seq_ac_ba~1 (
	.dataa(!\admin|ac_access_gnt~q ),
	.datab(!\dgrb|dgrb_ac_access_req~q ),
	.datac(!\dgwb|dgwb_ac_access_req~q ),
	.datad(!\admin|addr_cmd[1].ba[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_ac_ba~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_ba~1 .extended_lut = "off";
defparam \seq_ac_ba~1 .lut_mask = 64'h00EA00EA00EA00EA;
defparam \seq_ac_ba~1 .shared_arith = "off";

arriaii_lcell_comb \seq_ac_ba~2 (
	.dataa(!\admin|ac_access_gnt~q ),
	.datab(!\dgrb|dgrb_ac_access_req~q ),
	.datac(!\dgwb|dgwb_ac_access_req~q ),
	.datad(!\admin|addr_cmd[0].ba[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_ac_ba~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_ba~2 .extended_lut = "off";
defparam \seq_ac_ba~2 .lut_mask = 64'h00EA00EA00EA00EA;
defparam \seq_ac_ba~2 .shared_arith = "off";

arriaii_lcell_comb \seq_ac_ba~3 (
	.dataa(!\admin|ac_access_gnt~q ),
	.datab(!\dgrb|dgrb_ac_access_req~q ),
	.datac(!\dgwb|dgwb_ac_access_req~q ),
	.datad(!\admin|addr_cmd[1].ba[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_ac_ba~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_ba~3 .extended_lut = "off";
defparam \seq_ac_ba~3 .lut_mask = 64'h00EA00EA00EA00EA;
defparam \seq_ac_ba~3 .shared_arith = "off";

arriaii_lcell_comb \seq_ac_rst_n~0 (
	.dataa(!\admin|ac_access_gnt~q ),
	.datab(!\dgrb|dgrb_ac_access_req~q ),
	.datac(!\dgwb|dgwb_ac_access_req~q ),
	.datad(!\dgwb|sig_addr_cmd[0].rst_n~q ),
	.datae(!\admin|addr_cmd[0].rst_n~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_ac_rst_n~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_rst_n~0 .extended_lut = "off";
defparam \seq_ac_rst_n~0 .lut_mask = 64'h0015EAFF0015EAFF;
defparam \seq_ac_rst_n~0 .shared_arith = "off";

arriaii_lcell_comb \seq_rdp_reset_req_n~0 (
	.dataa(!seq_rdp_reset_req_n1),
	.datab(!\ctrl|state.s_rrp_sweep~q ),
	.datac(!\ctrl|master_ctrl_op_rec~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_rdp_reset_req_n~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_rdp_reset_req_n~0 .extended_lut = "off";
defparam \seq_rdp_reset_req_n~0 .lut_mask = 64'h7575757575757575;
defparam \seq_rdp_reset_req_n~0 .shared_arith = "off";

arriaii_lcell_comb \seq_ac_add_1t_ac_lat_internal~0 (
	.dataa(!\ctrl|ac_nt[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_ac_add_1t_ac_lat_internal~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_add_1t_ac_lat_internal~0 .extended_lut = "off";
defparam \seq_ac_add_1t_ac_lat_internal~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \seq_ac_add_1t_ac_lat_internal~0 .shared_arith = "off";

arriaii_lcell_comb \seq_pll_inc_dec_n~0 (
	.dataa(!\ctrl|state.s_was~q ),
	.datab(!\ctrl|state.s_prep_customer_mr_setup~q ),
	.datac(!\dgrb|seq_pll_inc_dec_n~q ),
	.datad(!\ctrl|Selector61~0_combout ),
	.datae(!\ctrl|WideOr35~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_pll_inc_dec_n~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_pll_inc_dec_n~0 .extended_lut = "off";
defparam \seq_pll_inc_dec_n~0 .lut_mask = 64'h0000000800000008;
defparam \seq_pll_inc_dec_n~0 .shared_arith = "off";

arriaii_lcell_comb \seq_pll_start_reconfig~0 (
	.dataa(!\ctrl|state.s_was~q ),
	.datab(!\ctrl|state.s_prep_customer_mr_setup~q ),
	.datac(!\ctrl|Selector61~0_combout ),
	.datad(!\ctrl|WideOr35~0_combout ),
	.datae(!\dgrb|seq_pll_start_reconfig~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_pll_start_reconfig~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_pll_start_reconfig~0 .extended_lut = "off";
defparam \seq_pll_start_reconfig~0 .lut_mask = 64'h0000000800000008;
defparam \seq_pll_start_reconfig~0 .shared_arith = "off";

arriaii_lcell_comb \seq_pll_select~0 (
	.dataa(!\ctrl|state.s_was~q ),
	.datab(!\ctrl|state.s_prep_customer_mr_setup~q ),
	.datac(!\ctrl|Selector61~0_combout ),
	.datad(!\ctrl|WideOr35~0_combout ),
	.datae(!\dgrb|seq_pll_select[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_pll_select~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_pll_select~0 .extended_lut = "off";
defparam \seq_pll_select~0 .lut_mask = 64'h0000000800000008;
defparam \seq_pll_select~0 .shared_arith = "off";

arriaii_lcell_comb \seq_pll_select~1 (
	.dataa(!\ctrl|state.s_was~q ),
	.datab(!\ctrl|state.s_prep_customer_mr_setup~q ),
	.datac(!\ctrl|Selector61~0_combout ),
	.datad(!\ctrl|WideOr35~0_combout ),
	.datae(!\dgrb|seq_pll_select[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_pll_select~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_pll_select~1 .extended_lut = "off";
defparam \seq_pll_select~1 .lut_mask = 64'h0000000800000008;
defparam \seq_pll_select~1 .shared_arith = "off";

dffeas \ac_mux:mem_clk_disable[1] (
	.clk(clk),
	.d(\ac_mux:mem_clk_disable[0]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_mux:mem_clk_disable[1]~q ),
	.prn(vcc));
defparam \ac_mux:mem_clk_disable[1] .is_wysiwyg = "true";
defparam \ac_mux:mem_clk_disable[1] .power_up = "low";

dffeas \ac_mux:mem_clk_disable[2] (
	.clk(clk),
	.d(\ac_mux:mem_clk_disable[1]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_mux:mem_clk_disable[2]~q ),
	.prn(vcc));
defparam \ac_mux:mem_clk_disable[2] .is_wysiwyg = "true";
defparam \ac_mux:mem_clk_disable[2] .power_up = "low";

arriaii_lcell_comb \seq_ac_cs_n~0 (
	.dataa(!\admin|ac_access_gnt~q ),
	.datab(!\dgrb|dgrb_ac_access_req~q ),
	.datac(!\dgwb|dgwb_ac_access_req~q ),
	.datad(!\ac_mux:mem_clk_disable[0]~q ),
	.datae(!\admin|addr_cmd[0].cs_n[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_ac_cs_n~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_cs_n~0 .extended_lut = "off";
defparam \seq_ac_cs_n~0 .lut_mask = 64'h000000EA000000EA;
defparam \seq_ac_cs_n~0 .shared_arith = "off";

arriaii_lcell_comb WideNor0(
	.dataa(!\ctrl|state.s_rrp_sweep~q ),
	.datab(!\ctrl|state.s_rdv~q ),
	.datac(!\ctrl|state.s_rrp_seek~q ),
	.datad(!\ctrl|state.s_adv_wr_lat~q ),
	.datae(!\ctrl|state.s_adv_rd_lat~q ),
	.dataf(!\ctrl|master_ctrl_op_rec~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideNor0.extended_lut = "off";
defparam WideNor0.lut_mask = 64'h7FFFFFFF00000000;
defparam WideNor0.shared_arith = "off";

arriaii_lcell_comb \seq_ac_ras_n[1]~1 (
	.dataa(!\admin|ac_access_gnt~q ),
	.datab(!\dgrb|dgrb_ac_access_req~q ),
	.datac(!\dgwb|dgwb_ac_access_req~q ),
	.datad(!\ac_mux:mem_clk_disable[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_ac_ras_n[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_ras_n[1]~1 .extended_lut = "off";
defparam \seq_ac_ras_n[1]~1 .lut_mask = 64'h00EF00EF00EF00EF;
defparam \seq_ac_ras_n[1]~1 .shared_arith = "off";

arriaii_lcell_comb \seq_ac_cas_n~0 (
	.dataa(!\seq_ac_ras_n[1]~0_combout ),
	.datab(!\ac_mux:mem_clk_disable[0]~q ),
	.datac(!\seq_ac_ras_n[1]~1_combout ),
	.datad(!\dgrb|sig_addr_cmd[0].addr[12]~q ),
	.datae(!\admin|addr_cmd[0].cas_n~q ),
	.dataf(!\dgwb|sig_addr_cmd[0].cas_n~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_ac_cas_n~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_cas_n~0 .extended_lut = "off";
defparam \seq_ac_cas_n~0 .lut_mask = 64'h2030223221312333;
defparam \seq_ac_cas_n~0 .shared_arith = "off";

dffeas \seq_ac_cas_n[0] (
	.clk(clk),
	.d(\seq_ac_cas_n~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_ac_cas_n[0]~q ),
	.prn(vcc));
defparam \seq_ac_cas_n[0] .is_wysiwyg = "true";
defparam \seq_ac_cas_n[0] .power_up = "low";

arriaii_lcell_comb \seq_ac_cas_n~1 (
	.dataa(!\seq_ac_ras_n[1]~0_combout ),
	.datab(!\ac_mux:mem_clk_disable[0]~q ),
	.datac(!\seq_ac_ras_n[1]~1_combout ),
	.datad(!\dgrb|sig_addr_cmd[0].addr[12]~q ),
	.datae(!\dgwb|sig_addr_cmd[0].cas_n~q ),
	.dataf(!\admin|addr_cmd[1].cas_n~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_ac_cas_n~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_cas_n~1 .extended_lut = "off";
defparam \seq_ac_cas_n~1 .lut_mask = 64'h2030213122322333;
defparam \seq_ac_cas_n~1 .shared_arith = "off";

dffeas \seq_ac_cas_n[1] (
	.clk(clk),
	.d(\seq_ac_cas_n~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_ac_cas_n[1]~q ),
	.prn(vcc));
defparam \seq_ac_cas_n[1] .is_wysiwyg = "true";
defparam \seq_ac_cas_n[1] .power_up = "low";

arriaii_lcell_comb \seq_ac_cs_n~1 (
	.dataa(!\seq_ac_ras_n[1]~0_combout ),
	.datab(!\ac_mux:mem_clk_disable[0]~q ),
	.datac(!\dgwb|sig_addr_cmd[1].cs_n[0]~q ),
	.datad(!\seq_ac_ras_n[1]~1_combout ),
	.datae(!\dgrb|sig_addr_cmd[1].cs_n[0]~q ),
	.dataf(!\admin|addr_cmd[1].cs_n[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_ac_cs_n~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_cs_n~1 .extended_lut = "off";
defparam \seq_ac_cs_n~1 .lut_mask = 64'h2201330122233323;
defparam \seq_ac_cs_n~1 .shared_arith = "off";

dffeas \seq_ac_cs_n[1] (
	.clk(clk),
	.d(\seq_ac_cs_n~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_ac_cs_n[1]~q ),
	.prn(vcc));
defparam \seq_ac_cs_n[1] .is_wysiwyg = "true";
defparam \seq_ac_cs_n[1] .power_up = "low";

arriaii_lcell_comb \seq_ac_ras_n~2 (
	.dataa(!\admin|ac_access_gnt~q ),
	.datab(!\dgrb|dgrb_ac_access_req~q ),
	.datac(!\dgwb|dgwb_ac_access_req~q ),
	.datad(!\ac_mux:mem_clk_disable[0]~q ),
	.datae(!\admin|addr_cmd[0].ras_n~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_ac_ras_n~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_ras_n~2 .extended_lut = "off";
defparam \seq_ac_ras_n~2 .lut_mask = 64'h000000EA000000EA;
defparam \seq_ac_ras_n~2 .shared_arith = "off";

dffeas \seq_ac_ras_n[0] (
	.clk(clk),
	.d(\seq_ac_ras_n~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_ac_ras_n[0]~q ),
	.prn(vcc));
defparam \seq_ac_ras_n[0] .is_wysiwyg = "true";
defparam \seq_ac_ras_n[0] .power_up = "low";

arriaii_lcell_comb \seq_ac_ras_n~3 (
	.dataa(!\admin|ac_access_gnt~q ),
	.datab(!\dgrb|dgrb_ac_access_req~q ),
	.datac(!\dgwb|dgwb_ac_access_req~q ),
	.datad(!\ac_mux:mem_clk_disable[0]~q ),
	.datae(!\admin|addr_cmd[1].ras_n~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_ac_ras_n~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_ras_n~3 .extended_lut = "off";
defparam \seq_ac_ras_n~3 .lut_mask = 64'h000000EA000000EA;
defparam \seq_ac_ras_n~3 .shared_arith = "off";

dffeas \seq_ac_ras_n[1] (
	.clk(clk),
	.d(\seq_ac_ras_n~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_ac_ras_n[1]~q ),
	.prn(vcc));
defparam \seq_ac_ras_n[1] .is_wysiwyg = "true";
defparam \seq_ac_ras_n[1] .power_up = "low";

arriaii_lcell_comb \seq_ac_we_n~0 (
	.dataa(!\seq_ac_ras_n[1]~0_combout ),
	.datab(!\ac_mux:mem_clk_disable[0]~q ),
	.datac(!\seq_ac_ras_n[1]~1_combout ),
	.datad(!\dgwb|sig_addr_cmd[0].cas_n~q ),
	.datae(!\admin|addr_cmd[0].we_n~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_ac_we_n~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_we_n~0 .extended_lut = "off";
defparam \seq_ac_we_n~0 .lut_mask = 64'h00010E0F00010E0F;
defparam \seq_ac_we_n~0 .shared_arith = "off";

dffeas \seq_ac_we_n[0] (
	.clk(clk),
	.d(\seq_ac_we_n~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_ac_we_n[0]~q ),
	.prn(vcc));
defparam \seq_ac_we_n[0] .is_wysiwyg = "true";
defparam \seq_ac_we_n[0] .power_up = "low";

arriaii_lcell_comb \seq_ac_we_n~1 (
	.dataa(!\seq_ac_ras_n[1]~0_combout ),
	.datab(!\ac_mux:mem_clk_disable[0]~q ),
	.datac(!\seq_ac_ras_n[1]~1_combout ),
	.datad(!\dgwb|sig_addr_cmd[0].cas_n~q ),
	.datae(!\admin|addr_cmd[1].we_n~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_ac_we_n~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_ac_we_n~1 .extended_lut = "off";
defparam \seq_ac_we_n~1 .lut_mask = 64'h00010E0F00010E0F;
defparam \seq_ac_we_n~1 .shared_arith = "off";

dffeas \seq_ac_we_n[1] (
	.clk(clk),
	.d(\seq_ac_we_n~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_ac_we_n[1]~q ),
	.prn(vcc));
defparam \seq_ac_we_n[1] .is_wysiwyg = "true";
defparam \seq_ac_we_n[1] .power_up = "low";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_admin (
	clk,
	rst_n,
	ctl_init_fail,
	ctl_init_success,
	curr_cmdcmd_prep_customer_mr_setup,
	curr_cmdcmd_init_dram,
	curr_cmdcmd_prog_cal_mr,
	WideOr0,
	admin_ctrlcommand_done,
	ac_access_gnt1,
	seq_ac_sel1,
	ac_muxctrl_broadcast_rcommand_req,
	dgrb_ac_access_req,
	dgwb_ac_access_req,
	addr_cmd0cs_n0,
	addr_cmd1cs_n0,
	addr_cmd0cke0,
	addr_cmd0addr0,
	addr_cmd1addr0,
	addr_cmd0addr1,
	addr_cmd1addr1,
	addr_cmd0addr8,
	addr_cmd1addr8,
	addr_cmd0addr10,
	addr_cmd1addr10,
	addr_cmd0ba0,
	addr_cmd1ba0,
	addr_cmd0ba1,
	addr_cmd1ba1,
	addr_cmd0ras_n,
	addr_cmd1ras_n,
	addr_cmd0cas_n,
	addr_cmd1cas_n,
	addr_cmd0we_n,
	addr_cmd1we_n,
	addr_cmd0rst_n,
	dgb_ac_access_req,
	admin_ctrlcommand_ack)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	rst_n;
input 	ctl_init_fail;
input 	ctl_init_success;
input 	curr_cmdcmd_prep_customer_mr_setup;
input 	curr_cmdcmd_init_dram;
input 	curr_cmdcmd_prog_cal_mr;
input 	WideOr0;
output 	admin_ctrlcommand_done;
output 	ac_access_gnt1;
output 	seq_ac_sel1;
input 	ac_muxctrl_broadcast_rcommand_req;
input 	dgrb_ac_access_req;
input 	dgwb_ac_access_req;
output 	addr_cmd0cs_n0;
output 	addr_cmd1cs_n0;
output 	addr_cmd0cke0;
output 	addr_cmd0addr0;
output 	addr_cmd1addr0;
output 	addr_cmd0addr1;
output 	addr_cmd1addr1;
output 	addr_cmd0addr8;
output 	addr_cmd1addr8;
output 	addr_cmd0addr10;
output 	addr_cmd1addr10;
output 	addr_cmd0ba0;
output 	addr_cmd1ba0;
output 	addr_cmd0ba1;
output 	addr_cmd1ba1;
output 	addr_cmd0ras_n;
output 	addr_cmd1ras_n;
output 	addr_cmd0cas_n;
output 	addr_cmd1cas_n;
output 	addr_cmd0we_n;
output 	addr_cmd1we_n;
output 	addr_cmd0rst_n;
input 	dgb_ac_access_req;
output 	admin_ctrlcommand_ack;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~5_sumout ;
wire \Add0~9_sumout ;
wire \Add0~13_sumout ;
wire \Add0~17_sumout ;
wire \refresh_count~10_combout ;
wire \refresh_count[3]~q ;
wire \refresh_count~11_combout ;
wire \refresh_count[2]~q ;
wire \refresh_count~9_combout ;
wire \refresh_count[1]~q ;
wire \refresh_count~8_combout ;
wire \refresh_count[0]~q ;
wire \Add0~2 ;
wire \Add0~6 ;
wire \Add0~10 ;
wire \Add0~14 ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \refresh_count~3_combout ;
wire \refresh_count[5]~q ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \refresh_count~4_combout ;
wire \refresh_count[6]~q ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \refresh_count~5_combout ;
wire \refresh_count[7]~q ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \refresh_count~7_combout ;
wire \refresh_count[8]~q ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \refresh_count~6_combout ;
wire \refresh_count[9]~q ;
wire \Equal0~0_combout ;
wire \Equal0~1_combout ;
wire \state~38_combout ;
wire \state.s_reset~0_combout ;
wire \state.s_reset~q ;
wire \WideOr34~0_combout ;
wire \Selector431~0_combout ;
wire \ac_state.s_9~q ;
wire \Selector432~0_combout ;
wire \ac_state.s_10~q ;
wire \Selector433~1_combout ;
wire \ac_state.s_11~q ;
wire \Selector434~0_combout ;
wire \ac_state.s_12~q ;
wire \Selector3~0_combout ;
wire \state~43_combout ;
wire \state~50_combout ;
wire \state~36_combout ;
wire \state~40_combout ;
wire \state~41_combout ;
wire \state.s_program_cal_mrs~q ;
wire \ac_state~19_combout ;
wire \stage_counter[17]~1_combout ;
wire \process_12~0_combout ;
wire \ac_state~20_combout ;
wire \ac_state~24_combout ;
wire \ac_state.s_3~q ;
wire \ac_state~23_combout ;
wire \ac_state.s_4~q ;
wire \ac_state~22_combout ;
wire \ac_state.s_5~q ;
wire \WideOr32~combout ;
wire \Selector421~1_combout ;
wire \per_cs_init_seen[0]~q ;
wire \mem_init_complete~q ;
wire \state~51_combout ;
wire \state~52_combout ;
wire \state.s_topup_refresh~q ;
wire \state~48_combout ;
wire \state.s_topup_refresh_done~q ;
wire \state~42_combout ;
wire \Selector15~0_combout ;
wire \command_started~q ;
wire \admin_req_extended~0_combout ;
wire \admin_req_extended~q ;
wire \state~44_combout ;
wire \state.s_prog_user_mrs~q ;
wire \ac_state~21_combout ;
wire \ac_state.s_6~q ;
wire \Selector429~0_combout ;
wire \ac_state.s_7~q ;
wire \Selector430~0_combout ;
wire \ac_state.s_8~q ;
wire \WideOr16~combout ;
wire \ac_state.s_1~0_combout ;
wire \ac_state.s_1~q ;
wire \cal_complete~combout ;
wire \state~56_combout ;
wire \state~61_combout ;
wire \state.s_zq_cal_short~q ;
wire \state~45_combout ;
wire \state.s_access_act~q ;
wire \state~34_combout ;
wire \state.s_access~q ;
wire \state~46_combout ;
wire \state~47_combout ;
wire \state.s_dummy_wait~q ;
wire \state~53_combout ;
wire \state~54_combout ;
wire \state.s_refresh~q ;
wire \state~55_combout ;
wire \state.s_access_precharge~q ;
wire \Selector422~1_combout ;
wire \Selector424~0_combout ;
wire \ac_state.s_2~q ;
wire \WideNor1~0_combout ;
wire \WideNor1~1_combout ;
wire \Selector595~0_combout ;
wire \Selector422~0_combout ;
wire \Selector422~2_combout ;
wire \Selector422~3_combout ;
wire \ac_state.s_0~q ;
wire \Selector433~0_combout ;
wire \addr_cmd~14_combout ;
wire \stage_counter[17]~2_combout ;
wire \stage_counter[17]~3_combout ;
wire \Selector448~0_combout ;
wire \Selector452~0_combout ;
wire \Selector472~2_combout ;
wire \Selector452~1_combout ;
wire \Selector452~2_combout ;
wire \Selector450~0_combout ;
wire \Selector450~1_combout ;
wire \Selector421~0_combout ;
wire \addr_cmd~57_combout ;
wire \Selector453~1_combout ;
wire \Add3~1_sumout ;
wire \Selector454~0_combout ;
wire \addr_cmd~7_combout ;
wire \Selector454~1_combout ;
wire \WideNor2~combout ;
wire \Selector595~3_combout ;
wire \Selector454~2_combout ;
wire \Selector454~3_combout ;
wire \Selector454~4_combout ;
wire \Selector454~5_combout ;
wire \stage_counter~37_combout ;
wire \stage_counter[0]~q ;
wire \Add3~2 ;
wire \Add3~5_sumout ;
wire \stage_counter~4_combout ;
wire \stage_counter[1]~q ;
wire \Add3~6 ;
wire \Add3~9_sumout ;
wire \stage_counter~5_combout ;
wire \stage_counter[2]~q ;
wire \Selector448~1_combout ;
wire \Selector451~0_combout ;
wire \Selector451~1_combout ;
wire \Add3~10 ;
wire \Add3~13_sumout ;
wire \stage_counter~6_combout ;
wire \stage_counter[3]~q ;
wire \Selector449~0_combout ;
wire \Selector449~1_combout ;
wire \Add3~14 ;
wire \Add3~17_sumout ;
wire \stage_counter~8_combout ;
wire \stage_counter[4]~q ;
wire \Add3~18 ;
wire \Add3~21_sumout ;
wire \stage_counter~7_combout ;
wire \stage_counter[5]~q ;
wire \stage_counter_zero~0_combout ;
wire \stage_counter[17]~9_combout ;
wire \stage_counter[17]~10_combout ;
wire \stage_counter[17]~11_combout ;
wire \stage_counter[17]~12_combout ;
wire \stage_counter[17]~18_combout ;
wire \Add3~22 ;
wire \Add3~25_sumout ;
wire \stage_counter~27_combout ;
wire \stage_counter[6]~q ;
wire \Add3~26 ;
wire \Add3~29_sumout ;
wire \stage_counter[8]~14_combout ;
wire \stage_counter~28_combout ;
wire \stage_counter~29_combout ;
wire \stage_counter[7]~q ;
wire \Add3~30 ;
wire \Add3~33_sumout ;
wire \stage_counter[8]~13_combout ;
wire \stage_counter~15_combout ;
wire \stage_counter~30_combout ;
wire \stage_counter~31_combout ;
wire \stage_counter[8]~q ;
wire \Add3~34 ;
wire \Add3~37_sumout ;
wire \stage_counter~32_combout ;
wire \stage_counter[9]~q ;
wire \Add3~38 ;
wire \Add3~41_sumout ;
wire \stage_counter~35_combout ;
wire \stage_counter~36_combout ;
wire \stage_counter[10]~q ;
wire \Add3~42 ;
wire \Add3~45_sumout ;
wire \stage_counter~33_combout ;
wire \stage_counter~34_combout ;
wire \stage_counter[11]~q ;
wire \Add3~46 ;
wire \Add3~49_sumout ;
wire \stage_counter~16_combout ;
wire \stage_counter~17_combout ;
wire \stage_counter[12]~q ;
wire \stage_counter~19_combout ;
wire \stage_counter~20_combout ;
wire \Add3~50 ;
wire \Add3~53_sumout ;
wire \stage_counter~21_combout ;
wire \stage_counter[13]~q ;
wire \Add3~54 ;
wire \Add3~57_sumout ;
wire \stage_counter~22_combout ;
wire \stage_counter[14]~q ;
wire \Add3~58 ;
wire \Add3~61_sumout ;
wire \stage_counter~23_combout ;
wire \stage_counter[17]~24_combout ;
wire \stage_counter[15]~q ;
wire \Add3~62 ;
wire \Add3~65_sumout ;
wire \stage_counter~26_combout ;
wire \stage_counter[16]~q ;
wire \Add3~66 ;
wire \Add3~69_sumout ;
wire \stage_counter~25_combout ;
wire \stage_counter[17]~q ;
wire \stage_counter_zero~1_combout ;
wire \stage_counter_zero~2_combout ;
wire \stage_counter_zero~3_combout ;
wire \stage_counter_zero~q ;
wire \stage_counter~0_combout ;
wire \Selector595~1_combout ;
wire \Selector595~2_combout ;
wire \finished_state~0_combout ;
wire \finished_state~q ;
wire \state~49_combout ;
wire \state.s_refresh_done~q ;
wire \Selector453~0_combout ;
wire \refresh_done~0_combout ;
wire \refresh_done~q ;
wire \initial_refresh_issued~0_combout ;
wire \initial_refresh_issued~q ;
wire \refresh_count[6]~0_combout ;
wire \refresh_count[6]~1_combout ;
wire \refresh_count~2_combout ;
wire \refresh_count[4]~q ;
wire \process_7~0_combout ;
wire \refresh_due~q ;
wire \num_stacked_refreshes~2_combout ;
wire \num_stacked_refreshes[0]~q ;
wire \num_stacked_refreshes~0_combout ;
wire \num_stacked_refreshes[2]~q ;
wire \num_stacked_refreshes~1_combout ;
wire \num_stacked_refreshes[1]~q ;
wire \LessThan0~0_combout ;
wire \refreshes_maxed~q ;
wire \state~35_combout ;
wire \state~57_combout ;
wire \state~58_combout ;
wire \state~59_combout ;
wire \state~60_combout ;
wire \state.s_idle~q ;
wire \state~62_combout ;
wire \state~37_combout ;
wire \state~39_combout ;
wire \state.s_run_init_seq~q ;
wire \command_done~0_combout ;
wire \command_done~q ;
wire \addr_cmd~0_combout ;
wire \addr_cmd~1_combout ;
wire \addr_cmd~2_combout ;
wire \addr_cmd~3_combout ;
wire \WideOr21~combout ;
wire \addr_cmd~4_combout ;
wire \addr_cmd~5_combout ;
wire \addr_cmd~6_combout ;
wire \addr_cmd~8_combout ;
wire \addr_cmd~9_combout ;
wire \addr_cmd~10_combout ;
wire \addr_cmd~11_combout ;
wire \addr_cmd~12_combout ;
wire \addr_cmd~13_combout ;
wire \addr_cmd~15_combout ;
wire \Selector468~0_combout ;
wire \Selector469~0_combout ;
wire \Selector468~1_combout ;
wire \Selector468~2_combout ;
wire \Selector469~1_combout ;
wire \Selector469~2_combout ;
wire \Selector469~3_combout ;
wire \addr_cmd~16_combout ;
wire \addr_cmd~17_combout ;
wire \addr_cmd~18_combout ;
wire \addr_cmd~19_combout ;
wire \addr_cmd~20_combout ;
wire \addr_cmd~21_combout ;
wire \Selector468~3_combout ;
wire \Selector468~4_combout ;
wire \addr_cmd~22_combout ;
wire \addr_cmd~23_combout ;
wire \addr_cmd~24_combout ;
wire \Selector469~4_combout ;
wire \Selector461~0_combout ;
wire \addr_cmd~25_combout ;
wire \addr_cmd~26_combout ;
wire \addr_cmd~27_combout ;
wire \Selector459~0_combout ;
wire \Selector459~1_combout ;
wire \Selector459~2_combout ;
wire \Selector459~3_combout ;
wire \addr_cmd~28_combout ;
wire \addr_cmd~29_combout ;
wire \addr_cmd~30_combout ;
wire \addr_cmd~31_combout ;
wire \addr_cmd~32_combout ;
wire \Selector472~0_combout ;
wire \Selector472~1_combout ;
wire \addr_cmd~33_combout ;
wire \addr_cmd~34_combout ;
wire \Selector471~0_combout ;
wire \Selector471~1_combout ;
wire \Selector471~2_combout ;
wire \addr_cmd~35_combout ;
wire \addr_cmd~36_combout ;
wire \addr_cmd~37_combout ;
wire \addr_cmd~38_combout ;
wire \addr_cmd~39_combout ;
wire \addr_cmd~40_combout ;
wire \addr_cmd~41_combout ;
wire \addr_cmd~42_combout ;
wire \addr_cmd~43_combout ;
wire \addr_cmd~44_combout ;
wire \addr_cmd~45_combout ;
wire \addr_cmd~46_combout ;
wire \addr_cmd~47_combout ;
wire \addr_cmd~48_combout ;
wire \addr_cmd~49_combout ;
wire \addr_cmd~50_combout ;
wire \addr_cmd~51_combout ;
wire \Selector473~0_combout ;
wire \Selector473~1_combout ;
wire \Selector473~2_combout ;
wire \Selector473~3_combout ;
wire \Selector473~4_combout ;
wire \addr_cmd~52_combout ;
wire \addr_cmd~53_combout ;
wire \addr_cmd~54_combout ;
wire \addr_cmd~55_combout ;
wire \addr_cmd~56_combout ;
wire \addr_cmd~58_combout ;
wire \addr_cmd~59_combout ;
wire \addr_cmd~60_combout ;
wire \addr_cmd~61_combout ;
wire \addr_cmd~62_combout ;
wire \addr_cmd~63_combout ;
wire \addr_cmd~64_combout ;
wire \addr_cmd~65_combout ;
wire \addr_cmd~66_combout ;
wire \addr_cmd~67_combout ;
wire \addr_cmd~68_combout ;


arriaii_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\refresh_count[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "off";

arriaii_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\refresh_count[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000000000FF00;
defparam \Add0~5 .shared_arith = "off";

arriaii_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\refresh_count[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000000000FF00;
defparam \Add0~9 .shared_arith = "off";

arriaii_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\refresh_count[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

arriaii_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\refresh_count[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \admin_ctrl.command_done (
	.clk(clk),
	.d(\command_done~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(admin_ctrlcommand_done),
	.prn(vcc));
defparam \admin_ctrl.command_done .is_wysiwyg = "true";
defparam \admin_ctrl.command_done .power_up = "low";

dffeas ac_access_gnt(
	.clk(clk),
	.d(\state.s_access~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ac_access_gnt1),
	.prn(vcc));
defparam ac_access_gnt.is_wysiwyg = "true";
defparam ac_access_gnt.power_up = "low";

dffeas seq_ac_sel(
	.clk(clk),
	.d(\cal_complete~combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_ac_sel1),
	.prn(vcc));
defparam seq_ac_sel.is_wysiwyg = "true";
defparam seq_ac_sel.power_up = "low";

dffeas \addr_cmd[0].cs_n[0] (
	.clk(clk),
	.d(\addr_cmd~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd0cs_n0),
	.prn(vcc));
defparam \addr_cmd[0].cs_n[0] .is_wysiwyg = "true";
defparam \addr_cmd[0].cs_n[0] .power_up = "low";

dffeas \addr_cmd[1].cs_n[0] (
	.clk(clk),
	.d(\addr_cmd~9_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd1cs_n0),
	.prn(vcc));
defparam \addr_cmd[1].cs_n[0] .is_wysiwyg = "true";
defparam \addr_cmd[1].cs_n[0] .power_up = "low";

dffeas \addr_cmd[0].cke[0] (
	.clk(clk),
	.d(\addr_cmd~12_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd0cke0),
	.prn(vcc));
defparam \addr_cmd[0].cke[0] .is_wysiwyg = "true";
defparam \addr_cmd[0].cke[0] .power_up = "low";

dffeas \addr_cmd[0].addr[0] (
	.clk(clk),
	.d(\addr_cmd~16_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd0addr0),
	.prn(vcc));
defparam \addr_cmd[0].addr[0] .is_wysiwyg = "true";
defparam \addr_cmd[0].addr[0] .power_up = "low";

dffeas \addr_cmd[1].addr[0] (
	.clk(clk),
	.d(\addr_cmd~20_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd1addr0),
	.prn(vcc));
defparam \addr_cmd[1].addr[0] .is_wysiwyg = "true";
defparam \addr_cmd[1].addr[0] .power_up = "low";

dffeas \addr_cmd[0].addr[1] (
	.clk(clk),
	.d(\addr_cmd~22_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd0addr1),
	.prn(vcc));
defparam \addr_cmd[0].addr[1] .is_wysiwyg = "true";
defparam \addr_cmd[0].addr[1] .power_up = "low";

dffeas \addr_cmd[1].addr[1] (
	.clk(clk),
	.d(\addr_cmd~23_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd1addr1),
	.prn(vcc));
defparam \addr_cmd[1].addr[1] .is_wysiwyg = "true";
defparam \addr_cmd[1].addr[1] .power_up = "low";

dffeas \addr_cmd[0].addr[8] (
	.clk(clk),
	.d(\addr_cmd~25_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd0addr8),
	.prn(vcc));
defparam \addr_cmd[0].addr[8] .is_wysiwyg = "true";
defparam \addr_cmd[0].addr[8] .power_up = "low";

dffeas \addr_cmd[1].addr[8] (
	.clk(clk),
	.d(\addr_cmd~26_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd1addr8),
	.prn(vcc));
defparam \addr_cmd[1].addr[8] .is_wysiwyg = "true";
defparam \addr_cmd[1].addr[8] .power_up = "low";

dffeas \addr_cmd[0].addr[10] (
	.clk(clk),
	.d(\addr_cmd~28_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd0addr10),
	.prn(vcc));
defparam \addr_cmd[0].addr[10] .is_wysiwyg = "true";
defparam \addr_cmd[0].addr[10] .power_up = "low";

dffeas \addr_cmd[1].addr[10] (
	.clk(clk),
	.d(\addr_cmd~31_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd1addr10),
	.prn(vcc));
defparam \addr_cmd[1].addr[10] .is_wysiwyg = "true";
defparam \addr_cmd[1].addr[10] .power_up = "low";

dffeas \addr_cmd[0].ba[0] (
	.clk(clk),
	.d(\addr_cmd~33_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd0ba0),
	.prn(vcc));
defparam \addr_cmd[0].ba[0] .is_wysiwyg = "true";
defparam \addr_cmd[0].ba[0] .power_up = "low";

dffeas \addr_cmd[1].ba[0] (
	.clk(clk),
	.d(\addr_cmd~34_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd1ba0),
	.prn(vcc));
defparam \addr_cmd[1].ba[0] .is_wysiwyg = "true";
defparam \addr_cmd[1].ba[0] .power_up = "low";

dffeas \addr_cmd[0].ba[1] (
	.clk(clk),
	.d(\addr_cmd~35_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd0ba1),
	.prn(vcc));
defparam \addr_cmd[0].ba[1] .is_wysiwyg = "true";
defparam \addr_cmd[0].ba[1] .power_up = "low";

dffeas \addr_cmd[1].ba[1] (
	.clk(clk),
	.d(\addr_cmd~36_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd1ba1),
	.prn(vcc));
defparam \addr_cmd[1].ba[1] .is_wysiwyg = "true";
defparam \addr_cmd[1].ba[1] .power_up = "low";

dffeas \addr_cmd[0].ras_n (
	.clk(clk),
	.d(\addr_cmd~47_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd0ras_n),
	.prn(vcc));
defparam \addr_cmd[0].ras_n .is_wysiwyg = "true";
defparam \addr_cmd[0].ras_n .power_up = "low";

dffeas \addr_cmd[1].ras_n (
	.clk(clk),
	.d(\addr_cmd~50_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd1ras_n),
	.prn(vcc));
defparam \addr_cmd[1].ras_n .is_wysiwyg = "true";
defparam \addr_cmd[1].ras_n .power_up = "low";

dffeas \addr_cmd[0].cas_n (
	.clk(clk),
	.d(\addr_cmd~52_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd0cas_n),
	.prn(vcc));
defparam \addr_cmd[0].cas_n .is_wysiwyg = "true";
defparam \addr_cmd[0].cas_n .power_up = "low";

dffeas \addr_cmd[1].cas_n (
	.clk(clk),
	.d(\addr_cmd~56_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd1cas_n),
	.prn(vcc));
defparam \addr_cmd[1].cas_n .is_wysiwyg = "true";
defparam \addr_cmd[1].cas_n .power_up = "low";

dffeas \addr_cmd[0].we_n (
	.clk(clk),
	.d(\addr_cmd~63_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd0we_n),
	.prn(vcc));
defparam \addr_cmd[0].we_n .is_wysiwyg = "true";
defparam \addr_cmd[0].we_n .power_up = "low";

dffeas \addr_cmd[1].we_n (
	.clk(clk),
	.d(\addr_cmd~66_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd1we_n),
	.prn(vcc));
defparam \addr_cmd[1].we_n .is_wysiwyg = "true";
defparam \addr_cmd[1].we_n .power_up = "low";

dffeas \addr_cmd[0].rst_n (
	.clk(clk),
	.d(\addr_cmd~68_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(addr_cmd0rst_n),
	.prn(vcc));
defparam \addr_cmd[0].rst_n .is_wysiwyg = "true";
defparam \addr_cmd[0].rst_n .power_up = "low";

dffeas \admin_ctrl.command_ack (
	.clk(clk),
	.d(\command_started~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(admin_ctrlcommand_ack),
	.prn(vcc));
defparam \admin_ctrl.command_ack .is_wysiwyg = "true";
defparam \admin_ctrl.command_ack .power_up = "low";

arriaii_lcell_comb \refresh_count~10 (
	.dataa(!\Add0~13_sumout ),
	.datab(!\refresh_count[6]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\refresh_count~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \refresh_count~10 .extended_lut = "off";
defparam \refresh_count~10 .lut_mask = 64'h1111111111111111;
defparam \refresh_count~10 .shared_arith = "off";

dffeas \refresh_count[3] (
	.clk(clk),
	.d(\refresh_count~10_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_count[3]~q ),
	.prn(vcc));
defparam \refresh_count[3] .is_wysiwyg = "true";
defparam \refresh_count[3] .power_up = "low";

arriaii_lcell_comb \refresh_count~11 (
	.dataa(!\Add0~9_sumout ),
	.datab(!\refresh_count[6]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\refresh_count~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \refresh_count~11 .extended_lut = "off";
defparam \refresh_count~11 .lut_mask = 64'h2222222222222222;
defparam \refresh_count~11 .shared_arith = "off";

dffeas \refresh_count[2] (
	.clk(clk),
	.d(\refresh_count~11_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_count[2]~q ),
	.prn(vcc));
defparam \refresh_count[2] .is_wysiwyg = "true";
defparam \refresh_count[2] .power_up = "low";

arriaii_lcell_comb \refresh_count~9 (
	.dataa(!\Add0~5_sumout ),
	.datab(!\refresh_count[6]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\refresh_count~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \refresh_count~9 .extended_lut = "off";
defparam \refresh_count~9 .lut_mask = 64'h2222222222222222;
defparam \refresh_count~9 .shared_arith = "off";

dffeas \refresh_count[1] (
	.clk(clk),
	.d(\refresh_count~9_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_count[1]~q ),
	.prn(vcc));
defparam \refresh_count[1] .is_wysiwyg = "true";
defparam \refresh_count[1] .power_up = "low";

arriaii_lcell_comb \refresh_count~8 (
	.dataa(!\Add0~1_sumout ),
	.datab(!\refresh_count[6]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\refresh_count~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \refresh_count~8 .extended_lut = "off";
defparam \refresh_count~8 .lut_mask = 64'h2222222222222222;
defparam \refresh_count~8 .shared_arith = "off";

dffeas \refresh_count[0] (
	.clk(clk),
	.d(\refresh_count~8_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_count[0]~q ),
	.prn(vcc));
defparam \refresh_count[0] .is_wysiwyg = "true";
defparam \refresh_count[0] .power_up = "low";

arriaii_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\refresh_count[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

arriaii_lcell_comb \refresh_count~3 (
	.dataa(!\refresh_count[6]~1_combout ),
	.datab(!\Add0~21_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\refresh_count~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \refresh_count~3 .extended_lut = "off";
defparam \refresh_count~3 .lut_mask = 64'h1111111111111111;
defparam \refresh_count~3 .shared_arith = "off";

dffeas \refresh_count[5] (
	.clk(clk),
	.d(\refresh_count~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_count[5]~q ),
	.prn(vcc));
defparam \refresh_count[5] .is_wysiwyg = "true";
defparam \refresh_count[5] .power_up = "low";

arriaii_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\refresh_count[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000000000FF00;
defparam \Add0~25 .shared_arith = "off";

arriaii_lcell_comb \refresh_count~4 (
	.dataa(!\refresh_count[6]~1_combout ),
	.datab(!\Add0~25_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\refresh_count~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \refresh_count~4 .extended_lut = "off";
defparam \refresh_count~4 .lut_mask = 64'h4444444444444444;
defparam \refresh_count~4 .shared_arith = "off";

dffeas \refresh_count[6] (
	.clk(clk),
	.d(\refresh_count~4_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_count[6]~q ),
	.prn(vcc));
defparam \refresh_count[6] .is_wysiwyg = "true";
defparam \refresh_count[6] .power_up = "low";

arriaii_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\refresh_count[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

arriaii_lcell_comb \refresh_count~5 (
	.dataa(!\refresh_count[6]~1_combout ),
	.datab(!\Add0~29_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\refresh_count~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \refresh_count~5 .extended_lut = "off";
defparam \refresh_count~5 .lut_mask = 64'h1111111111111111;
defparam \refresh_count~5 .shared_arith = "off";

dffeas \refresh_count[7] (
	.clk(clk),
	.d(\refresh_count~5_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_count[7]~q ),
	.prn(vcc));
defparam \refresh_count[7] .is_wysiwyg = "true";
defparam \refresh_count[7] .power_up = "low";

arriaii_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\refresh_count[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

arriaii_lcell_comb \refresh_count~7 (
	.dataa(!\refresh_count[6]~1_combout ),
	.datab(!\Add0~33_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\refresh_count~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \refresh_count~7 .extended_lut = "off";
defparam \refresh_count~7 .lut_mask = 64'h1111111111111111;
defparam \refresh_count~7 .shared_arith = "off";

dffeas \refresh_count[8] (
	.clk(clk),
	.d(\refresh_count~7_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_count[8]~q ),
	.prn(vcc));
defparam \refresh_count[8] .is_wysiwyg = "true";
defparam \refresh_count[8] .power_up = "low";

arriaii_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\refresh_count[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000000000FF00;
defparam \Add0~37 .shared_arith = "off";

arriaii_lcell_comb \refresh_count~6 (
	.dataa(!\refresh_count[6]~1_combout ),
	.datab(!\Add0~37_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\refresh_count~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \refresh_count~6 .extended_lut = "off";
defparam \refresh_count~6 .lut_mask = 64'h4444444444444444;
defparam \refresh_count~6 .shared_arith = "off";

dffeas \refresh_count[9] (
	.clk(clk),
	.d(\refresh_count~6_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_count[9]~q ),
	.prn(vcc));
defparam \refresh_count[9] .is_wysiwyg = "true";
defparam \refresh_count[9] .power_up = "low";

arriaii_lcell_comb \Equal0~0 (
	.dataa(!\refresh_count[6]~q ),
	.datab(!\refresh_count[7]~q ),
	.datac(!\refresh_count[9]~q ),
	.datad(!\refresh_count[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h0400040004000400;
defparam \Equal0~0 .shared_arith = "off";

arriaii_lcell_comb \Equal0~1 (
	.dataa(!\refresh_count[0]~q ),
	.datab(!\refresh_count[1]~q ),
	.datac(!\refresh_count[3]~q ),
	.datad(!\refresh_count[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~1 .extended_lut = "off";
defparam \Equal0~1 .lut_mask = 64'h0010001000100010;
defparam \Equal0~1 .shared_arith = "off";

arriaii_lcell_comb \state~38 (
	.dataa(!\state.s_access~q ),
	.datab(!ctl_init_fail),
	.datac(!ctl_init_success),
	.datad(!dgrb_ac_access_req),
	.datae(!dgwb_ac_access_req),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~38 .extended_lut = "off";
defparam \state~38 .lut_mask = 64'h80C0C08080C0C080;
defparam \state~38 .shared_arith = "off";

arriaii_lcell_comb \state.s_reset~0 (
	.dataa(!\state.s_reset~q ),
	.datab(!\state~62_combout ),
	.datac(!\state~38_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state.s_reset~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state.s_reset~0 .extended_lut = "off";
defparam \state.s_reset~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \state.s_reset~0 .shared_arith = "off";

dffeas \state.s_reset (
	.clk(clk),
	.d(\state.s_reset~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_reset~q ),
	.prn(vcc));
defparam \state.s_reset .is_wysiwyg = "true";
defparam \state.s_reset .power_up = "low";

arriaii_lcell_comb \WideOr34~0 (
	.dataa(!\state.s_access~q ),
	.datab(!\state.s_reset~q ),
	.datac(!\state.s_idle~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr34~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr34~0 .extended_lut = "off";
defparam \WideOr34~0 .lut_mask = 64'h2020202020202020;
defparam \WideOr34~0 .shared_arith = "off";

arriaii_lcell_comb \Selector431~0 (
	.dataa(!\ac_state.s_8~q ),
	.datab(!\ac_state.s_9~q ),
	.datac(!\WideOr34~0_combout ),
	.datad(!\Selector433~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector431~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector431~0 .extended_lut = "off";
defparam \Selector431~0 .lut_mask = 64'h3075307530753075;
defparam \Selector431~0 .shared_arith = "off";

dffeas \ac_state.s_9 (
	.clk(clk),
	.d(\Selector431~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\stage_counter~0_combout ),
	.q(\ac_state.s_9~q ),
	.prn(vcc));
defparam \ac_state.s_9 .is_wysiwyg = "true";
defparam \ac_state.s_9 .power_up = "low";

arriaii_lcell_comb \Selector432~0 (
	.dataa(!\ac_state.s_10~q ),
	.datab(!\ac_state.s_9~q ),
	.datac(!\WideOr34~0_combout ),
	.datad(!\Selector433~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector432~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector432~0 .extended_lut = "off";
defparam \Selector432~0 .lut_mask = 64'h5073507350735073;
defparam \Selector432~0 .shared_arith = "off";

dffeas \ac_state.s_10 (
	.clk(clk),
	.d(\Selector432~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\stage_counter~0_combout ),
	.q(\ac_state.s_10~q ),
	.prn(vcc));
defparam \ac_state.s_10 .is_wysiwyg = "true";
defparam \ac_state.s_10 .power_up = "low";

arriaii_lcell_comb \Selector433~1 (
	.dataa(!\ac_state.s_11~q ),
	.datab(!\ac_state.s_10~q ),
	.datac(!\WideOr34~0_combout ),
	.datad(!\Selector433~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector433~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector433~1 .extended_lut = "off";
defparam \Selector433~1 .lut_mask = 64'h5073507350735073;
defparam \Selector433~1 .shared_arith = "off";

dffeas \ac_state.s_11 (
	.clk(clk),
	.d(\Selector433~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\stage_counter~0_combout ),
	.q(\ac_state.s_11~q ),
	.prn(vcc));
defparam \ac_state.s_11 .is_wysiwyg = "true";
defparam \ac_state.s_11 .power_up = "low";

arriaii_lcell_comb \Selector434~0 (
	.dataa(!\state.s_run_init_seq~q ),
	.datab(!\ac_state.s_12~q ),
	.datac(!\ac_state.s_11~q ),
	.datad(!\WideOr34~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector434~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector434~0 .extended_lut = "off";
defparam \Selector434~0 .lut_mask = 64'h3705370537053705;
defparam \Selector434~0 .shared_arith = "off";

dffeas \ac_state.s_12 (
	.clk(clk),
	.d(\Selector434~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\stage_counter~0_combout ),
	.q(\ac_state.s_12~q ),
	.prn(vcc));
defparam \ac_state.s_12 .is_wysiwyg = "true";
defparam \ac_state.s_12 .power_up = "low";

arriaii_lcell_comb \Selector3~0 (
	.dataa(!curr_cmdcmd_init_dram),
	.datab(!\admin_req_extended~q ),
	.datac(!\state.s_reset~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'hE0E0E0E0E0E0E0E0;
defparam \Selector3~0 .shared_arith = "off";

arriaii_lcell_comb \state~43 (
	.dataa(!curr_cmdcmd_init_dram),
	.datab(!\finished_state~q ),
	.datac(!\admin_req_extended~q ),
	.datad(!\state.s_reset~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~43 .extended_lut = "off";
defparam \state~43 .lut_mask = 64'h0133013301330133;
defparam \state~43 .shared_arith = "off";

arriaii_lcell_comb \state~50 (
	.dataa(!curr_cmdcmd_prep_customer_mr_setup),
	.datab(!dgb_ac_access_req),
	.datac(!\admin_req_extended~q ),
	.datad(!\state.s_idle~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~50_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~50 .extended_lut = "off";
defparam \state~50 .lut_mask = 64'h0037003700370037;
defparam \state~50 .shared_arith = "off";

arriaii_lcell_comb \state~36 (
	.dataa(!dgb_ac_access_req),
	.datab(!\state.s_idle~q ),
	.datac(!\state~35_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~36 .extended_lut = "off";
defparam \state~36 .lut_mask = 64'h3131313131313131;
defparam \state~36 .shared_arith = "off";

arriaii_lcell_comb \state~40 (
	.dataa(!curr_cmdcmd_prog_cal_mr),
	.datab(!dgb_ac_access_req),
	.datac(!\admin_req_extended~q ),
	.datad(!\state~36_combout ),
	.datae(!\state~38_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~40 .extended_lut = "off";
defparam \state~40 .lut_mask = 64'h0000000400000004;
defparam \state~40 .shared_arith = "off";

arriaii_lcell_comb \state~41 (
	.dataa(!\finished_state~q ),
	.datab(!\state~38_combout ),
	.datac(!dgb_ac_access_req),
	.datad(!\state.s_idle~q ),
	.datae(!\state~35_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~41 .extended_lut = "off";
defparam \state~41 .lut_mask = 64'hDDFFDDDFDDFFDDDF;
defparam \state~41 .shared_arith = "off";

dffeas \state.s_program_cal_mrs (
	.clk(clk),
	.d(\state~40_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state~41_combout ),
	.q(\state.s_program_cal_mrs~q ),
	.prn(vcc));
defparam \state.s_program_cal_mrs .is_wysiwyg = "true";
defparam \state.s_program_cal_mrs .power_up = "low";

arriaii_lcell_comb \ac_state~19 (
	.dataa(!\state.s_access~q ),
	.datab(!\state.s_reset~q ),
	.datac(!\stage_counter_zero~q ),
	.datad(!\state.s_idle~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_state~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_state~19 .extended_lut = "off";
defparam \ac_state~19 .lut_mask = 64'h2000200020002000;
defparam \ac_state~19 .shared_arith = "off";

arriaii_lcell_comb \stage_counter[17]~1 (
	.dataa(!\state.s_program_cal_mrs~q ),
	.datab(!\state.s_prog_user_mrs~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter[17]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter[17]~1 .extended_lut = "off";
defparam \stage_counter[17]~1 .lut_mask = 64'h8888888888888888;
defparam \stage_counter[17]~1 .shared_arith = "off";

arriaii_lcell_comb \process_12~0 (
	.dataa(!\ac_state.s_12~q ),
	.datab(!\ac_state.s_0~q ),
	.datac(!\ac_state.s_11~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\process_12~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \process_12~0 .extended_lut = "off";
defparam \process_12~0 .lut_mask = 64'h2020202020202020;
defparam \process_12~0 .shared_arith = "off";

arriaii_lcell_comb \ac_state~20 (
	.dataa(!\state.s_run_init_seq~q ),
	.datab(!\stage_counter[17]~1_combout ),
	.datac(!\process_12~0_combout ),
	.datad(!\ac_state~19_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_state~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_state~20 .extended_lut = "off";
defparam \ac_state~20 .lut_mask = 64'h0072007200720072;
defparam \ac_state~20 .shared_arith = "off";

arriaii_lcell_comb \ac_state~24 (
	.dataa(!\ac_state.s_2~q ),
	.datab(!\ac_state.s_3~q ),
	.datac(!\ac_state~19_combout ),
	.datad(!\ac_state~20_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_state~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_state~24 .extended_lut = "off";
defparam \ac_state~24 .lut_mask = 64'h3500350035003500;
defparam \ac_state~24 .shared_arith = "off";

dffeas \ac_state.s_3 (
	.clk(clk),
	.d(\ac_state~24_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_state.s_3~q ),
	.prn(vcc));
defparam \ac_state.s_3 .is_wysiwyg = "true";
defparam \ac_state.s_3 .power_up = "low";

arriaii_lcell_comb \ac_state~23 (
	.dataa(!\ac_state.s_4~q ),
	.datab(!\ac_state.s_3~q ),
	.datac(!\ac_state~19_combout ),
	.datad(!\ac_state~20_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_state~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_state~23 .extended_lut = "off";
defparam \ac_state~23 .lut_mask = 64'h5300530053005300;
defparam \ac_state~23 .shared_arith = "off";

dffeas \ac_state.s_4 (
	.clk(clk),
	.d(\ac_state~23_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_state.s_4~q ),
	.prn(vcc));
defparam \ac_state.s_4 .is_wysiwyg = "true";
defparam \ac_state.s_4 .power_up = "low";

arriaii_lcell_comb \ac_state~22 (
	.dataa(!\ac_state.s_5~q ),
	.datab(!\ac_state.s_4~q ),
	.datac(!\ac_state~19_combout ),
	.datad(!\ac_state~20_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_state~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_state~22 .extended_lut = "off";
defparam \ac_state~22 .lut_mask = 64'h5300530053005300;
defparam \ac_state~22 .shared_arith = "off";

dffeas \ac_state.s_5 (
	.clk(clk),
	.d(\ac_state~22_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_state.s_5~q ),
	.prn(vcc));
defparam \ac_state.s_5 .is_wysiwyg = "true";
defparam \ac_state.s_5 .power_up = "low";

arriaii_lcell_comb WideOr32(
	.dataa(!\state.s_access~q ),
	.datab(!\state.s_idle~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr32~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr32.extended_lut = "off";
defparam WideOr32.lut_mask = 64'h8888888888888888;
defparam WideOr32.shared_arith = "off";

arriaii_lcell_comb \Selector421~1 (
	.dataa(!\state.s_run_init_seq~q ),
	.datab(!\state.s_program_cal_mrs~q ),
	.datac(!\ac_state.s_5~q ),
	.datad(!\WideOr32~combout ),
	.datae(!\per_cs_init_seen[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector421~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector421~1 .extended_lut = "off";
defparam \Selector421~1 .lut_mask = 64'h0303FFBB0303FFBB;
defparam \Selector421~1 .shared_arith = "off";

dffeas \per_cs_init_seen[0] (
	.clk(clk),
	.d(\Selector421~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\stage_counter~0_combout ),
	.q(\per_cs_init_seen[0]~q ),
	.prn(vcc));
defparam \per_cs_init_seen[0] .is_wysiwyg = "true";
defparam \per_cs_init_seen[0] .power_up = "low";

dffeas mem_init_complete(
	.clk(clk),
	.d(\per_cs_init_seen[0]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_init_complete~q ),
	.prn(vcc));
defparam mem_init_complete.is_wysiwyg = "true";
defparam mem_init_complete.power_up = "low";

arriaii_lcell_comb \state~51 (
	.dataa(!\finished_state~q ),
	.datab(!\state.s_program_cal_mrs~q ),
	.datac(!\state.s_topup_refresh_done~q ),
	.datad(!\refreshes_maxed~q ),
	.datae(!\mem_init_complete~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~51 .extended_lut = "off";
defparam \state~51 .lut_mask = 64'h0500150005001500;
defparam \state~51 .shared_arith = "off";

arriaii_lcell_comb \state~52 (
	.dataa(!\cal_complete~combout ),
	.datab(!\state.s_topup_refresh~q ),
	.datac(!\state~43_combout ),
	.datad(!\state~50_combout ),
	.datae(!\state~51_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~52 .extended_lut = "off";
defparam \state~52 .lut_mask = 64'h20AAAAAA20AAAAAA;
defparam \state~52 .shared_arith = "off";

dffeas \state.s_topup_refresh (
	.clk(clk),
	.d(\state~52_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_topup_refresh~q ),
	.prn(vcc));
defparam \state.s_topup_refresh .is_wysiwyg = "true";
defparam \state.s_topup_refresh .power_up = "low";

arriaii_lcell_comb \state~48 (
	.dataa(!\cal_complete~combout ),
	.datab(!\finished_state~q ),
	.datac(!\Selector3~0_combout ),
	.datad(!\state.s_topup_refresh_done~q ),
	.datae(!\state.s_topup_refresh~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~48 .extended_lut = "off";
defparam \state~48 .lut_mask = 64'h008A22AA008A22AA;
defparam \state~48 .shared_arith = "off";

dffeas \state.s_topup_refresh_done (
	.clk(clk),
	.d(\state~48_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_topup_refresh_done~q ),
	.prn(vcc));
defparam \state.s_topup_refresh_done .is_wysiwyg = "true";
defparam \state.s_topup_refresh_done .power_up = "low";

arriaii_lcell_comb \state~42 (
	.dataa(!curr_cmdcmd_prep_customer_mr_setup),
	.datab(!\finished_state~q ),
	.datac(!\state.s_topup_refresh_done~q ),
	.datad(!\refreshes_maxed~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~42 .extended_lut = "off";
defparam \state~42 .lut_mask = 64'h0001000100010001;
defparam \state~42 .shared_arith = "off";

arriaii_lcell_comb \Selector15~0 (
	.dataa(!\state.s_idle~q ),
	.datab(!dgb_ac_access_req),
	.datac(!\state.s_reset~q ),
	.datad(!\state~42_combout ),
	.datae(!curr_cmdcmd_init_dram),
	.dataf(!\admin_req_extended~q ),
	.datag(!curr_cmdcmd_prog_cal_mr),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector15~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector15~0 .extended_lut = "on";
defparam \Selector15~0 .lut_mask = 64'h0000000004FFF4FF;
defparam \Selector15~0 .shared_arith = "off";

dffeas command_started(
	.clk(clk),
	.d(\Selector15~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\command_started~q ),
	.prn(vcc));
defparam command_started.is_wysiwyg = "true";
defparam command_started.power_up = "low";

arriaii_lcell_comb \admin_req_extended~0 (
	.dataa(!WideOr0),
	.datab(!ac_muxctrl_broadcast_rcommand_req),
	.datac(!\admin_req_extended~q ),
	.datad(!\command_started~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\admin_req_extended~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \admin_req_extended~0 .extended_lut = "off";
defparam \admin_req_extended~0 .lut_mask = 64'h2F222F222F222F22;
defparam \admin_req_extended~0 .shared_arith = "off";

dffeas admin_req_extended(
	.clk(clk),
	.d(\admin_req_extended~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\admin_req_extended~q ),
	.prn(vcc));
defparam admin_req_extended.is_wysiwyg = "true";
defparam admin_req_extended.power_up = "low";

arriaii_lcell_comb \state~44 (
	.dataa(!\cal_complete~combout ),
	.datab(!\state.s_prog_user_mrs~q ),
	.datac(!\admin_req_extended~q ),
	.datad(!\state~42_combout ),
	.datae(!\state~43_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~44 .extended_lut = "off";
defparam \state~44 .lut_mask = 64'h222A000A222A000A;
defparam \state~44 .shared_arith = "off";

dffeas \state.s_prog_user_mrs (
	.clk(clk),
	.d(\state~44_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_prog_user_mrs~q ),
	.prn(vcc));
defparam \state.s_prog_user_mrs .is_wysiwyg = "true";
defparam \state.s_prog_user_mrs .power_up = "low";

arriaii_lcell_comb \ac_state~21 (
	.dataa(!\ac_state.s_6~q ),
	.datab(!\ac_state.s_5~q ),
	.datac(!\ac_state~19_combout ),
	.datad(!\ac_state~20_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_state~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_state~21 .extended_lut = "off";
defparam \ac_state~21 .lut_mask = 64'h5300530053005300;
defparam \ac_state~21 .shared_arith = "off";

dffeas \ac_state.s_6 (
	.clk(clk),
	.d(\ac_state~21_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_state.s_6~q ),
	.prn(vcc));
defparam \ac_state.s_6 .is_wysiwyg = "true";
defparam \ac_state.s_6 .power_up = "low";

arriaii_lcell_comb \Selector429~0 (
	.dataa(!\state.s_run_init_seq~q ),
	.datab(!\state.s_prog_user_mrs~q ),
	.datac(!\ac_state.s_6~q ),
	.datad(!\ac_state.s_7~q ),
	.datae(!\WideOr34~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector429~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector429~0 .extended_lut = "off";
defparam \Selector429~0 .lut_mask = 64'h07FF070707FF0707;
defparam \Selector429~0 .shared_arith = "off";

dffeas \ac_state.s_7 (
	.clk(clk),
	.d(\Selector429~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\stage_counter~0_combout ),
	.q(\ac_state.s_7~q ),
	.prn(vcc));
defparam \ac_state.s_7 .is_wysiwyg = "true";
defparam \ac_state.s_7 .power_up = "low";

arriaii_lcell_comb \Selector430~0 (
	.dataa(!\ac_state.s_7~q ),
	.datab(!\ac_state.s_8~q ),
	.datac(!\WideOr34~0_combout ),
	.datad(!\Selector433~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector430~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector430~0 .extended_lut = "off";
defparam \Selector430~0 .lut_mask = 64'h3075307530753075;
defparam \Selector430~0 .shared_arith = "off";

dffeas \ac_state.s_8 (
	.clk(clk),
	.d(\Selector430~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\stage_counter~0_combout ),
	.q(\ac_state.s_8~q ),
	.prn(vcc));
defparam \ac_state.s_8 .is_wysiwyg = "true";
defparam \ac_state.s_8 .power_up = "low";

arriaii_lcell_comb WideOr16(
	.dataa(!\ac_state.s_12~q ),
	.datab(!\ac_state.s_11~q ),
	.datac(!\ac_state.s_10~q ),
	.datad(!\ac_state.s_8~q ),
	.datae(!\ac_state.s_9~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr16~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr16.extended_lut = "off";
defparam WideOr16.lut_mask = 64'h8000000080000000;
defparam WideOr16.shared_arith = "off";

arriaii_lcell_comb \ac_state.s_1~0 (
	.dataa(!\ac_state.s_1~q ),
	.datab(!\ac_state.s_0~q ),
	.datac(!\ac_state~19_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_state.s_1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_state.s_1~0 .extended_lut = "off";
defparam \ac_state.s_1~0 .lut_mask = 64'h5C5C5C5C5C5C5C5C;
defparam \ac_state.s_1~0 .shared_arith = "off";

dffeas \ac_state.s_1 (
	.clk(clk),
	.d(\ac_state.s_1~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_state.s_1~q ),
	.prn(vcc));
defparam \ac_state.s_1 .is_wysiwyg = "true";
defparam \ac_state.s_1 .power_up = "low";

arriaii_lcell_comb cal_complete(
	.dataa(!ctl_init_fail),
	.datab(!ctl_init_success),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cal_complete~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam cal_complete.extended_lut = "off";
defparam cal_complete.lut_mask = 64'h7777777777777777;
defparam cal_complete.shared_arith = "off";

arriaii_lcell_comb \state~56 (
	.dataa(!curr_cmdcmd_prep_customer_mr_setup),
	.datab(!\finished_state~q ),
	.datac(!\admin_req_extended~q ),
	.datad(!\state.s_topup_refresh_done~q ),
	.datae(!\refreshes_maxed~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~56_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~56 .extended_lut = "off";
defparam \state~56 .lut_mask = 64'h0000003200000032;
defparam \state~56 .shared_arith = "off";

arriaii_lcell_comb \state~61 (
	.dataa(!\cal_complete~combout ),
	.datab(!dgb_ac_access_req),
	.datac(!\state.s_zq_cal_short~q ),
	.datad(!\state~43_combout ),
	.datae(!\state~56_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~61_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~61 .extended_lut = "off";
defparam \state~61 .lut_mask = 64'h0A002A220A002A22;
defparam \state~61 .shared_arith = "off";

dffeas \state.s_zq_cal_short (
	.clk(clk),
	.d(\state~61_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_zq_cal_short~q ),
	.prn(vcc));
defparam \state.s_zq_cal_short .is_wysiwyg = "true";
defparam \state.s_zq_cal_short .power_up = "low";

arriaii_lcell_comb \state~45 (
	.dataa(!\cal_complete~combout ),
	.datab(!\finished_state~q ),
	.datac(!\state.s_access_act~q ),
	.datad(!\Selector3~0_combout ),
	.datae(!\state.s_zq_cal_short~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~45 .extended_lut = "off";
defparam \state~45 .lut_mask = 64'h080A2A2A080A2A2A;
defparam \state~45 .shared_arith = "off";

dffeas \state.s_access_act (
	.clk(clk),
	.d(\state~45_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_access_act~q ),
	.prn(vcc));
defparam \state.s_access_act .is_wysiwyg = "true";
defparam \state.s_access_act .power_up = "low";

arriaii_lcell_comb \state~34 (
	.dataa(!\cal_complete~combout ),
	.datab(!\state.s_access~q ),
	.datac(!\finished_state~q ),
	.datad(!\state.s_access_act~q ),
	.datae(!dgb_ac_access_req),
	.dataf(!\Selector3~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~34 .extended_lut = "off";
defparam \state~34 .lut_mask = 64'h000A222A222A222A;
defparam \state~34 .shared_arith = "off";

dffeas \state.s_access (
	.clk(clk),
	.d(\state~34_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_access~q ),
	.prn(vcc));
defparam \state.s_access .is_wysiwyg = "true";
defparam \state.s_access .power_up = "low";

arriaii_lcell_comb \state~46 (
	.dataa(!WideOr0),
	.datab(!\cal_complete~combout ),
	.datac(!\state.s_access~q ),
	.datad(!\admin_req_extended~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~46 .extended_lut = "off";
defparam \state~46 .lut_mask = 64'hC040C040C040C040;
defparam \state~46 .shared_arith = "off";

arriaii_lcell_comb \state~47 (
	.dataa(!dgb_ac_access_req),
	.datab(!\state.s_idle~q ),
	.datac(!\state~35_combout ),
	.datad(!\state~46_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~47 .extended_lut = "off";
defparam \state~47 .lut_mask = 64'h0020002000200020;
defparam \state~47 .shared_arith = "off";

dffeas \state.s_dummy_wait (
	.clk(clk),
	.d(\state~47_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state~41_combout ),
	.q(\state.s_dummy_wait~q ),
	.prn(vcc));
defparam \state.s_dummy_wait .is_wysiwyg = "true";
defparam \state.s_dummy_wait .power_up = "low";

arriaii_lcell_comb \state~53 (
	.dataa(!\finished_state~q ),
	.datab(!\state.s_dummy_wait~q ),
	.datac(!\state.s_refresh_done~q ),
	.datad(!\refreshes_maxed~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~53_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~53 .extended_lut = "off";
defparam \state~53 .lut_mask = 64'h1511151115111511;
defparam \state~53 .shared_arith = "off";

arriaii_lcell_comb \state~54 (
	.dataa(!\cal_complete~combout ),
	.datab(!\state.s_refresh~q ),
	.datac(!\state~43_combout ),
	.datad(!\state~53_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~54_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~54 .extended_lut = "off";
defparam \state~54 .lut_mask = 64'h20AA20AA20AA20AA;
defparam \state~54 .shared_arith = "off";

dffeas \state.s_refresh (
	.clk(clk),
	.d(\state~54_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_refresh~q ),
	.prn(vcc));
defparam \state.s_refresh .is_wysiwyg = "true";
defparam \state.s_refresh .power_up = "low";

arriaii_lcell_comb \state~55 (
	.dataa(!\cal_complete~combout ),
	.datab(!\state.s_access~q ),
	.datac(!\finished_state~q ),
	.datad(!dgb_ac_access_req),
	.datae(!\state.s_access_precharge~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~55_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~55 .extended_lut = "off";
defparam \state~55 .lut_mask = 64'h2200A2A02200A2A0;
defparam \state~55 .shared_arith = "off";

dffeas \state.s_access_precharge (
	.clk(clk),
	.d(\state~55_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_access_precharge~q ),
	.prn(vcc));
defparam \state.s_access_precharge .is_wysiwyg = "true";
defparam \state.s_access_precharge .power_up = "low";

arriaii_lcell_comb \Selector422~1 (
	.dataa(!\state.s_access_act~q ),
	.datab(!\state.s_topup_refresh~q ),
	.datac(!\state.s_refresh~q ),
	.datad(!\state.s_access_precharge~q ),
	.datae(!\state.s_zq_cal_short~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector422~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector422~1 .extended_lut = "off";
defparam \Selector422~1 .lut_mask = 64'h8000000080000000;
defparam \Selector422~1 .shared_arith = "off";

arriaii_lcell_comb \Selector424~0 (
	.dataa(!\state.s_run_init_seq~q ),
	.datab(!\stage_counter[17]~1_combout ),
	.datac(!\ac_state.s_1~q ),
	.datad(!\ac_state.s_2~q ),
	.datae(!\Selector422~1_combout ),
	.dataf(!\WideOr34~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector424~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector424~0 .extended_lut = "off";
defparam \Selector424~0 .lut_mask = 64'h0FFF0DFF0F0F0D0D;
defparam \Selector424~0 .shared_arith = "off";

dffeas \ac_state.s_2 (
	.clk(clk),
	.d(\Selector424~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\stage_counter~0_combout ),
	.q(\ac_state.s_2~q ),
	.prn(vcc));
defparam \ac_state.s_2 .is_wysiwyg = "true";
defparam \ac_state.s_2 .power_up = "low";

arriaii_lcell_comb \WideNor1~0 (
	.dataa(!\ac_state.s_5~q ),
	.datab(!\ac_state.s_4~q ),
	.datac(!\ac_state.s_2~q ),
	.datad(!\ac_state.s_3~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor1~0 .extended_lut = "off";
defparam \WideNor1~0 .lut_mask = 64'h8000800080008000;
defparam \WideNor1~0 .shared_arith = "off";

arriaii_lcell_comb \WideNor1~1 (
	.dataa(!\ac_state.s_1~q ),
	.datab(!\ac_state.s_0~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor1~1 .extended_lut = "off";
defparam \WideNor1~1 .lut_mask = 64'h2222222222222222;
defparam \WideNor1~1 .shared_arith = "off";

arriaii_lcell_comb \Selector595~0 (
	.dataa(!\state.s_run_init_seq~q ),
	.datab(!\ac_state.s_12~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector595~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector595~0 .extended_lut = "off";
defparam \Selector595~0 .lut_mask = 64'h1111111111111111;
defparam \Selector595~0 .shared_arith = "off";

arriaii_lcell_comb \Selector422~0 (
	.dataa(!\state.s_program_cal_mrs~q ),
	.datab(!\ac_state.s_6~q ),
	.datac(!\WideNor1~0_combout ),
	.datad(!\WideNor1~1_combout ),
	.datae(!\Selector595~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector422~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector422~0 .extended_lut = "off";
defparam \Selector422~0 .lut_mask = 64'hEEEA0000EEEA0000;
defparam \Selector422~0 .shared_arith = "off";

arriaii_lcell_comb \Selector422~2 (
	.dataa(!\addr_cmd~14_combout ),
	.datab(!\ac_state.s_1~q ),
	.datac(!\ac_state.s_0~q ),
	.datad(!\Selector422~1_combout ),
	.datae(!\WideOr34~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector422~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector422~2 .extended_lut = "off";
defparam \Selector422~2 .lut_mask = 64'h0105F1F50105F1F5;
defparam \Selector422~2 .shared_arith = "off";

arriaii_lcell_comb \Selector422~3 (
	.dataa(!\state.s_prog_user_mrs~q ),
	.datab(!\ac_state.s_7~q ),
	.datac(!\WideOr16~combout ),
	.datad(!\Selector422~0_combout ),
	.datae(!\Selector422~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector422~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector422~3 .extended_lut = "off";
defparam \Selector422~3 .lut_mask = 64'h000000AE000000AE;
defparam \Selector422~3 .shared_arith = "off";

dffeas \ac_state.s_0 (
	.clk(clk),
	.d(\Selector422~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\stage_counter~0_combout ),
	.q(\ac_state.s_0~q ),
	.prn(vcc));
defparam \ac_state.s_0 .is_wysiwyg = "true";
defparam \ac_state.s_0 .power_up = "low";

arriaii_lcell_comb \Selector433~0 (
	.dataa(!\state.s_run_init_seq~q ),
	.datab(!\ac_state.s_12~q ),
	.datac(!\ac_state.s_0~q ),
	.datad(!\ac_state.s_11~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector433~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector433~0 .extended_lut = "off";
defparam \Selector433~0 .lut_mask = 64'h0400040004000400;
defparam \Selector433~0 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~14 (
	.dataa(!\state.s_dummy_wait~q ),
	.datab(!\state.s_topup_refresh_done~q ),
	.datac(!\state.s_refresh_done~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~14 .extended_lut = "off";
defparam \addr_cmd~14 .lut_mask = 64'h8080808080808080;
defparam \addr_cmd~14 .shared_arith = "off";

arriaii_lcell_comb \stage_counter[17]~2 (
	.dataa(!\state.s_program_cal_mrs~q ),
	.datab(!\ac_state.s_6~q ),
	.datac(!\WideNor1~0_combout ),
	.datad(!\WideNor1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter[17]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter[17]~2 .extended_lut = "off";
defparam \stage_counter[17]~2 .lut_mask = 64'h0004000400040004;
defparam \stage_counter[17]~2 .shared_arith = "off";

arriaii_lcell_comb \stage_counter[17]~3 (
	.dataa(!\state.s_prog_user_mrs~q ),
	.datab(!\WideOr16~combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter[17]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter[17]~3 .extended_lut = "off";
defparam \stage_counter[17]~3 .lut_mask = 64'h4444444444444444;
defparam \stage_counter[17]~3 .shared_arith = "off";

arriaii_lcell_comb \Selector448~0 (
	.dataa(!\WideNor2~combout ),
	.datab(!\Selector422~1_combout ),
	.datac(!\stage_counter[17]~2_combout ),
	.datad(!\stage_counter[17]~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector448~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector448~0 .extended_lut = "off";
defparam \Selector448~0 .lut_mask = 64'hB000B000B000B000;
defparam \Selector448~0 .shared_arith = "off";

arriaii_lcell_comb \Selector452~0 (
	.dataa(!\state.s_reset~q ),
	.datab(!\addr_cmd~14_combout ),
	.datac(!\ac_state.s_1~q ),
	.datad(!\stage_counter[2]~q ),
	.datae(!\Selector448~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector452~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector452~0 .extended_lut = "off";
defparam \Selector452~0 .lut_mask = 64'h0055004000550040;
defparam \Selector452~0 .shared_arith = "off";

arriaii_lcell_comb \Selector472~2 (
	.dataa(!\ac_state.s_2~q ),
	.datab(!\ac_state.s_3~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector472~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector472~2 .extended_lut = "off";
defparam \Selector472~2 .lut_mask = 64'h8888888888888888;
defparam \Selector472~2 .shared_arith = "off";

arriaii_lcell_comb \Selector452~1 (
	.dataa(!\state.s_program_cal_mrs~q ),
	.datab(!\state.s_prog_user_mrs~q ),
	.datac(!\ac_state.s_1~q ),
	.datad(!\ac_state.s_4~q ),
	.datae(!\Selector472~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector452~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector452~1 .extended_lut = "off";
defparam \Selector452~1 .lut_mask = 64'h8888FAC88888FAC8;
defparam \Selector452~1 .shared_arith = "off";

arriaii_lcell_comb \Selector452~2 (
	.dataa(!\state.s_run_init_seq~q ),
	.datab(!\state.s_access_act~q ),
	.datac(!\addr_cmd~14_combout ),
	.datad(!\ac_state.s_0~q ),
	.datae(!\Selector452~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector452~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector452~2 .extended_lut = "off";
defparam \Selector452~2 .lut_mask = 64'h000008FF000008FF;
defparam \Selector452~2 .shared_arith = "off";

arriaii_lcell_comb \Selector450~0 (
	.dataa(!\state.s_dummy_wait~q ),
	.datab(!\state.s_topup_refresh_done~q ),
	.datac(!\state.s_refresh_done~q ),
	.datad(!\ac_state.s_1~q ),
	.datae(!\ac_state.s_0~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector450~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector450~0 .extended_lut = "off";
defparam \Selector450~0 .lut_mask = 64'h3F007F003F007F00;
defparam \Selector450~0 .shared_arith = "off";

arriaii_lcell_comb \Selector450~1 (
	.dataa(!\state.s_reset~q ),
	.datab(!\Selector448~0_combout ),
	.datac(!\Selector450~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector450~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector450~1 .extended_lut = "off";
defparam \Selector450~1 .lut_mask = 64'h4545454545454545;
defparam \Selector450~1 .shared_arith = "off";

arriaii_lcell_comb \Selector421~0 (
	.dataa(!\state.s_program_cal_mrs~q ),
	.datab(!\ac_state.s_5~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector421~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector421~0 .extended_lut = "off";
defparam \Selector421~0 .lut_mask = 64'h1111111111111111;
defparam \Selector421~0 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~57 (
	.dataa(!\ac_state.s_1~q ),
	.datab(!\state.s_zq_cal_short~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~57_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~57 .extended_lut = "off";
defparam \addr_cmd~57 .lut_mask = 64'h1111111111111111;
defparam \addr_cmd~57 .shared_arith = "off";

arriaii_lcell_comb \Selector453~1 (
	.dataa(!\state.s_run_init_seq~q ),
	.datab(!\ac_state.s_11~q ),
	.datac(!\Selector421~0_combout ),
	.datad(!\addr_cmd~57_combout ),
	.datae(!\Selector453~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector453~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector453~1 .extended_lut = "off";
defparam \Selector453~1 .lut_mask = 64'hE0000000E0000000;
defparam \Selector453~1 .shared_arith = "off";

arriaii_lcell_comb \Add3~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\stage_counter[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~1_sumout ),
	.cout(\Add3~2 ),
	.shareout());
defparam \Add3~1 .extended_lut = "off";
defparam \Add3~1 .lut_mask = 64'h00000000000000FF;
defparam \Add3~1 .shared_arith = "off";

arriaii_lcell_comb \Selector454~0 (
	.dataa(!\state.s_reset~q ),
	.datab(!\addr_cmd~14_combout ),
	.datac(!\ac_state.s_1~q ),
	.datad(!\ac_state.s_0~q ),
	.datae(!\stage_counter[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector454~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector454~0 .extended_lut = "off";
defparam \Selector454~0 .lut_mask = 64'h0C0C0C4C0C0C0C4C;
defparam \Selector454~0 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~7 (
	.dataa(!\state.s_topup_refresh~q ),
	.datab(!\state.s_refresh~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~7 .extended_lut = "off";
defparam \addr_cmd~7 .lut_mask = 64'h8888888888888888;
defparam \addr_cmd~7 .shared_arith = "off";

arriaii_lcell_comb \Selector454~1 (
	.dataa(!\state.s_reset~q ),
	.datab(!\addr_cmd~7_combout ),
	.datac(!\stage_counter[17]~2_combout ),
	.datad(!\stage_counter[17]~3_combout ),
	.datae(!\stage_counter[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector454~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector454~1 .extended_lut = "off";
defparam \Selector454~1 .lut_mask = 64'h0000455500004555;
defparam \Selector454~1 .shared_arith = "off";

arriaii_lcell_comb WideNor2(
	.dataa(!\ac_state.s_1~q ),
	.datab(!\ac_state.s_2~q ),
	.datac(!\ac_state.s_0~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor2~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideNor2.extended_lut = "off";
defparam WideNor2.lut_mask = 64'h0808080808080808;
defparam WideNor2.shared_arith = "off";

arriaii_lcell_comb \Selector595~3 (
	.dataa(!\state.s_access_act~q ),
	.datab(!\state.s_access_precharge~q ),
	.datac(!\state.s_zq_cal_short~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector595~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector595~3 .extended_lut = "off";
defparam \Selector595~3 .lut_mask = 64'h8080808080808080;
defparam \Selector595~3 .shared_arith = "off";

arriaii_lcell_comb \Selector454~2 (
	.dataa(!\state.s_reset~q ),
	.datab(!\ac_state.s_2~q ),
	.datac(!\WideNor1~1_combout ),
	.datad(!\Selector595~3_combout ),
	.datae(!\stage_counter[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector454~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector454~2 .extended_lut = "off";
defparam \Selector454~2 .lut_mask = 64'h3300370033003700;
defparam \Selector454~2 .shared_arith = "off";

arriaii_lcell_comb \Selector454~3 (
	.dataa(!\state.s_run_init_seq~q ),
	.datab(!\state.s_prog_user_mrs~q ),
	.datac(!\ac_state.s_12~q ),
	.datad(!\ac_state.s_0~q ),
	.datae(!\ac_state.s_11~q ),
	.dataf(!\state.s_zq_cal_short~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector454~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector454~3 .extended_lut = "off";
defparam \Selector454~3 .lut_mask = 64'h88AA88FA00AA00FA;
defparam \Selector454~3 .shared_arith = "off";

arriaii_lcell_comb \Selector454~4 (
	.dataa(!\state.s_program_cal_mrs~q ),
	.datab(!\state.s_prog_user_mrs~q ),
	.datac(!\ac_state.s_6~q ),
	.datad(!\ac_state.s_7~q ),
	.datae(!\Selector454~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector454~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector454~4 .extended_lut = "off";
defparam \Selector454~4 .lut_mask = 64'h0000F8C80000F8C8;
defparam \Selector454~4 .shared_arith = "off";

arriaii_lcell_comb \Selector454~5 (
	.dataa(!\addr_cmd~7_combout ),
	.datab(!\WideNor2~combout ),
	.datac(!\WideOr34~0_combout ),
	.datad(!\Selector454~2_combout ),
	.datae(!\Selector454~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector454~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector454~5 .extended_lut = "off";
defparam \Selector454~5 .lut_mask = 64'h0000070000000700;
defparam \Selector454~5 .shared_arith = "off";

arriaii_lcell_comb \stage_counter~37 (
	.dataa(!\stage_counter~0_combout ),
	.datab(!\Add3~1_sumout ),
	.datac(!\Selector454~0_combout ),
	.datad(!\Selector454~1_combout ),
	.datae(!\Selector454~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter~37 .extended_lut = "off";
defparam \stage_counter~37 .lut_mask = 64'h7777277777772777;
defparam \stage_counter~37 .shared_arith = "off";

dffeas \stage_counter[0] (
	.clk(clk),
	.d(\stage_counter~37_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\stage_counter[0]~q ),
	.prn(vcc));
defparam \stage_counter[0] .is_wysiwyg = "true";
defparam \stage_counter[0] .power_up = "low";

arriaii_lcell_comb \Add3~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\stage_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~5_sumout ),
	.cout(\Add3~6 ),
	.shareout());
defparam \Add3~5 .extended_lut = "off";
defparam \Add3~5 .lut_mask = 64'h00000000000000FF;
defparam \Add3~5 .shared_arith = "off";

arriaii_lcell_comb \stage_counter~4 (
	.dataa(!\stage_counter~0_combout ),
	.datab(!\stage_counter[1]~q ),
	.datac(!\Selector450~1_combout ),
	.datad(!\Selector453~1_combout ),
	.datae(!\Add3~5_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter~4 .extended_lut = "off";
defparam \stage_counter~4 .lut_mask = 64'h5501FFAB5501FFAB;
defparam \stage_counter~4 .shared_arith = "off";

dffeas \stage_counter[1] (
	.clk(clk),
	.d(\stage_counter~4_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\stage_counter[1]~q ),
	.prn(vcc));
defparam \stage_counter[1] .is_wysiwyg = "true";
defparam \stage_counter[1] .power_up = "low";

arriaii_lcell_comb \Add3~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\stage_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~9_sumout ),
	.cout(\Add3~10 ),
	.shareout());
defparam \Add3~9 .extended_lut = "off";
defparam \Add3~9 .lut_mask = 64'h00000000000000FF;
defparam \Add3~9 .shared_arith = "off";

arriaii_lcell_comb \stage_counter~5 (
	.dataa(!\stage_counter~0_combout ),
	.datab(!\Selector433~0_combout ),
	.datac(!\Selector452~0_combout ),
	.datad(!\Selector452~2_combout ),
	.datae(!\Add3~9_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter~5 .extended_lut = "off";
defparam \stage_counter~5 .lut_mask = 64'h5515FFBF5515FFBF;
defparam \stage_counter~5 .shared_arith = "off";

dffeas \stage_counter[2] (
	.clk(clk),
	.d(\stage_counter~5_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\stage_counter[2]~q ),
	.prn(vcc));
defparam \stage_counter[2] .is_wysiwyg = "true";
defparam \stage_counter[2] .power_up = "low";

arriaii_lcell_comb \Selector448~1 (
	.dataa(!\state.s_reset~q ),
	.datab(!\addr_cmd~14_combout ),
	.datac(!\WideNor1~1_combout ),
	.datad(!\Selector448~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector448~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector448~1 .extended_lut = "off";
defparam \Selector448~1 .lut_mask = 64'h5504550455045504;
defparam \Selector448~1 .shared_arith = "off";

arriaii_lcell_comb \Selector451~0 (
	.dataa(!\state.s_prog_user_mrs~q ),
	.datab(!\state.s_access_act~q ),
	.datac(!\ac_state.s_1~q ),
	.datad(!\ac_state.s_5~q ),
	.datae(!\ac_state.s_0~q ),
	.dataf(!\state.s_access_precharge~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector451~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector451~0 .extended_lut = "off";
defparam \Selector451~0 .lut_mask = 64'hF8A8F8A80000F0A0;
defparam \Selector451~0 .shared_arith = "off";

arriaii_lcell_comb \Selector451~1 (
	.dataa(!\state.s_program_cal_mrs~q ),
	.datab(!\ac_state.s_4~q ),
	.datac(!\ac_state.s_0~q ),
	.datad(!\Selector433~0_combout ),
	.datae(!\Selector451~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector451~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector451~1 .extended_lut = "off";
defparam \Selector451~1 .lut_mask = 64'h0000AE000000AE00;
defparam \Selector451~1 .shared_arith = "off";

arriaii_lcell_comb \Add3~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\stage_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~13_sumout ),
	.cout(\Add3~14 ),
	.shareout());
defparam \Add3~13 .extended_lut = "off";
defparam \Add3~13 .lut_mask = 64'h00000000000000FF;
defparam \Add3~13 .shared_arith = "off";

arriaii_lcell_comb \stage_counter~6 (
	.dataa(!\stage_counter~0_combout ),
	.datab(!\stage_counter[3]~q ),
	.datac(!\Selector448~1_combout ),
	.datad(!\Selector451~1_combout ),
	.datae(!\Add3~13_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter~6 .extended_lut = "off";
defparam \stage_counter~6 .lut_mask = 64'h5501FFAB5501FFAB;
defparam \stage_counter~6 .shared_arith = "off";

dffeas \stage_counter[3] (
	.clk(clk),
	.d(\stage_counter~6_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\stage_counter[3]~q ),
	.prn(vcc));
defparam \stage_counter[3] .is_wysiwyg = "true";
defparam \stage_counter[3] .power_up = "low";

arriaii_lcell_comb \Selector449~0 (
	.dataa(!\state.s_run_init_seq~q ),
	.datab(!\state.s_topup_refresh_done~q ),
	.datac(!\state.s_refresh_done~q ),
	.datad(!\ac_state.s_0~q ),
	.datae(!\ac_state.s_11~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector449~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector449~0 .extended_lut = "off";
defparam \Selector449~0 .lut_mask = 64'h80FF80AA80FF80AA;
defparam \Selector449~0 .shared_arith = "off";

arriaii_lcell_comb \Selector449~1 (
	.dataa(!\state.s_run_init_seq~q ),
	.datab(!\state.s_topup_refresh_done~q ),
	.datac(!\state.s_refresh_done~q ),
	.datad(!\ac_state.s_0~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector449~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector449~1 .extended_lut = "off";
defparam \Selector449~1 .lut_mask = 64'h7F007F007F007F00;
defparam \Selector449~1 .shared_arith = "off";

arriaii_lcell_comb \Add3~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\stage_counter[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~17_sumout ),
	.cout(\Add3~18 ),
	.shareout());
defparam \Add3~17 .extended_lut = "off";
defparam \Add3~17 .lut_mask = 64'h00000000000000FF;
defparam \Add3~17 .shared_arith = "off";

arriaii_lcell_comb \stage_counter~8 (
	.dataa(!\stage_counter~0_combout ),
	.datab(!\stage_counter[4]~q ),
	.datac(!\Selector450~1_combout ),
	.datad(!\Selector449~1_combout ),
	.datae(!\Add3~17_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter~8 .extended_lut = "off";
defparam \stage_counter~8 .lut_mask = 64'h0155ABFF0155ABFF;
defparam \stage_counter~8 .shared_arith = "off";

dffeas \stage_counter[4] (
	.clk(clk),
	.d(\stage_counter~8_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\stage_counter[4]~q ),
	.prn(vcc));
defparam \stage_counter[4] .is_wysiwyg = "true";
defparam \stage_counter[4] .power_up = "low";

arriaii_lcell_comb \Add3~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\stage_counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~21_sumout ),
	.cout(\Add3~22 ),
	.shareout());
defparam \Add3~21 .extended_lut = "off";
defparam \Add3~21 .lut_mask = 64'h00000000000000FF;
defparam \Add3~21 .shared_arith = "off";

arriaii_lcell_comb \stage_counter~7 (
	.dataa(!\stage_counter~0_combout ),
	.datab(!\stage_counter[5]~q ),
	.datac(!\Selector450~1_combout ),
	.datad(!\Selector449~0_combout ),
	.datae(!\Add3~21_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter~7 .extended_lut = "off";
defparam \stage_counter~7 .lut_mask = 64'h5501FFAB5501FFAB;
defparam \stage_counter~7 .shared_arith = "off";

dffeas \stage_counter[5] (
	.clk(clk),
	.d(\stage_counter~7_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\stage_counter[5]~q ),
	.prn(vcc));
defparam \stage_counter[5] .is_wysiwyg = "true";
defparam \stage_counter[5] .power_up = "low";

arriaii_lcell_comb \stage_counter_zero~0 (
	.dataa(!\stage_counter[1]~q ),
	.datab(!\stage_counter[2]~q ),
	.datac(!\stage_counter[3]~q ),
	.datad(!\stage_counter[5]~q ),
	.datae(!\stage_counter[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter_zero~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter_zero~0 .extended_lut = "off";
defparam \stage_counter_zero~0 .lut_mask = 64'h8000000080000000;
defparam \stage_counter_zero~0 .shared_arith = "off";

arriaii_lcell_comb \stage_counter[17]~9 (
	.dataa(!\stage_counter[17]~1_combout ),
	.datab(!\WideNor2~combout ),
	.datac(!\Selector422~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter[17]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter[17]~9 .extended_lut = "off";
defparam \stage_counter[17]~9 .lut_mask = 64'h1010101010101010;
defparam \stage_counter[17]~9 .shared_arith = "off";

arriaii_lcell_comb \stage_counter[17]~10 (
	.dataa(!\stage_counter[17]~1_combout ),
	.datab(!\addr_cmd~14_combout ),
	.datac(!\WideNor1~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter[17]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter[17]~10 .extended_lut = "off";
defparam \stage_counter[17]~10 .lut_mask = 64'h0404040404040404;
defparam \stage_counter[17]~10 .shared_arith = "off";

arriaii_lcell_comb \stage_counter[17]~11 (
	.dataa(!\state.s_program_cal_mrs~q ),
	.datab(!\state.s_prog_user_mrs~q ),
	.datac(!\WideOr16~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter[17]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter[17]~11 .extended_lut = "off";
defparam \stage_counter[17]~11 .lut_mask = 64'h2020202020202020;
defparam \stage_counter[17]~11 .shared_arith = "off";

arriaii_lcell_comb \stage_counter[17]~12 (
	.dataa(!\state.s_access~q ),
	.datab(!\state.s_run_init_seq~q ),
	.datac(!\state.s_reset~q ),
	.datad(!\state.s_idle~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter[17]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter[17]~12 .extended_lut = "off";
defparam \stage_counter[17]~12 .lut_mask = 64'h0800080008000800;
defparam \stage_counter[17]~12 .shared_arith = "off";

arriaii_lcell_comb \stage_counter[17]~18 (
	.dataa(!\stage_counter[17]~2_combout ),
	.datab(!\stage_counter[17]~9_combout ),
	.datac(!\stage_counter[17]~10_combout ),
	.datad(!\stage_counter[17]~11_combout ),
	.datae(!\stage_counter[17]~12_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter[17]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter[17]~18 .extended_lut = "off";
defparam \stage_counter[17]~18 .lut_mask = 64'h00007FFF00007FFF;
defparam \stage_counter[17]~18 .shared_arith = "off";

arriaii_lcell_comb \Add3~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\stage_counter[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~25_sumout ),
	.cout(\Add3~26 ),
	.shareout());
defparam \Add3~25 .extended_lut = "off";
defparam \Add3~25 .lut_mask = 64'h00000000000000FF;
defparam \Add3~25 .shared_arith = "off";

arriaii_lcell_comb \stage_counter~27 (
	.dataa(!\stage_counter~0_combout ),
	.datab(!\addr_cmd~57_combout ),
	.datac(!\stage_counter[6]~q ),
	.datad(!\Selector433~0_combout ),
	.datae(!\Selector448~1_combout ),
	.dataf(!\Add3~25_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter~27 .extended_lut = "off";
defparam \stage_counter~27 .lut_mask = 64'h11551555BBFFBFFF;
defparam \stage_counter~27 .shared_arith = "off";

dffeas \stage_counter[6] (
	.clk(clk),
	.d(\stage_counter~27_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\stage_counter[6]~q ),
	.prn(vcc));
defparam \stage_counter[6] .is_wysiwyg = "true";
defparam \stage_counter[6] .power_up = "low";

arriaii_lcell_comb \Add3~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\stage_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~29_sumout ),
	.cout(\Add3~30 ),
	.shareout());
defparam \Add3~29 .extended_lut = "off";
defparam \Add3~29 .lut_mask = 64'h00000000000000FF;
defparam \Add3~29 .shared_arith = "off";

arriaii_lcell_comb \stage_counter[8]~14 (
	.dataa(!\state.s_run_init_seq~q ),
	.datab(!\state.s_reset~q ),
	.datac(!\stage_counter_zero~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter[8]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter[8]~14 .extended_lut = "off";
defparam \stage_counter[8]~14 .lut_mask = 64'h1313131313131313;
defparam \stage_counter[8]~14 .shared_arith = "off";

arriaii_lcell_comb \stage_counter~28 (
	.dataa(!\state.s_reset~q ),
	.datab(!\stage_counter[7]~q ),
	.datac(!\Add3~29_sumout ),
	.datad(!\stage_counter[8]~14_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter~28 .extended_lut = "off";
defparam \stage_counter~28 .lut_mask = 64'h110F110F110F110F;
defparam \stage_counter~28 .shared_arith = "off";

arriaii_lcell_comb \stage_counter~29 (
	.dataa(!\state.s_run_init_seq~q ),
	.datab(!\state.s_reset~q ),
	.datac(!\stage_counter_zero~q ),
	.datad(!\ac_state.s_11~q ),
	.datae(!\stage_counter[17]~18_combout ),
	.dataf(!\stage_counter~28_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter~29 .extended_lut = "off";
defparam \stage_counter~29 .lut_mask = 64'h001000100313FFFF;
defparam \stage_counter~29 .shared_arith = "off";

dffeas \stage_counter[7] (
	.clk(clk),
	.d(\stage_counter~29_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\stage_counter[7]~q ),
	.prn(vcc));
defparam \stage_counter[7] .is_wysiwyg = "true";
defparam \stage_counter[7] .power_up = "low";

arriaii_lcell_comb \Add3~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\stage_counter[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~33_sumout ),
	.cout(\Add3~34 ),
	.shareout());
defparam \Add3~33 .extended_lut = "off";
defparam \Add3~33 .lut_mask = 64'h00000000000000FF;
defparam \Add3~33 .shared_arith = "off";

arriaii_lcell_comb \stage_counter[8]~13 (
	.dataa(!\stage_counter~0_combout ),
	.datab(!\stage_counter[17]~2_combout ),
	.datac(!\stage_counter[17]~9_combout ),
	.datad(!\stage_counter[17]~10_combout ),
	.datae(!\stage_counter[17]~11_combout ),
	.dataf(!\stage_counter[17]~12_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter[8]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter[8]~13 .extended_lut = "off";
defparam \stage_counter[8]~13 .lut_mask = 64'h5555555540000000;
defparam \stage_counter[8]~13 .shared_arith = "off";

arriaii_lcell_comb \stage_counter~15 (
	.dataa(!\ac_state.s_12~q ),
	.datab(!\ac_state.s_0~q ),
	.datac(!\ac_state.s_11~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter~15 .extended_lut = "off";
defparam \stage_counter~15 .lut_mask = 64'h1313131313131313;
defparam \stage_counter~15 .shared_arith = "off";

arriaii_lcell_comb \stage_counter~30 (
	.dataa(!\state.s_reset~q ),
	.datab(!\stage_counter[8]~q ),
	.datac(!\stage_counter[8]~13_combout ),
	.datad(!\stage_counter[8]~14_combout ),
	.datae(!\stage_counter~15_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter~30 .extended_lut = "off";
defparam \stage_counter~30 .lut_mask = 64'h100F1000100F1000;
defparam \stage_counter~30 .shared_arith = "off";

arriaii_lcell_comb \stage_counter~31 (
	.dataa(!\stage_counter~0_combout ),
	.datab(!\Add3~33_sumout ),
	.datac(!\stage_counter~30_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter~31 .extended_lut = "off";
defparam \stage_counter~31 .lut_mask = 64'h2F2F2F2F2F2F2F2F;
defparam \stage_counter~31 .shared_arith = "off";

dffeas \stage_counter[8] (
	.clk(clk),
	.d(\stage_counter~31_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\stage_counter[8]~q ),
	.prn(vcc));
defparam \stage_counter[8] .is_wysiwyg = "true";
defparam \stage_counter[8] .power_up = "low";

arriaii_lcell_comb \Add3~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\stage_counter[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~37_sumout ),
	.cout(\Add3~38 ),
	.shareout());
defparam \Add3~37 .extended_lut = "off";
defparam \Add3~37 .lut_mask = 64'h00000000000000FF;
defparam \Add3~37 .shared_arith = "off";

arriaii_lcell_comb \stage_counter~32 (
	.dataa(!\stage_counter~0_combout ),
	.datab(!\Selector421~0_combout ),
	.datac(!\stage_counter[9]~q ),
	.datad(!\Selector448~1_combout ),
	.datae(!\Add3~37_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter~32 .extended_lut = "off";
defparam \stage_counter~32 .lut_mask = 64'h1115BBBF1115BBBF;
defparam \stage_counter~32 .shared_arith = "off";

dffeas \stage_counter[9] (
	.clk(clk),
	.d(\stage_counter~32_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\stage_counter[9]~q ),
	.prn(vcc));
defparam \stage_counter[9] .is_wysiwyg = "true";
defparam \stage_counter[9] .power_up = "low";

arriaii_lcell_comb \Add3~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\stage_counter[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~41_sumout ),
	.cout(\Add3~42 ),
	.shareout());
defparam \Add3~41 .extended_lut = "off";
defparam \Add3~41 .lut_mask = 64'h00000000000000FF;
defparam \Add3~41 .shared_arith = "off";

arriaii_lcell_comb \stage_counter~35 (
	.dataa(!\state.s_reset~q ),
	.datab(!\stage_counter[10]~q ),
	.datac(!\stage_counter[8]~13_combout ),
	.datad(!\stage_counter[8]~14_combout ),
	.datae(!\stage_counter~15_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter~35 .extended_lut = "off";
defparam \stage_counter~35 .lut_mask = 64'h100F1000100F1000;
defparam \stage_counter~35 .shared_arith = "off";

arriaii_lcell_comb \stage_counter~36 (
	.dataa(!\stage_counter~0_combout ),
	.datab(!\Add3~41_sumout ),
	.datac(!\stage_counter~35_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter~36 .extended_lut = "off";
defparam \stage_counter~36 .lut_mask = 64'h2F2F2F2F2F2F2F2F;
defparam \stage_counter~36 .shared_arith = "off";

dffeas \stage_counter[10] (
	.clk(clk),
	.d(\stage_counter~36_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\stage_counter[10]~q ),
	.prn(vcc));
defparam \stage_counter[10] .is_wysiwyg = "true";
defparam \stage_counter[10] .power_up = "low";

arriaii_lcell_comb \Add3~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\stage_counter[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~45_sumout ),
	.cout(\Add3~46 ),
	.shareout());
defparam \Add3~45 .extended_lut = "off";
defparam \Add3~45 .lut_mask = 64'h00000000000000FF;
defparam \Add3~45 .shared_arith = "off";

arriaii_lcell_comb \stage_counter~33 (
	.dataa(!\state.s_reset~q ),
	.datab(!\process_12~0_combout ),
	.datac(!\stage_counter[11]~q ),
	.datad(!\stage_counter[8]~13_combout ),
	.datae(!\stage_counter[8]~14_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter~33 .extended_lut = "off";
defparam \stage_counter~33 .lut_mask = 64'h0500003305000033;
defparam \stage_counter~33 .shared_arith = "off";

arriaii_lcell_comb \stage_counter~34 (
	.dataa(!\stage_counter~0_combout ),
	.datab(!\Add3~45_sumout ),
	.datac(!\stage_counter~33_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter~34 .extended_lut = "off";
defparam \stage_counter~34 .lut_mask = 64'h2F2F2F2F2F2F2F2F;
defparam \stage_counter~34 .shared_arith = "off";

dffeas \stage_counter[11] (
	.clk(clk),
	.d(\stage_counter~34_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\stage_counter[11]~q ),
	.prn(vcc));
defparam \stage_counter[11] .is_wysiwyg = "true";
defparam \stage_counter[11] .power_up = "low";

arriaii_lcell_comb \Add3~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\stage_counter[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~49_sumout ),
	.cout(\Add3~50 ),
	.shareout());
defparam \Add3~49 .extended_lut = "off";
defparam \Add3~49 .lut_mask = 64'h00000000000000FF;
defparam \Add3~49 .shared_arith = "off";

arriaii_lcell_comb \stage_counter~16 (
	.dataa(!\state.s_reset~q ),
	.datab(!\stage_counter[12]~q ),
	.datac(!\stage_counter[8]~13_combout ),
	.datad(!\stage_counter[8]~14_combout ),
	.datae(!\stage_counter~15_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter~16 .extended_lut = "off";
defparam \stage_counter~16 .lut_mask = 64'h100F1000100F1000;
defparam \stage_counter~16 .shared_arith = "off";

arriaii_lcell_comb \stage_counter~17 (
	.dataa(!\stage_counter~0_combout ),
	.datab(!\Add3~49_sumout ),
	.datac(!\stage_counter~16_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter~17 .extended_lut = "off";
defparam \stage_counter~17 .lut_mask = 64'h2F2F2F2F2F2F2F2F;
defparam \stage_counter~17 .shared_arith = "off";

dffeas \stage_counter[12] (
	.clk(clk),
	.d(\stage_counter~17_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\stage_counter[12]~q ),
	.prn(vcc));
defparam \stage_counter[12] .is_wysiwyg = "true";
defparam \stage_counter[12] .power_up = "low";

arriaii_lcell_comb \stage_counter~19 (
	.dataa(!\state.s_run_init_seq~q ),
	.datab(!\state.s_reset~q ),
	.datac(!\stage_counter_zero~q ),
	.datad(!\stage_counter[17]~18_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter~19 .extended_lut = "off";
defparam \stage_counter~19 .lut_mask = 64'h0020002000200020;
defparam \stage_counter~19 .shared_arith = "off";

arriaii_lcell_comb \stage_counter~20 (
	.dataa(!\state.s_run_init_seq~q ),
	.datab(!\state.s_reset~q ),
	.datac(!\stage_counter_zero~q ),
	.datad(!\ac_state.s_0~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter~20 .extended_lut = "off";
defparam \stage_counter~20 .lut_mask = 64'h1000100010001000;
defparam \stage_counter~20 .shared_arith = "off";

arriaii_lcell_comb \Add3~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\stage_counter[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~53_sumout ),
	.cout(\Add3~54 ),
	.shareout());
defparam \Add3~53 .extended_lut = "off";
defparam \Add3~53 .lut_mask = 64'h00000000000000FF;
defparam \Add3~53 .shared_arith = "off";

arriaii_lcell_comb \stage_counter~21 (
	.dataa(!\stage_counter~0_combout ),
	.datab(!\stage_counter[13]~q ),
	.datac(!\stage_counter~19_combout ),
	.datad(!\stage_counter~20_combout ),
	.datae(!\Add3~53_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter~21 .extended_lut = "off";
defparam \stage_counter~21 .lut_mask = 64'h03FFABFF03FFABFF;
defparam \stage_counter~21 .shared_arith = "off";

dffeas \stage_counter[13] (
	.clk(clk),
	.d(\stage_counter~21_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\stage_counter[13]~q ),
	.prn(vcc));
defparam \stage_counter[13] .is_wysiwyg = "true";
defparam \stage_counter[13] .power_up = "low";

arriaii_lcell_comb \Add3~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\stage_counter[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~57_sumout ),
	.cout(\Add3~58 ),
	.shareout());
defparam \Add3~57 .extended_lut = "off";
defparam \Add3~57 .lut_mask = 64'h00000000000000FF;
defparam \Add3~57 .shared_arith = "off";

arriaii_lcell_comb \stage_counter~22 (
	.dataa(!\stage_counter~0_combout ),
	.datab(!\stage_counter[14]~q ),
	.datac(!\stage_counter~19_combout ),
	.datad(!\stage_counter~20_combout ),
	.datae(!\Add3~57_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter~22 .extended_lut = "off";
defparam \stage_counter~22 .lut_mask = 64'h03FFABFF03FFABFF;
defparam \stage_counter~22 .shared_arith = "off";

dffeas \stage_counter[14] (
	.clk(clk),
	.d(\stage_counter~22_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\stage_counter[14]~q ),
	.prn(vcc));
defparam \stage_counter[14] .is_wysiwyg = "true";
defparam \stage_counter[14] .power_up = "low";

arriaii_lcell_comb \Add3~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\stage_counter[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~61_sumout ),
	.cout(\Add3~62 ),
	.shareout());
defparam \Add3~61 .extended_lut = "off";
defparam \Add3~61 .lut_mask = 64'h00000000000000FF;
defparam \Add3~61 .shared_arith = "off";

arriaii_lcell_comb \stage_counter~23 (
	.dataa(!\stage_counter~0_combout ),
	.datab(!\Add3~61_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter~23 .extended_lut = "off";
defparam \stage_counter~23 .lut_mask = 64'h2222222222222222;
defparam \stage_counter~23 .shared_arith = "off";

arriaii_lcell_comb \stage_counter[17]~24 (
	.dataa(!\stage_counter~0_combout ),
	.datab(!\stage_counter[17]~2_combout ),
	.datac(!\stage_counter[17]~9_combout ),
	.datad(!\stage_counter[17]~10_combout ),
	.datae(!\stage_counter[17]~11_combout ),
	.dataf(!\stage_counter[17]~12_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter[17]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter[17]~24 .extended_lut = "off";
defparam \stage_counter[17]~24 .lut_mask = 64'hFFFFFFFFEAAAAAAA;
defparam \stage_counter[17]~24 .shared_arith = "off";

dffeas \stage_counter[15] (
	.clk(clk),
	.d(\stage_counter~23_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\stage_counter[17]~24_combout ),
	.q(\stage_counter[15]~q ),
	.prn(vcc));
defparam \stage_counter[15] .is_wysiwyg = "true";
defparam \stage_counter[15] .power_up = "low";

arriaii_lcell_comb \Add3~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\stage_counter[16]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~65_sumout ),
	.cout(\Add3~66 ),
	.shareout());
defparam \Add3~65 .extended_lut = "off";
defparam \Add3~65 .lut_mask = 64'h00000000000000FF;
defparam \Add3~65 .shared_arith = "off";

arriaii_lcell_comb \stage_counter~26 (
	.dataa(!\stage_counter~0_combout ),
	.datab(!\Add3~65_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter~26 .extended_lut = "off";
defparam \stage_counter~26 .lut_mask = 64'h2222222222222222;
defparam \stage_counter~26 .shared_arith = "off";

dffeas \stage_counter[16] (
	.clk(clk),
	.d(\stage_counter~26_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\stage_counter[17]~24_combout ),
	.q(\stage_counter[16]~q ),
	.prn(vcc));
defparam \stage_counter[16] .is_wysiwyg = "true";
defparam \stage_counter[16] .power_up = "low";

arriaii_lcell_comb \Add3~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\stage_counter[17]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~69_sumout ),
	.cout(),
	.shareout());
defparam \Add3~69 .extended_lut = "off";
defparam \Add3~69 .lut_mask = 64'h00000000000000FF;
defparam \Add3~69 .shared_arith = "off";

arriaii_lcell_comb \stage_counter~25 (
	.dataa(!\stage_counter~0_combout ),
	.datab(!\Add3~69_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter~25 .extended_lut = "off";
defparam \stage_counter~25 .lut_mask = 64'h2222222222222222;
defparam \stage_counter~25 .shared_arith = "off";

dffeas \stage_counter[17] (
	.clk(clk),
	.d(\stage_counter~25_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\stage_counter[17]~24_combout ),
	.q(\stage_counter[17]~q ),
	.prn(vcc));
defparam \stage_counter[17] .is_wysiwyg = "true";
defparam \stage_counter[17] .power_up = "low";

arriaii_lcell_comb \stage_counter_zero~1 (
	.dataa(!\stage_counter[13]~q ),
	.datab(!\stage_counter[14]~q ),
	.datac(!\stage_counter[15]~q ),
	.datad(!\stage_counter[17]~q ),
	.datae(!\stage_counter[16]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter_zero~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter_zero~1 .extended_lut = "off";
defparam \stage_counter_zero~1 .lut_mask = 64'h8000000080000000;
defparam \stage_counter_zero~1 .shared_arith = "off";

arriaii_lcell_comb \stage_counter_zero~2 (
	.dataa(!\stage_counter[7]~q ),
	.datab(!\stage_counter[8]~q ),
	.datac(!\stage_counter[9]~q ),
	.datad(!\stage_counter[11]~q ),
	.datae(!\stage_counter[10]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter_zero~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter_zero~2 .extended_lut = "off";
defparam \stage_counter_zero~2 .lut_mask = 64'h8000000080000000;
defparam \stage_counter_zero~2 .shared_arith = "off";

arriaii_lcell_comb \stage_counter_zero~3 (
	.dataa(!\stage_counter~0_combout ),
	.datab(!\stage_counter_zero~0_combout ),
	.datac(!\stage_counter[12]~q ),
	.datad(!\stage_counter_zero~1_combout ),
	.datae(!\stage_counter[6]~q ),
	.dataf(!\stage_counter_zero~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter_zero~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter_zero~3 .extended_lut = "off";
defparam \stage_counter_zero~3 .lut_mask = 64'hFFFFFFFFFFDFFFFF;
defparam \stage_counter_zero~3 .shared_arith = "off";

dffeas stage_counter_zero(
	.clk(clk),
	.d(\stage_counter_zero~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\stage_counter_zero~q ),
	.prn(vcc));
defparam stage_counter_zero.is_wysiwyg = "true";
defparam stage_counter_zero.power_up = "low";

arriaii_lcell_comb \stage_counter~0 (
	.dataa(!\state.s_reset~q ),
	.datab(!\stage_counter_zero~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stage_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stage_counter~0 .extended_lut = "off";
defparam \stage_counter~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \stage_counter~0 .shared_arith = "off";

arriaii_lcell_comb \Selector595~1 (
	.dataa(!\state.s_program_cal_mrs~q ),
	.datab(!\state.s_prog_user_mrs~q ),
	.datac(!\ac_state.s_6~q ),
	.datad(!\ac_state.s_7~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector595~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector595~1 .extended_lut = "off";
defparam \Selector595~1 .lut_mask = 64'h0537053705370537;
defparam \Selector595~1 .shared_arith = "off";

arriaii_lcell_comb \Selector595~2 (
	.dataa(!\ac_state.s_2~q ),
	.datab(!\Selector595~0_combout ),
	.datac(!\Selector422~1_combout ),
	.datad(!\Selector595~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector595~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector595~2 .extended_lut = "off";
defparam \Selector595~2 .lut_mask = 64'h8C008C008C008C00;
defparam \Selector595~2 .shared_arith = "off";

arriaii_lcell_comb \finished_state~0 (
	.dataa(!\addr_cmd~14_combout ),
	.datab(!\stage_counter~0_combout ),
	.datac(!\ac_state.s_1~q ),
	.datad(!\Selector595~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\finished_state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \finished_state~0 .extended_lut = "off";
defparam \finished_state~0 .lut_mask = 64'h3302330233023302;
defparam \finished_state~0 .shared_arith = "off";

dffeas finished_state(
	.clk(clk),
	.d(\finished_state~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\finished_state~q ),
	.prn(vcc));
defparam finished_state.is_wysiwyg = "true";
defparam finished_state.power_up = "low";

arriaii_lcell_comb \state~49 (
	.dataa(!\cal_complete~combout ),
	.datab(!\finished_state~q ),
	.datac(!\Selector3~0_combout ),
	.datad(!\state.s_refresh_done~q ),
	.datae(!\state.s_refresh~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~49 .extended_lut = "off";
defparam \state~49 .lut_mask = 64'h008A22AA008A22AA;
defparam \state~49 .shared_arith = "off";

dffeas \state.s_refresh_done (
	.clk(clk),
	.d(\state~49_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_refresh_done~q ),
	.prn(vcc));
defparam \state.s_refresh_done .is_wysiwyg = "true";
defparam \state.s_refresh_done .power_up = "low";

arriaii_lcell_comb \Selector453~0 (
	.dataa(!\state.s_topup_refresh_done~q ),
	.datab(!\state.s_refresh_done~q ),
	.datac(!\ac_state.s_0~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector453~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector453~0 .extended_lut = "off";
defparam \Selector453~0 .lut_mask = 64'h7070707070707070;
defparam \Selector453~0 .shared_arith = "off";

arriaii_lcell_comb \refresh_done~0 (
	.dataa(!\stage_counter~0_combout ),
	.datab(!\Selector453~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\refresh_done~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \refresh_done~0 .extended_lut = "off";
defparam \refresh_done~0 .lut_mask = 64'h1111111111111111;
defparam \refresh_done~0 .shared_arith = "off";

dffeas refresh_done(
	.clk(clk),
	.d(\refresh_done~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_done~q ),
	.prn(vcc));
defparam refresh_done.is_wysiwyg = "true";
defparam refresh_done.power_up = "low";

arriaii_lcell_comb \initial_refresh_issued~0 (
	.dataa(!\cal_complete~combout ),
	.datab(!\state.s_topup_refresh_done~q ),
	.datac(!\state.s_refresh_done~q ),
	.datad(!\initial_refresh_issued~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\initial_refresh_issued~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \initial_refresh_issued~0 .extended_lut = "off";
defparam \initial_refresh_issued~0 .lut_mask = 64'h2AAA2AAA2AAA2AAA;
defparam \initial_refresh_issued~0 .shared_arith = "off";

dffeas initial_refresh_issued(
	.clk(clk),
	.d(\initial_refresh_issued~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\initial_refresh_issued~q ),
	.prn(vcc));
defparam initial_refresh_issued.is_wysiwyg = "true";
defparam initial_refresh_issued.power_up = "low";

arriaii_lcell_comb \refresh_count[6]~0 (
	.dataa(!ctl_init_fail),
	.datab(!ctl_init_success),
	.datac(!\refreshes_maxed~q ),
	.datad(!\refresh_done~q ),
	.datae(!\initial_refresh_issued~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\refresh_count[6]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \refresh_count[6]~0 .extended_lut = "off";
defparam \refresh_count[6]~0 .lut_mask = 64'h0000888000008880;
defparam \refresh_count[6]~0 .shared_arith = "off";

arriaii_lcell_comb \refresh_count[6]~1 (
	.dataa(!\refresh_count[4]~q ),
	.datab(!\refresh_count[5]~q ),
	.datac(!\Equal0~0_combout ),
	.datad(!\Equal0~1_combout ),
	.datae(!\refresh_count[6]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\refresh_count[6]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \refresh_count[6]~1 .extended_lut = "off";
defparam \refresh_count[6]~1 .lut_mask = 64'h0000FFF70000FFF7;
defparam \refresh_count[6]~1 .shared_arith = "off";

arriaii_lcell_comb \refresh_count~2 (
	.dataa(!\Add0~17_sumout ),
	.datab(!\refresh_count[6]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\refresh_count~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \refresh_count~2 .extended_lut = "off";
defparam \refresh_count~2 .lut_mask = 64'h1111111111111111;
defparam \refresh_count~2 .shared_arith = "off";

dffeas \refresh_count[4] (
	.clk(clk),
	.d(\refresh_count~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_count[4]~q ),
	.prn(vcc));
defparam \refresh_count[4] .is_wysiwyg = "true";
defparam \refresh_count[4] .power_up = "low";

arriaii_lcell_comb \process_7~0 (
	.dataa(!\cal_complete~combout ),
	.datab(!\refresh_count[4]~q ),
	.datac(!\refresh_count[5]~q ),
	.datad(!\Equal0~0_combout ),
	.datae(!\Equal0~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\process_7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \process_7~0 .extended_lut = "off";
defparam \process_7~0 .lut_mask = 64'h0000008000000080;
defparam \process_7~0 .shared_arith = "off";

dffeas refresh_due(
	.clk(clk),
	.d(\process_7~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refresh_due~q ),
	.prn(vcc));
defparam refresh_due.is_wysiwyg = "true";
defparam refresh_due.power_up = "low";

arriaii_lcell_comb \num_stacked_refreshes~2 (
	.dataa(!\cal_complete~combout ),
	.datab(!\num_stacked_refreshes[2]~q ),
	.datac(!\num_stacked_refreshes[1]~q ),
	.datad(!\num_stacked_refreshes[0]~q ),
	.datae(!\refresh_due~q ),
	.dataf(!\refresh_done~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\num_stacked_refreshes~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \num_stacked_refreshes~2 .extended_lut = "off";
defparam \num_stacked_refreshes~2 .lut_mask = 64'h00AA2A00AA02AA00;
defparam \num_stacked_refreshes~2 .shared_arith = "off";

dffeas \num_stacked_refreshes[0] (
	.clk(clk),
	.d(\num_stacked_refreshes~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\num_stacked_refreshes[0]~q ),
	.prn(vcc));
defparam \num_stacked_refreshes[0] .is_wysiwyg = "true";
defparam \num_stacked_refreshes[0] .power_up = "low";

arriaii_lcell_comb \num_stacked_refreshes~0 (
	.dataa(!\cal_complete~combout ),
	.datab(!\num_stacked_refreshes[2]~q ),
	.datac(!\num_stacked_refreshes[1]~q ),
	.datad(!\num_stacked_refreshes[0]~q ),
	.datae(!\refresh_due~q ),
	.dataf(!\refresh_done~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\num_stacked_refreshes~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \num_stacked_refreshes~0 .extended_lut = "off";
defparam \num_stacked_refreshes~0 .lut_mask = 64'h22220222222A0222;
defparam \num_stacked_refreshes~0 .shared_arith = "off";

dffeas \num_stacked_refreshes[2] (
	.clk(clk),
	.d(\num_stacked_refreshes~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\num_stacked_refreshes[2]~q ),
	.prn(vcc));
defparam \num_stacked_refreshes[2] .is_wysiwyg = "true";
defparam \num_stacked_refreshes[2] .power_up = "low";

arriaii_lcell_comb \num_stacked_refreshes~1 (
	.dataa(!\cal_complete~combout ),
	.datab(!\num_stacked_refreshes[2]~q ),
	.datac(!\num_stacked_refreshes[1]~q ),
	.datad(!\num_stacked_refreshes[0]~q ),
	.datae(!\refresh_due~q ),
	.dataf(!\refresh_done~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\num_stacked_refreshes~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \num_stacked_refreshes~1 .extended_lut = "off";
defparam \num_stacked_refreshes~1 .lut_mask = 64'h0A0A200A0AA2200A;
defparam \num_stacked_refreshes~1 .shared_arith = "off";

dffeas \num_stacked_refreshes[1] (
	.clk(clk),
	.d(\num_stacked_refreshes~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\num_stacked_refreshes[1]~q ),
	.prn(vcc));
defparam \num_stacked_refreshes[1] .is_wysiwyg = "true";
defparam \num_stacked_refreshes[1] .power_up = "low";

arriaii_lcell_comb \LessThan0~0 (
	.dataa(!\num_stacked_refreshes[2]~q ),
	.datab(!\num_stacked_refreshes[1]~q ),
	.datac(!\num_stacked_refreshes[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h0101010101010101;
defparam \LessThan0~0 .shared_arith = "off";

dffeas refreshes_maxed(
	.clk(clk),
	.d(\LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\refreshes_maxed~q ),
	.prn(vcc));
defparam refreshes_maxed.is_wysiwyg = "true";
defparam refreshes_maxed.power_up = "low";

arriaii_lcell_comb \state~35 (
	.dataa(!\admin_req_extended~q ),
	.datab(!\refreshes_maxed~q ),
	.datac(!\mem_init_complete~q ),
	.datad(!curr_cmdcmd_prep_customer_mr_setup),
	.datae(!curr_cmdcmd_init_dram),
	.dataf(!curr_cmdcmd_prog_cal_mr),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~35 .extended_lut = "off";
defparam \state~35 .lut_mask = 64'hF3A2A2A2A2A2A2A2;
defparam \state~35 .shared_arith = "off";

arriaii_lcell_comb \state~57 (
	.dataa(!\finished_state~q ),
	.datab(!\state.s_program_cal_mrs~q ),
	.datac(!\state.s_refresh_done~q ),
	.datad(!\refreshes_maxed~q ),
	.datae(!\mem_init_complete~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~57_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~57 .extended_lut = "off";
defparam \state~57 .lut_mask = 64'h1115001511150015;
defparam \state~57 .shared_arith = "off";

arriaii_lcell_comb \state~58 (
	.dataa(!\finished_state~q ),
	.datab(!\state.s_run_init_seq~q ),
	.datac(!\state.s_prog_user_mrs~q ),
	.datad(!\state.s_access_precharge~q ),
	.datae(!\state.s_idle~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~58_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~58 .extended_lut = "off";
defparam \state~58 .lut_mask = 64'hEAAAC000EAAAC000;
defparam \state~58 .shared_arith = "off";

arriaii_lcell_comb \state~59 (
	.dataa(!\cal_complete~combout ),
	.datab(!\Selector3~0_combout ),
	.datac(!\state.s_idle~q ),
	.datad(!\state~57_combout ),
	.datae(!\state~58_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~59_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~59 .extended_lut = "off";
defparam \state~59 .lut_mask = 64'h0000A8000000A800;
defparam \state~59 .shared_arith = "off";

arriaii_lcell_comb \state~60 (
	.dataa(!dgb_ac_access_req),
	.datab(!\state.s_idle~q ),
	.datac(!\state~35_combout ),
	.datad(!\state~56_combout ),
	.datae(!\state~59_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~60_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~60 .extended_lut = "off";
defparam \state~60 .lut_mask = 64'hFFFF02AAFFFF02AA;
defparam \state~60 .shared_arith = "off";

dffeas \state.s_idle (
	.clk(clk),
	.d(\state~60_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_idle~q ),
	.prn(vcc));
defparam \state.s_idle .is_wysiwyg = "true";
defparam \state.s_idle .power_up = "low";

arriaii_lcell_comb \state~62 (
	.dataa(!\state.s_access~q ),
	.datab(!\state.s_idle~q ),
	.datac(!\finished_state~q ),
	.datad(!\state~36_combout ),
	.datae(!\state.s_reset~q ),
	.dataf(!curr_cmdcmd_init_dram),
	.datag(!\admin_req_extended~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~62_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~62 .extended_lut = "on";
defparam \state~62 .lut_mask = 64'h00FF08FF0FFF08FF;
defparam \state~62 .shared_arith = "off";

arriaii_lcell_comb \state~37 (
	.dataa(!curr_cmdcmd_init_dram),
	.datab(!dgb_ac_access_req),
	.datac(!\admin_req_extended~q ),
	.datad(!\state.s_reset~q ),
	.datae(!\state.s_idle~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~37 .extended_lut = "off";
defparam \state~37 .lut_mask = 64'h0500040405000404;
defparam \state~37 .shared_arith = "off";

arriaii_lcell_comb \state~39 (
	.dataa(!\state.s_run_init_seq~q ),
	.datab(!\state~62_combout ),
	.datac(!\state~37_combout ),
	.datad(!\state~38_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~39 .extended_lut = "off";
defparam \state~39 .lut_mask = 64'h0047004700470047;
defparam \state~39 .shared_arith = "off";

dffeas \state.s_run_init_seq (
	.clk(clk),
	.d(\state~39_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_run_init_seq~q ),
	.prn(vcc));
defparam \state.s_run_init_seq .is_wysiwyg = "true";
defparam \state.s_run_init_seq .power_up = "low";

arriaii_lcell_comb \command_done~0 (
	.dataa(!\finished_state~q ),
	.datab(!\state.s_run_init_seq~q ),
	.datac(!\state.s_program_cal_mrs~q ),
	.datad(!\state.s_prog_user_mrs~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\command_done~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \command_done~0 .extended_lut = "off";
defparam \command_done~0 .lut_mask = 64'h1555155515551555;
defparam \command_done~0 .shared_arith = "off";

dffeas command_done(
	.clk(clk),
	.d(\command_done~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\command_done~q ),
	.prn(vcc));
defparam command_done.is_wysiwyg = "true";
defparam command_done.power_up = "low";

arriaii_lcell_comb \addr_cmd~0 (
	.dataa(!\state.s_reset~q ),
	.datab(!\state.s_dummy_wait~q ),
	.datac(!\state.s_topup_refresh_done~q ),
	.datad(!\state.s_refresh_done~q ),
	.datae(!\stage_counter_zero~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~0 .extended_lut = "off";
defparam \addr_cmd~0 .lut_mask = 64'h4000000040000000;
defparam \addr_cmd~0 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~1 (
	.dataa(!\ac_state.s_1~q ),
	.datab(!\state.s_topup_refresh~q ),
	.datac(!\state.s_refresh~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~1 .extended_lut = "off";
defparam \addr_cmd~1 .lut_mask = 64'h2A2A2A2A2A2A2A2A;
defparam \addr_cmd~1 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~2 (
	.dataa(!addr_cmd0cs_n0),
	.datab(!\state.s_run_init_seq~q ),
	.datac(!\addr_cmd~0_combout ),
	.datad(!\ac_state.s_12~q ),
	.datae(!\addr_cmd~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~2 .extended_lut = "off";
defparam \addr_cmd~2 .lut_mask = 64'h1011111110111111;
defparam \addr_cmd~2 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~3 (
	.dataa(!\state.s_program_cal_mrs~q ),
	.datab(!\ac_state.s_1~q ),
	.datac(!\ac_state.s_6~q ),
	.datad(!\WideNor1~0_combout ),
	.datae(!\ac_state.s_0~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~3 .extended_lut = "off";
defparam \addr_cmd~3 .lut_mask = 64'h5555054555550545;
defparam \addr_cmd~3 .shared_arith = "off";

arriaii_lcell_comb WideOr21(
	.dataa(!\ac_state.s_6~q ),
	.datab(!\ac_state.s_7~q ),
	.datac(!\WideOr16~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr21~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr21.extended_lut = "off";
defparam WideOr21.lut_mask = 64'h0808080808080808;
defparam WideOr21.shared_arith = "off";

arriaii_lcell_comb \addr_cmd~4 (
	.dataa(!\ac_state.s_1~q ),
	.datab(!\ac_state.s_2~q ),
	.datac(!\ac_state.s_0~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~4 .extended_lut = "off";
defparam \addr_cmd~4 .lut_mask = 64'hC4C4C4C4C4C4C4C4;
defparam \addr_cmd~4 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~5 (
	.dataa(!\state.s_run_init_seq~q ),
	.datab(!\ac_state.s_12~q ),
	.datac(!\ac_state.s_0~q ),
	.datad(!\state.s_access_precharge~q ),
	.datae(!\addr_cmd~4_combout ),
	.dataf(!\WideOr32~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~5 .extended_lut = "off";
defparam \addr_cmd~5 .lut_mask = 64'h00000000BB00BB0B;
defparam \addr_cmd~5 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~6 (
	.dataa(!\state.s_prog_user_mrs~q ),
	.datab(!\ac_state.s_0~q ),
	.datac(!\addr_cmd~3_combout ),
	.datad(!\WideOr21~combout ),
	.datae(!\addr_cmd~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~6 .extended_lut = "off";
defparam \addr_cmd~6 .lut_mask = 64'h0000A0B00000A0B0;
defparam \addr_cmd~6 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~8 (
	.dataa(!\state.s_access_act~q ),
	.datab(!\addr_cmd~0_combout ),
	.datac(!\ac_state.s_1~q ),
	.datad(!\addr_cmd~7_combout ),
	.datae(!\state.s_zq_cal_short~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~8 .extended_lut = "off";
defparam \addr_cmd~8 .lut_mask = 64'h0323030303230303;
defparam \addr_cmd~8 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~9 (
	.dataa(!addr_cmd1cs_n0),
	.datab(!\state.s_run_init_seq~q ),
	.datac(!\stage_counter~0_combout ),
	.datad(!\addr_cmd~6_combout ),
	.datae(!\addr_cmd~8_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~9 .extended_lut = "off";
defparam \addr_cmd~9 .lut_mask = 64'h1011D0DD1011D0DD;
defparam \addr_cmd~9 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~10 (
	.dataa(!addr_cmd0cke0),
	.datab(!\state.s_run_init_seq~q ),
	.datac(!\state.s_reset~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~10 .extended_lut = "off";
defparam \addr_cmd~10 .lut_mask = 64'h1D1D1D1D1D1D1D1D;
defparam \addr_cmd~10 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~11 (
	.dataa(!\state.s_run_init_seq~q ),
	.datab(!\addr_cmd~0_combout ),
	.datac(!\addr_cmd~1_combout ),
	.datad(!\ac_state.s_11~q ),
	.datae(!\addr_cmd~10_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~11 .extended_lut = "off";
defparam \addr_cmd~11 .lut_mask = 64'h2030AAFF2030AAFF;
defparam \addr_cmd~11 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~12 (
	.dataa(!\stage_counter~0_combout ),
	.datab(!\ac_state.s_12~q ),
	.datac(!\addr_cmd~10_combout ),
	.datad(!\addr_cmd~11_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~12 .extended_lut = "off";
defparam \addr_cmd~12 .lut_mask = 64'h0BFF0BFF0BFF0BFF;
defparam \addr_cmd~12 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~13 (
	.dataa(!addr_cmd0addr0),
	.datab(!addr_cmd1addr0),
	.datac(!\state.s_run_init_seq~q ),
	.datad(!\state.s_reset~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~13 .extended_lut = "off";
defparam \addr_cmd~13 .lut_mask = 64'h0035003500350035;
defparam \addr_cmd~13 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~15 (
	.dataa(!\state.s_prog_user_mrs~q ),
	.datab(!\state.s_reset~q ),
	.datac(!\addr_cmd~14_combout ),
	.datad(!\WideOr21~combout ),
	.datae(!\Selector422~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~15 .extended_lut = "off";
defparam \addr_cmd~15 .lut_mask = 64'h0000020300000203;
defparam \addr_cmd~15 .shared_arith = "off";

arriaii_lcell_comb \Selector468~0 (
	.dataa(!\addr_cmd~1_combout ),
	.datab(!\state.s_access_precharge~q ),
	.datac(!\addr_cmd~4_combout ),
	.datad(!\addr_cmd~15_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector468~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector468~0 .extended_lut = "off";
defparam \Selector468~0 .lut_mask = 64'h008A008A008A008A;
defparam \Selector468~0 .shared_arith = "off";

arriaii_lcell_comb \Selector469~0 (
	.dataa(!\state.s_program_cal_mrs~q ),
	.datab(!\state.s_prog_user_mrs~q ),
	.datac(!\state.s_access_precharge~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector469~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector469~0 .extended_lut = "off";
defparam \Selector469~0 .lut_mask = 64'h8080808080808080;
defparam \Selector469~0 .shared_arith = "off";

arriaii_lcell_comb \Selector468~1 (
	.dataa(!\state.s_run_init_seq~q ),
	.datab(!\ac_state.s_11~q ),
	.datac(!\WideOr32~combout ),
	.datad(!\process_12~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector468~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector468~1 .extended_lut = "off";
defparam \Selector468~1 .lut_mask = 64'h0E0A0E0A0E0A0E0A;
defparam \Selector468~1 .shared_arith = "off";

arriaii_lcell_comb \Selector468~2 (
	.dataa(!\ac_state.s_1~q ),
	.datab(!\addr_cmd~7_combout ),
	.datac(!\ac_state.s_0~q ),
	.datad(!\Selector469~0_combout ),
	.datae(!\Selector468~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector468~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector468~2 .extended_lut = "off";
defparam \Selector468~2 .lut_mask = 64'h00000BBB00000BBB;
defparam \Selector468~2 .shared_arith = "off";

arriaii_lcell_comb \Selector469~1 (
	.dataa(!\state.s_access_act~q ),
	.datab(!\state.s_reset~q ),
	.datac(!\ac_state.s_1~q ),
	.datad(!\state.s_zq_cal_short~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector469~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector469~1 .extended_lut = "off";
defparam \Selector469~1 .lut_mask = 64'h1030103010301030;
defparam \Selector469~1 .shared_arith = "off";

arriaii_lcell_comb \Selector469~2 (
	.dataa(!\state.s_program_cal_mrs~q ),
	.datab(!\state.s_prog_user_mrs~q ),
	.datac(!\ac_state.s_5~q ),
	.datad(!\ac_state.s_4~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector469~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector469~2 .extended_lut = "off";
defparam \Selector469~2 .lut_mask = 64'h0357035703570357;
defparam \Selector469~2 .shared_arith = "off";

arriaii_lcell_comb \Selector469~3 (
	.dataa(!addr_cmd0addr0),
	.datab(!addr_cmd1addr0),
	.datac(!\state.s_run_init_seq~q ),
	.datad(!\Selector469~1_combout ),
	.datae(!\Selector469~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector469~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector469~3 .extended_lut = "off";
defparam \Selector469~3 .lut_mask = 64'hFFCA0000FFCA0000;
defparam \Selector469~3 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~16 (
	.dataa(!addr_cmd1addr0),
	.datab(!\stage_counter~0_combout ),
	.datac(!\addr_cmd~13_combout ),
	.datad(!\Selector468~0_combout ),
	.datae(!\Selector468~2_combout ),
	.dataf(!\Selector469~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~16 .extended_lut = "off";
defparam \addr_cmd~16 .lut_mask = 64'h3F3F3F3F1F1D0F0C;
defparam \addr_cmd~16 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~17 (
	.dataa(!\state.s_reset~q ),
	.datab(!\stage_counter_zero~q ),
	.datac(!\state.s_access_precharge~q ),
	.datad(!\addr_cmd~4_combout ),
	.datae(!\addr_cmd~15_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~17 .extended_lut = "off";
defparam \addr_cmd~17 .lut_mask = 64'h5555151155551511;
defparam \addr_cmd~17 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~18 (
	.dataa(!\state.s_reset~q ),
	.datab(!\ac_state.s_1~q ),
	.datac(!\state.s_topup_refresh~q ),
	.datad(!\state.s_refresh~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~18 .extended_lut = "off";
defparam \addr_cmd~18 .lut_mask = 64'hF888F888F888F888;
defparam \addr_cmd~18 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~19 (
	.dataa(!\ac_state.s_0~q ),
	.datab(!\Selector469~0_combout ),
	.datac(!\Selector468~1_combout ),
	.datad(!\Selector469~1_combout ),
	.datae(!\addr_cmd~18_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~19 .extended_lut = "off";
defparam \addr_cmd~19 .lut_mask = 64'h0000070000000700;
defparam \addr_cmd~19 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~20 (
	.dataa(!addr_cmd1addr0),
	.datab(!\stage_counter~0_combout ),
	.datac(!\Selector469~2_combout ),
	.datad(!\addr_cmd~17_combout ),
	.datae(!\addr_cmd~19_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~20 .extended_lut = "off";
defparam \addr_cmd~20 .lut_mask = 64'h1357035713570357;
defparam \addr_cmd~20 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~21 (
	.dataa(!addr_cmd0addr1),
	.datab(!addr_cmd1addr1),
	.datac(!\state.s_run_init_seq~q ),
	.datad(!\state.s_reset~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~21 .extended_lut = "off";
defparam \addr_cmd~21 .lut_mask = 64'h0035003500350035;
defparam \addr_cmd~21 .shared_arith = "off";

arriaii_lcell_comb \Selector468~3 (
	.dataa(!\state.s_program_cal_mrs~q ),
	.datab(!\state.s_prog_user_mrs~q ),
	.datac(!\ac_state.s_4~q ),
	.datad(!\ac_state.s_3~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector468~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector468~3 .extended_lut = "off";
defparam \Selector468~3 .lut_mask = 64'h0357035703570357;
defparam \Selector468~3 .shared_arith = "off";

arriaii_lcell_comb \Selector468~4 (
	.dataa(!addr_cmd0addr1),
	.datab(!addr_cmd1addr1),
	.datac(!\state.s_run_init_seq~q ),
	.datad(!\Selector469~1_combout ),
	.datae(!\Selector468~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector468~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector468~4 .extended_lut = "off";
defparam \Selector468~4 .lut_mask = 64'hFFCA0000FFCA0000;
defparam \Selector468~4 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~22 (
	.dataa(!addr_cmd1addr1),
	.datab(!\stage_counter~0_combout ),
	.datac(!\Selector468~0_combout ),
	.datad(!\Selector468~2_combout ),
	.datae(!\addr_cmd~21_combout ),
	.dataf(!\Selector468~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~22 .extended_lut = "off";
defparam \addr_cmd~22 .lut_mask = 64'h3333FFFF1100FDFC;
defparam \addr_cmd~22 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~23 (
	.dataa(!addr_cmd1addr1),
	.datab(!\stage_counter~0_combout ),
	.datac(!\addr_cmd~17_combout ),
	.datad(!\addr_cmd~19_combout ),
	.datae(!\Selector468~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~23 .extended_lut = "off";
defparam \addr_cmd~23 .lut_mask = 64'h1505373715053737;
defparam \addr_cmd~23 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~24 (
	.dataa(!addr_cmd0addr8),
	.datab(!addr_cmd1addr8),
	.datac(!\state.s_run_init_seq~q ),
	.datad(!\state.s_reset~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~24 .extended_lut = "off";
defparam \addr_cmd~24 .lut_mask = 64'h0035003500350035;
defparam \addr_cmd~24 .shared_arith = "off";

arriaii_lcell_comb \Selector469~4 (
	.dataa(!\state.s_program_cal_mrs~q ),
	.datab(!\ac_state.s_4~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector469~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector469~4 .extended_lut = "off";
defparam \Selector469~4 .lut_mask = 64'h1111111111111111;
defparam \Selector469~4 .shared_arith = "off";

arriaii_lcell_comb \Selector461~0 (
	.dataa(!addr_cmd0addr8),
	.datab(!addr_cmd1addr8),
	.datac(!\state.s_run_init_seq~q ),
	.datad(!\Selector468~2_combout ),
	.datae(!\Selector469~1_combout ),
	.dataf(!\Selector469~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector461~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector461~0 .extended_lut = "off";
defparam \Selector461~0 .lut_mask = 64'hCCFFC8CA00000000;
defparam \Selector461~0 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~25 (
	.dataa(!\stage_counter~0_combout ),
	.datab(!\Selector468~0_combout ),
	.datac(!\addr_cmd~24_combout ),
	.datad(!\Selector461~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~25 .extended_lut = "off";
defparam \addr_cmd~25 .lut_mask = 64'h5F0E5F0E5F0E5F0E;
defparam \addr_cmd~25 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~26 (
	.dataa(!addr_cmd1addr8),
	.datab(!\stage_counter~0_combout ),
	.datac(!\Selector469~4_combout ),
	.datad(!\addr_cmd~17_combout ),
	.datae(!\addr_cmd~19_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~26 .extended_lut = "off";
defparam \addr_cmd~26 .lut_mask = 64'h1357035713570357;
defparam \addr_cmd~26 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~27 (
	.dataa(!addr_cmd0addr10),
	.datab(!addr_cmd1addr10),
	.datac(!\state.s_run_init_seq~q ),
	.datad(!\state.s_reset~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~27 .extended_lut = "off";
defparam \addr_cmd~27 .lut_mask = 64'h0035003500350035;
defparam \addr_cmd~27 .shared_arith = "off";

arriaii_lcell_comb \Selector459~0 (
	.dataa(!addr_cmd1addr10),
	.datab(!\ac_state.s_0~q ),
	.datac(!\state.s_access_precharge~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector459~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector459~0 .extended_lut = "off";
defparam \Selector459~0 .lut_mask = 64'h0707070707070707;
defparam \Selector459~0 .shared_arith = "off";

arriaii_lcell_comb \Selector459~1 (
	.dataa(!\stage_counter[17]~1_combout ),
	.datab(!\ac_state.s_1~q ),
	.datac(!\addr_cmd~7_combout ),
	.datad(!\ac_state.s_0~q ),
	.datae(!\Selector468~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector459~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector459~1 .extended_lut = "off";
defparam \Selector459~1 .lut_mask = 64'h000045CF000045CF;
defparam \Selector459~1 .shared_arith = "off";

arriaii_lcell_comb \Selector459~2 (
	.dataa(!\state.s_prog_user_mrs~q ),
	.datab(!\ac_state.s_1~q ),
	.datac(!\addr_cmd~4_combout ),
	.datad(!\Selector459~0_combout ),
	.datae(!\Selector421~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector459~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector459~2 .extended_lut = "off";
defparam \Selector459~2 .lut_mask = 64'hEEE00000EEE00000;
defparam \Selector459~2 .shared_arith = "off";

arriaii_lcell_comb \Selector459~3 (
	.dataa(!addr_cmd0addr10),
	.datab(!addr_cmd1addr10),
	.datac(!\state.s_run_init_seq~q ),
	.datad(!\Selector469~1_combout ),
	.datae(!\Selector459~1_combout ),
	.dataf(!\Selector459~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector459~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector459~3 .extended_lut = "off";
defparam \Selector459~3 .lut_mask = 64'h00000000CCC8FFCA;
defparam \Selector459~3 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~28 (
	.dataa(!\stage_counter~0_combout ),
	.datab(!\addr_cmd~1_combout ),
	.datac(!\addr_cmd~15_combout ),
	.datad(!\addr_cmd~27_combout ),
	.datae(!\Selector459~0_combout ),
	.dataf(!\Selector459~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~28 .extended_lut = "off";
defparam \addr_cmd~28 .lut_mask = 64'h55FF55FF00FB00FF;
defparam \addr_cmd~28 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~29 (
	.dataa(!\stage_counter[17]~1_combout ),
	.datab(!\ac_state.s_0~q ),
	.datac(!\Selector468~1_combout ),
	.datad(!\Selector469~1_combout ),
	.datae(!\addr_cmd~18_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~29 .extended_lut = "off";
defparam \addr_cmd~29 .lut_mask = 64'h0000070000000700;
defparam \addr_cmd~29 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~30 (
	.dataa(!addr_cmd1addr10),
	.datab(!\state.s_reset~q ),
	.datac(!\stage_counter_zero~q ),
	.datad(!\state.s_access_precharge~q ),
	.datae(!\addr_cmd~15_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~30 .extended_lut = "off";
defparam \addr_cmd~30 .lut_mask = 64'h1111011111110111;
defparam \addr_cmd~30 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~31 (
	.dataa(!addr_cmd1addr10),
	.datab(!\stage_counter~0_combout ),
	.datac(!\Selector459~2_combout ),
	.datad(!\addr_cmd~29_combout ),
	.datae(!\addr_cmd~30_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~31 .extended_lut = "off";
defparam \addr_cmd~31 .lut_mask = 64'h3130FFFF3130FFFF;
defparam \addr_cmd~31 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~32 (
	.dataa(!addr_cmd0ba0),
	.datab(!addr_cmd1ba0),
	.datac(!\state.s_run_init_seq~q ),
	.datad(!\state.s_reset~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~32 .extended_lut = "off";
defparam \addr_cmd~32 .lut_mask = 64'h0035003500350035;
defparam \addr_cmd~32 .shared_arith = "off";

arriaii_lcell_comb \Selector472~0 (
	.dataa(!\state.s_program_cal_mrs~q ),
	.datab(!\state.s_prog_user_mrs~q ),
	.datac(!\ac_state.s_4~q ),
	.datad(!\ac_state.s_2~q ),
	.datae(!\ac_state.s_3~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector472~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector472~0 .extended_lut = "off";
defparam \Selector472~0 .lut_mask = 64'hFCA88888FCA88888;
defparam \Selector472~0 .shared_arith = "off";

arriaii_lcell_comb \Selector472~1 (
	.dataa(!addr_cmd0ba0),
	.datab(!addr_cmd1ba0),
	.datac(!\state.s_run_init_seq~q ),
	.datad(!\Selector469~1_combout ),
	.datae(!\Selector472~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector472~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector472~1 .extended_lut = "off";
defparam \Selector472~1 .lut_mask = 64'h0000FFCA0000FFCA;
defparam \Selector472~1 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~33 (
	.dataa(!addr_cmd1ba0),
	.datab(!\stage_counter~0_combout ),
	.datac(!\Selector468~0_combout ),
	.datad(!\Selector468~2_combout ),
	.datae(!\addr_cmd~32_combout ),
	.dataf(!\Selector472~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~33 .extended_lut = "off";
defparam \addr_cmd~33 .lut_mask = 64'h3333FFFF1100FDFC;
defparam \addr_cmd~33 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~34 (
	.dataa(!addr_cmd1ba0),
	.datab(!\stage_counter~0_combout ),
	.datac(!\addr_cmd~17_combout ),
	.datad(!\addr_cmd~19_combout ),
	.datae(!\Selector472~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~34 .extended_lut = "off";
defparam \addr_cmd~34 .lut_mask = 64'h3737150537371505;
defparam \addr_cmd~34 .shared_arith = "off";

arriaii_lcell_comb \Selector471~0 (
	.dataa(!addr_cmd0ba1),
	.datab(!addr_cmd1ba1),
	.datac(!\state.s_run_init_seq~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector471~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector471~0 .extended_lut = "off";
defparam \Selector471~0 .lut_mask = 64'h3535353535353535;
defparam \Selector471~0 .shared_arith = "off";

arriaii_lcell_comb \Selector471~1 (
	.dataa(!\state.s_program_cal_mrs~q ),
	.datab(!\state.s_prog_user_mrs~q ),
	.datac(!\ac_state.s_1~q ),
	.datad(!\ac_state.s_2~q ),
	.datae(!\ac_state.s_3~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector471~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector471~1 .extended_lut = "off";
defparam \Selector471~1 .lut_mask = 64'hFA88C888FA88C888;
defparam \Selector471~1 .shared_arith = "off";

arriaii_lcell_comb \Selector471~2 (
	.dataa(!addr_cmd1ba1),
	.datab(!\Selector468~2_combout ),
	.datac(!\Selector469~1_combout ),
	.datad(!\Selector471~0_combout ),
	.datae(!\Selector471~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector471~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector471~2 .extended_lut = "off";
defparam \Selector471~2 .lut_mask = 64'h0000BBB00000BBB0;
defparam \Selector471~2 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~35 (
	.dataa(!\state.s_reset~q ),
	.datab(!\stage_counter~0_combout ),
	.datac(!\Selector468~0_combout ),
	.datad(!\Selector471~0_combout ),
	.datae(!\Selector471~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~35 .extended_lut = "off";
defparam \addr_cmd~35 .lut_mask = 64'h3377005433770054;
defparam \addr_cmd~35 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~36 (
	.dataa(!addr_cmd1ba1),
	.datab(!\stage_counter~0_combout ),
	.datac(!\addr_cmd~17_combout ),
	.datad(!\addr_cmd~19_combout ),
	.datae(!\Selector471~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~36 .extended_lut = "off";
defparam \addr_cmd~36 .lut_mask = 64'h3737150537371505;
defparam \addr_cmd~36 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~37 (
	.dataa(!addr_cmd1ras_n),
	.datab(!\state.s_prog_user_mrs~q ),
	.datac(!\ac_state.s_0~q ),
	.datad(!\state.s_access_precharge~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~37 .extended_lut = "off";
defparam \addr_cmd~37 .lut_mask = 64'hECA0ECA0ECA0ECA0;
defparam \addr_cmd~37 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~38 (
	.dataa(!\state.s_access_act~q ),
	.datab(!\state.s_topup_refresh~q ),
	.datac(!\state.s_refresh~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~38 .extended_lut = "off";
defparam \addr_cmd~38 .lut_mask = 64'h8080808080808080;
defparam \addr_cmd~38 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~39 (
	.dataa(!\state.s_program_cal_mrs~q ),
	.datab(!\addr_cmd~0_combout ),
	.datac(!\ac_state.s_6~q ),
	.datad(!\WideNor1~0_combout ),
	.datae(!\WideNor1~1_combout ),
	.dataf(!\addr_cmd~38_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~39 .extended_lut = "off";
defparam \addr_cmd~39 .lut_mask = 64'h0000000032323222;
defparam \addr_cmd~39 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~40 (
	.dataa(!\state.s_reset~q ),
	.datab(!\stage_counter~0_combout ),
	.datac(!\ac_state.s_1~q ),
	.datad(!\state.s_zq_cal_short~q ),
	.datae(!\addr_cmd~37_combout ),
	.dataf(!\addr_cmd~39_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~40 .extended_lut = "off";
defparam \addr_cmd~40 .lut_mask = 64'h5555555555550010;
defparam \addr_cmd~40 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~41 (
	.dataa(!addr_cmd0ras_n),
	.datab(!addr_cmd1ras_n),
	.datac(!\state.s_run_init_seq~q ),
	.datad(!\addr_cmd~40_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~41 .extended_lut = "off";
defparam \addr_cmd~41 .lut_mask = 64'h0035003500350035;
defparam \addr_cmd~41 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~42 (
	.dataa(!addr_cmd0ras_n),
	.datab(!\state.s_run_init_seq~q ),
	.datac(!\state.s_reset~q ),
	.datad(!\ac_state.s_12~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~42 .extended_lut = "off";
defparam \addr_cmd~42 .lut_mask = 64'h0001000100010001;
defparam \addr_cmd~42 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~43 (
	.dataa(!addr_cmd1ras_n),
	.datab(!\state.s_program_cal_mrs~q ),
	.datac(!\ac_state.s_0~q ),
	.datad(!\Selector468~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~43 .extended_lut = "off";
defparam \addr_cmd~43 .lut_mask = 64'h5510551055105510;
defparam \addr_cmd~43 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~44 (
	.dataa(!\state.s_prog_user_mrs~q ),
	.datab(!\WideOr21~combout ),
	.datac(!\state.s_access_precharge~q ),
	.datad(!\addr_cmd~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~44 .extended_lut = "off";
defparam \addr_cmd~44 .lut_mask = 64'h111F111F111F111F;
defparam \addr_cmd~44 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~45 (
	.dataa(!\state.s_program_cal_mrs~q ),
	.datab(!\ac_state.s_1~q ),
	.datac(!\ac_state.s_4~q ),
	.datad(!\Selector472~2_combout ),
	.datae(!\addr_cmd~38_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~45 .extended_lut = "off";
defparam \addr_cmd~45 .lut_mask = 64'h88C8AAEA88C8AAEA;
defparam \addr_cmd~45 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~46 (
	.dataa(!addr_cmd1ras_n),
	.datab(!\ac_state.s_0~q ),
	.datac(!\addr_cmd~44_combout ),
	.datad(!\addr_cmd~45_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~46 .extended_lut = "off";
defparam \addr_cmd~46 .lut_mask = 64'h00F800F800F800F8;
defparam \addr_cmd~46 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~47 (
	.dataa(!\stage_counter~0_combout ),
	.datab(!\addr_cmd~41_combout ),
	.datac(!\addr_cmd~42_combout ),
	.datad(!\addr_cmd~43_combout ),
	.datae(!\addr_cmd~46_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~47 .extended_lut = "off";
defparam \addr_cmd~47 .lut_mask = 64'h7F7F3F7F7F7F3F7F;
defparam \addr_cmd~47 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~48 (
	.dataa(!\state.s_program_cal_mrs~q ),
	.datab(!\state.s_reset~q ),
	.datac(!\ac_state.s_1~q ),
	.datad(!\ac_state.s_0~q ),
	.datae(!\state.s_zq_cal_short~q ),
	.dataf(!\Selector468~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~48 .extended_lut = "off";
defparam \addr_cmd~48 .lut_mask = 64'h00000000AAFF8ACF;
defparam \addr_cmd~48 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~49 (
	.dataa(!\state.s_prog_user_mrs~q ),
	.datab(!\state.s_access_precharge~q ),
	.datac(!\Selector595~0_combout ),
	.datad(!\addr_cmd~39_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~49 .extended_lut = "off";
defparam \addr_cmd~49 .lut_mask = 64'h0080008000800080;
defparam \addr_cmd~49 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~50 (
	.dataa(!addr_cmd1ras_n),
	.datab(!\state.s_reset~q ),
	.datac(!\stage_counter_zero~q ),
	.datad(!\addr_cmd~46_combout ),
	.datae(!\addr_cmd~48_combout ),
	.dataf(!\addr_cmd~49_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~50_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~50 .extended_lut = "off";
defparam \addr_cmd~50 .lut_mask = 64'hFD55FD11FC54FC00;
defparam \addr_cmd~50 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~51 (
	.dataa(!addr_cmd0cas_n),
	.datab(!addr_cmd1cas_n),
	.datac(!\state.s_run_init_seq~q ),
	.datad(!\state.s_reset~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~51 .extended_lut = "off";
defparam \addr_cmd~51 .lut_mask = 64'h0035003500350035;
defparam \addr_cmd~51 .shared_arith = "off";

arriaii_lcell_comb \Selector473~0 (
	.dataa(!\addr_cmd~7_combout ),
	.datab(!\state.s_access_precharge~q ),
	.datac(!\addr_cmd~4_combout ),
	.datad(!\addr_cmd~15_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector473~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector473~0 .extended_lut = "off";
defparam \Selector473~0 .lut_mask = 64'h0045004500450045;
defparam \Selector473~0 .shared_arith = "off";

arriaii_lcell_comb \Selector473~1 (
	.dataa(!addr_cmd1cas_n),
	.datab(!\state.s_program_cal_mrs~q ),
	.datac(!\ac_state.s_0~q ),
	.datad(!\state.s_access_precharge~q ),
	.datae(!\Selector468~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector473~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector473~1 .extended_lut = "off";
defparam \Selector473~1 .lut_mask = 64'h5555105055551050;
defparam \Selector473~1 .shared_arith = "off";

arriaii_lcell_comb \Selector473~2 (
	.dataa(!\state.s_program_cal_mrs~q ),
	.datab(!\ac_state.s_1~q ),
	.datac(!\addr_cmd~7_combout ),
	.datad(!\ac_state.s_4~q ),
	.datae(!\Selector472~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector473~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector473~2 .extended_lut = "off";
defparam \Selector473~2 .lut_mask = 64'h8A8ACE8A8A8ACE8A;
defparam \Selector473~2 .shared_arith = "off";

arriaii_lcell_comb \Selector473~3 (
	.dataa(!addr_cmd0cas_n),
	.datab(!addr_cmd1cas_n),
	.datac(!\state.s_run_init_seq~q ),
	.datad(!\Selector469~1_combout ),
	.datae(!\Selector473~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector473~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector473~3 .extended_lut = "off";
defparam \Selector473~3 .lut_mask = 64'h0000FFCA0000FFCA;
defparam \Selector473~3 .shared_arith = "off";

arriaii_lcell_comb \Selector473~4 (
	.dataa(!addr_cmd1cas_n),
	.datab(!\state.s_prog_user_mrs~q ),
	.datac(!\WideNor1~0_combout ),
	.datad(!\ac_state.s_0~q ),
	.datae(!\Selector473~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector473~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector473~4 .extended_lut = "off";
defparam \Selector473~4 .lut_mask = 64'h0000CECF0000CECF;
defparam \Selector473~4 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~52 (
	.dataa(!\stage_counter~0_combout ),
	.datab(!\addr_cmd~51_combout ),
	.datac(!\Selector473~0_combout ),
	.datad(!\Selector473~1_combout ),
	.datae(!\Selector473~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~52 .extended_lut = "off";
defparam \addr_cmd~52 .lut_mask = 64'h7777327777773277;
defparam \addr_cmd~52 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~53 (
	.dataa(!\stage_counter~0_combout ),
	.datab(!\ac_state.s_0~q ),
	.datac(!\Selector469~0_combout ),
	.datad(!\Selector468~1_combout ),
	.datae(!\Selector469~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~53_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~53 .extended_lut = "off";
defparam \addr_cmd~53 .lut_mask = 64'h5540555555405555;
defparam \addr_cmd~53 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~54 (
	.dataa(!\stage_counter~0_combout ),
	.datab(!\addr_cmd~7_combout ),
	.datac(!\state.s_access_precharge~q ),
	.datad(!\addr_cmd~4_combout ),
	.datae(!\addr_cmd~15_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~54_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~54 .extended_lut = "off";
defparam \addr_cmd~54 .lut_mask = 64'h0000101100001011;
defparam \addr_cmd~54 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~55 (
	.dataa(!\state.s_prog_user_mrs~q ),
	.datab(!\stage_counter~0_combout ),
	.datac(!\WideNor1~0_combout ),
	.datad(!\Selector473~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~55_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~55 .extended_lut = "off";
defparam \addr_cmd~55 .lut_mask = 64'h3310331033103310;
defparam \addr_cmd~55 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~56 (
	.dataa(!addr_cmd1cas_n),
	.datab(!\state.s_reset~q ),
	.datac(!\addr_cmd~53_combout ),
	.datad(!\addr_cmd~54_combout ),
	.datae(!\addr_cmd~55_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~56_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~56 .extended_lut = "off";
defparam \addr_cmd~56 .lut_mask = 64'h1505FFFF1505FFFF;
defparam \addr_cmd~56 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~58 (
	.dataa(!\state.s_program_cal_mrs~q ),
	.datab(!\ac_state.s_6~q ),
	.datac(!\WideNor1~0_combout ),
	.datad(!\WideNor1~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~58_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~58 .extended_lut = "off";
defparam \addr_cmd~58 .lut_mask = 64'h4440444044404440;
defparam \addr_cmd~58 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~59 (
	.dataa(!addr_cmd1we_n),
	.datab(!\ac_state.s_0~q ),
	.datac(!\addr_cmd~44_combout ),
	.datad(!\addr_cmd~57_combout ),
	.datae(!\addr_cmd~58_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~59_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~59 .extended_lut = "off";
defparam \addr_cmd~59 .lut_mask = 64'hF8008800F8008800;
defparam \addr_cmd~59 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~60 (
	.dataa(!addr_cmd1we_n),
	.datab(!\addr_cmd~0_combout ),
	.datac(!\ac_state.s_0~q ),
	.datad(!\state.s_zq_cal_short~q ),
	.datae(!\Selector469~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~60_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~60 .extended_lut = "off";
defparam \addr_cmd~60 .lut_mask = 64'h2000330020003300;
defparam \addr_cmd~60 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~61 (
	.dataa(!\state.s_reset~q ),
	.datab(!\stage_counter_zero~q ),
	.datac(!\ac_state.s_1~q ),
	.datad(!\addr_cmd~38_combout ),
	.datae(!\addr_cmd~60_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~61_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~61 .extended_lut = "off";
defparam \addr_cmd~61 .lut_mask = 64'h5555400055554000;
defparam \addr_cmd~61 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~62 (
	.dataa(!addr_cmd0we_n),
	.datab(!addr_cmd1we_n),
	.datac(!\state.s_run_init_seq~q ),
	.datad(!\state.s_reset~q ),
	.datae(!\ac_state.s_12~q ),
	.dataf(!\addr_cmd~61_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~62_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~62 .extended_lut = "off";
defparam \addr_cmd~62 .lut_mask = 64'h0000000535353535;
defparam \addr_cmd~62 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~63 (
	.dataa(!addr_cmd1we_n),
	.datab(!\stage_counter~0_combout ),
	.datac(!\Selector468~1_combout ),
	.datad(!\addr_cmd~59_combout ),
	.datae(!\addr_cmd~62_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~63_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~63 .extended_lut = "off";
defparam \addr_cmd~63 .lut_mask = 64'h3310FFFF3310FFFF;
defparam \addr_cmd~63 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~64 (
	.dataa(!\state.s_reset~q ),
	.datab(!\ac_state.s_1~q ),
	.datac(!\Selector468~1_combout ),
	.datad(!\addr_cmd~38_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~64_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~64 .extended_lut = "off";
defparam \addr_cmd~64 .lut_mask = 64'h0B0F0B0F0B0F0B0F;
defparam \addr_cmd~64 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~65 (
	.dataa(!\addr_cmd~14_combout ),
	.datab(!\stage_counter_zero~q ),
	.datac(!\state.s_zq_cal_short~q ),
	.datad(!\Selector595~0_combout ),
	.datae(!\Selector469~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~65_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~65 .extended_lut = "off";
defparam \addr_cmd~65 .lut_mask = 64'h0000400000004000;
defparam \addr_cmd~65 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~66 (
	.dataa(!addr_cmd1we_n),
	.datab(!\state.s_reset~q ),
	.datac(!\stage_counter_zero~q ),
	.datad(!\addr_cmd~59_combout ),
	.datae(!\addr_cmd~64_combout ),
	.dataf(!\addr_cmd~65_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~66_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~66 .extended_lut = "off";
defparam \addr_cmd~66 .lut_mask = 64'hFD55FD11FC54FC00;
defparam \addr_cmd~66 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~67 (
	.dataa(!\addr_cmd~14_combout ),
	.datab(!\stage_counter_zero~q ),
	.datac(!\ac_state.s_12~q ),
	.datad(!\addr_cmd~1_combout ),
	.datae(!\ac_state.s_0~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~67_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~67 .extended_lut = "off";
defparam \addr_cmd~67 .lut_mask = 64'h0000400000004000;
defparam \addr_cmd~67 .shared_arith = "off";

arriaii_lcell_comb \addr_cmd~68 (
	.dataa(!\state.s_run_init_seq~q ),
	.datab(!addr_cmd0rst_n),
	.datac(!\state.s_reset~q ),
	.datad(!\stage_counter_zero~q ),
	.datae(!\ac_state.s_0~q ),
	.dataf(!\addr_cmd~67_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\addr_cmd~68_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \addr_cmd~68 .extended_lut = "off";
defparam \addr_cmd~68 .lut_mask = 64'h0A0B1B1B0F0F1F1F;
defparam \addr_cmd~68 .shared_arith = "off";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_ctrl (
	clk,
	rst_n,
	ctl_init_fail1,
	ctl_init_success1,
	states_rrp_sweep,
	states_rdv,
	states_rrp_seek,
	states_was,
	states_adv_wr_lat,
	states_adv_rd_lat,
	states_prep_customer_mr_setup,
	master_ctrl_op_rec,
	ac_nt_0,
	dgrb_ctrl_ac_nt_good,
	Selector61,
	WideOr35,
	dgrb_ctrlcommand_done,
	curr_cmdcmd_was,
	curr_cmdcmd_write_btp,
	curr_cmdcmd_write_mtp,
	curr_ctrlcommand_ack,
	curr_cmdcmd_idle,
	curr_cmdcmd_prep_customer_mr_setup,
	curr_cmdcmd_init_dram,
	curr_cmdcmd_prog_cal_mr,
	WideOr0,
	dgwb_ctrlcommand_done,
	admin_ctrlcommand_done,
	dgrb_ctrlcommand_err,
	WideOr21,
	Selector611,
	master_ctrl_op_rec1,
	master_ctrl_op_rec2,
	master_ctrl_op_rec3,
	dgrb_ctrlcommand_ack,
	dgwb_ctrlcommand_ack,
	admin_ctrlcommand_ack,
	master_ctrl_op_rec4,
	master_ctrl_op_rec5,
	master_ctrl_op_rec6,
	Selector60,
	master_ctrl_op_rec7,
	master_ctrl_op_rec8,
	ctrl_op_reccommand_opmtp_almt,
	ctrl_op_reccommand_opsingle_bit,
	dgrb_ctrlcommand_result_5,
	dgrb_ctrlcommand_result_2,
	dgrb_ctrlcommand_result_1,
	dgrb_ctrlcommand_result_0,
	dgrb_ctrlcommand_result_3,
	dgrb_ctrlcommand_result_4,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	clk;
input 	rst_n;
output 	ctl_init_fail1;
output 	ctl_init_success1;
output 	states_rrp_sweep;
output 	states_rdv;
output 	states_rrp_seek;
output 	states_was;
output 	states_adv_wr_lat;
output 	states_adv_rd_lat;
output 	states_prep_customer_mr_setup;
output 	master_ctrl_op_rec;
output 	ac_nt_0;
input 	dgrb_ctrl_ac_nt_good;
output 	Selector61;
output 	WideOr35;
input 	dgrb_ctrlcommand_done;
output 	curr_cmdcmd_was;
output 	curr_cmdcmd_write_btp;
output 	curr_cmdcmd_write_mtp;
output 	curr_ctrlcommand_ack;
output 	curr_cmdcmd_idle;
output 	curr_cmdcmd_prep_customer_mr_setup;
output 	curr_cmdcmd_init_dram;
output 	curr_cmdcmd_prog_cal_mr;
output 	WideOr0;
input 	dgwb_ctrlcommand_done;
input 	admin_ctrlcommand_done;
input 	dgrb_ctrlcommand_err;
output 	WideOr21;
output 	Selector611;
output 	master_ctrl_op_rec1;
output 	master_ctrl_op_rec2;
output 	master_ctrl_op_rec3;
input 	dgrb_ctrlcommand_ack;
input 	dgwb_ctrlcommand_ack;
input 	admin_ctrlcommand_ack;
output 	master_ctrl_op_rec4;
output 	master_ctrl_op_rec5;
output 	master_ctrl_op_rec6;
output 	Selector60;
output 	master_ctrl_op_rec7;
output 	master_ctrl_op_rec8;
output 	ctrl_op_reccommand_opmtp_almt;
output 	ctrl_op_reccommand_opsingle_bit;
input 	dgrb_ctrlcommand_result_5;
input 	dgrb_ctrlcommand_result_2;
input 	dgrb_ctrlcommand_result_1;
input 	dgrb_ctrlcommand_result_0;
input 	dgrb_ctrlcommand_result_3;
input 	dgrb_ctrlcommand_result_4;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~2_cout ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \last_state.s_prog_cal_mr~q ;
wire \last_state.s_write_mtp~q ;
wire \last_state.s_was~q ;
wire \last_state.s_adv_wr_lat~q ;
wire \last_state.s_adv_rd_lat~q ;
wire \WideNor1~4_combout ;
wire \last_state.s_prep_customer_mr_setup~q ;
wire \hold_state~q ;
wire \hold_state~0_combout ;
wire \dll_lock_counter[4]~q ;
wire \dll_lock_counter[5]~q ;
wire \dll_lock_counter[6]~q ;
wire \dll_lock_counter[7]~q ;
wire \dll_lock_counter[9]~q ;
wire \dll_lock_counter[8]~q ;
wire \Equal0~0_combout ;
wire \mtp_almt:dvw_size_a0[5]~q ;
wire \mtp_almt:dvw_size_a0[2]~q ;
wire \mtp_almt:dvw_size_a1[2]~q ;
wire \mtp_almt:dvw_size_a0[1]~q ;
wire \mtp_almt:dvw_size_a1[1]~q ;
wire \mtp_almt:dvw_size_a0[0]~q ;
wire \mtp_almt:dvw_size_a1[0]~q ;
wire \LessThan0~0_combout ;
wire \curr_ctrl.command_result[2]~q ;
wire \curr_ctrl.command_result[1]~q ;
wire \curr_ctrl.command_result[0]~q ;
wire \Selector7~0_combout ;
wire \Selector8~0_combout ;
wire \Selector9~0_combout ;
wire \dll_lock_counter[4]~1_combout ;
wire \dll_lock_counter[5]~2_combout ;
wire \dll_lock_counter[6]~3_combout ;
wire \dll_lock_counter[9]~4_combout ;
wire \Selector1~0_combout ;
wire \curr_ctrl.command_done~q ;
wire \Selector10~0_combout ;
wire \curr_ctrl.command_err~q ;
wire \Add1~1_sumout ;
wire \timeout_counter~0_combout ;
wire \timeout_counter_clear~0_combout ;
wire \state~34_combout ;
wire \state.s_phy_initialise~q ;
wire \state~33_combout ;
wire \state.s_init_dram~q ;
wire \flag_done_timeout~0_combout ;
wire \flag_done_timeout~q ;
wire \state~48_combout ;
wire \Add7~1_sumout ;
wire \milisecond_tick_gen_count[0]~0_combout ;
wire \milisecond_tick_gen_count[0]~q ;
wire \Add7~2 ;
wire \Add7~5_sumout ;
wire \milisecond_tick_gen_count[1]~1_combout ;
wire \milisecond_tick_gen_count[1]~q ;
wire \Add7~6 ;
wire \Add7~9_sumout ;
wire \milisecond_tick_gen_count[2]~2_combout ;
wire \milisecond_tick_gen_count[2]~q ;
wire \Add7~10 ;
wire \Add7~13_sumout ;
wire \milisecond_tick_gen_count[3]~3_combout ;
wire \milisecond_tick_gen_count[3]~q ;
wire \Add7~14 ;
wire \Add7~17_sumout ;
wire \milisecond_tick_gen_count[4]~5_combout ;
wire \milisecond_tick_gen_count[4]~q ;
wire \Add7~18 ;
wire \Add7~21_sumout ;
wire \milisecond_tick_gen_count[5]~4_combout ;
wire \milisecond_tick_gen_count[5]~q ;
wire \Equal4~0_combout ;
wire \Add7~22 ;
wire \Add7~25_sumout ;
wire \milisecond_tick_gen_count[6]~12_combout ;
wire \milisecond_tick_gen_count[6]~q ;
wire \Add7~26 ;
wire \Add7~29_sumout ;
wire \milisecond_tick_gen_count[7]~13_combout ;
wire \milisecond_tick_gen_count[7]~q ;
wire \Add7~30 ;
wire \Add7~33_sumout ;
wire \milisecond_tick_gen_count[8]~14_combout ;
wire \milisecond_tick_gen_count[8]~q ;
wire \Add7~34 ;
wire \Add7~37_sumout ;
wire \milisecond_tick_gen_count[9]~15_combout ;
wire \milisecond_tick_gen_count[9]~q ;
wire \Add7~38 ;
wire \Add7~41_sumout ;
wire \milisecond_tick_gen_count[10]~17_combout ;
wire \milisecond_tick_gen_count[10]~q ;
wire \Add7~42 ;
wire \Add7~45_sumout ;
wire \milisecond_tick_gen_count[11]~16_combout ;
wire \milisecond_tick_gen_count[11]~q ;
wire \Add7~46 ;
wire \Add7~49_sumout ;
wire \milisecond_tick_gen_count[12]~6_combout ;
wire \milisecond_tick_gen_count[12]~q ;
wire \Add7~50 ;
wire \Add7~53_sumout ;
wire \milisecond_tick_gen_count[13]~7_combout ;
wire \milisecond_tick_gen_count[13]~q ;
wire \Add7~54 ;
wire \Add7~57_sumout ;
wire \milisecond_tick_gen_count[14]~8_combout ;
wire \milisecond_tick_gen_count[14]~q ;
wire \Add7~58 ;
wire \Add7~61_sumout ;
wire \milisecond_tick_gen_count[15]~9_combout ;
wire \milisecond_tick_gen_count[15]~q ;
wire \Add7~62 ;
wire \Add7~65_sumout ;
wire \milisecond_tick_gen_count[16]~11_combout ;
wire \milisecond_tick_gen_count[16]~q ;
wire \Add7~66 ;
wire \Add7~69_sumout ;
wire \milisecond_tick_gen_count[17]~10_combout ;
wire \milisecond_tick_gen_count[17]~q ;
wire \Equal4~1_combout ;
wire \Equal4~2_combout ;
wire \Equal4~3_combout ;
wire \Add6~1_sumout ;
wire \last_state.s_operational~q ;
wire \process_16~0_combout ;
wire \tracking_ms_counter[0]~0_combout ;
wire \tracking_ms_counter[0]~q ;
wire \Add6~2 ;
wire \Add6~5_sumout ;
wire \tracking_ms_counter[1]~q ;
wire \Add6~6 ;
wire \Add6~9_sumout ;
wire \tracking_ms_counter[2]~q ;
wire \Add6~10 ;
wire \Add6~13_sumout ;
wire \tracking_ms_counter[3]~q ;
wire \Add6~14 ;
wire \Add6~17_sumout ;
wire \tracking_ms_counter[4]~q ;
wire \Add6~18 ;
wire \Add6~21_sumout ;
wire \tracking_ms_counter[5]~q ;
wire \Add6~22 ;
wire \Add6~25_sumout ;
wire \tracking_ms_counter[6]~q ;
wire \Add6~26 ;
wire \Add6~29_sumout ;
wire \tracking_ms_counter~1_combout ;
wire \tracking_ms_counter[7]~q ;
wire \Equal5~0_combout ;
wire \Equal5~1_combout ;
wire \tracking_update_due~0_combout ;
wire \tracking_update_due~q ;
wire \state~31_combout ;
wire \state.s_tracking~q ;
wire \state~32_combout ;
wire \state.s_operational~q ;
wire \last_state.s_tracking~q ;
wire \last_state.s_non_operational~q ;
wire \WideNor1~5_combout ;
wire \state~49_combout ;
wire \state.s_poa~q ;
wire \last_state.s_poa~q ;
wire \state~51_combout ;
wire \state.s_tracking_setup~q ;
wire \last_state.s_tracking_setup~q ;
wire \WideNor1~6_combout ;
wire \WideNor1~7_combout ;
wire \state~38_combout ;
wire \state.s_write_mtp~q ;
wire \Selector34~0_combout ;
wire \state.s_reset~q ;
wire \state~37_combout ;
wire \state.s_cal~q ;
wire \Selector36~0_combout ;
wire \ac_nt_almts_checked~q ;
wire \mtp_almts_checked[1]~0_combout ;
wire \mtp_almts_checked[1]~q ;
wire \mtp_almt:dvw_size_a0[0]~0_combout ;
wire \mtp_almts_checked[0]~q ;
wire \state~41_combout ;
wire \state~42_combout ;
wire \state.s_read_mtp~q ;
wire \state~39_combout ;
wire \state~40_combout ;
wire \state.s_rrp_reset~q ;
wire \last_state.s_rrp_reset~q ;
wire \last_state.s_read_mtp~q ;
wire \WideNor1~2_combout ;
wire \last_state.s_rrp_sweep~q ;
wire \last_state.s_rdv~q ;
wire \last_state.s_rrp_seek~q ;
wire \WideNor1~3_combout ;
wire \timeout_counter_enable~1_combout ;
wire \timeout_counter_enable~2_combout ;
wire \timeout_counter_enable~0_combout ;
wire \timeout_counter_clear~q ;
wire \timeout_counter_enable~q ;
wire \Add1~14 ;
wire \Add1~17_sumout ;
wire \timeout_counter~11_combout ;
wire \timeout_counter[4]~q ;
wire \Add1~18 ;
wire \Add1~21_sumout ;
wire \timeout_counter~12_combout ;
wire \timeout_counter[5]~q ;
wire \Add1~22 ;
wire \Add1~25_sumout ;
wire \timeout_counter~13_combout ;
wire \timeout_counter[6]~q ;
wire \Add1~26 ;
wire \Add1~29_sumout ;
wire \timeout_counter~15_combout ;
wire \timeout_counter[7]~q ;
wire \Add1~30 ;
wire \Add1~33_sumout ;
wire \timeout_counter~14_combout ;
wire \timeout_counter[8]~q ;
wire \Equal1~1_combout ;
wire \Add1~34 ;
wire \Add1~37_sumout ;
wire \timeout_counter~4_combout ;
wire \timeout_counter[9]~q ;
wire \Add1~38 ;
wire \Add1~41_sumout ;
wire \timeout_counter~5_combout ;
wire \timeout_counter[10]~q ;
wire \Add1~42 ;
wire \Add1~45_sumout ;
wire \timeout_counter~6_combout ;
wire \timeout_counter[11]~q ;
wire \Add1~46 ;
wire \Add1~49_sumout ;
wire \timeout_counter~7_combout ;
wire \timeout_counter[12]~q ;
wire \Add1~50 ;
wire \Add1~53_sumout ;
wire \timeout_counter~9_combout ;
wire \timeout_counter[13]~q ;
wire \Add1~54 ;
wire \Add1~57_sumout ;
wire \timeout_counter~8_combout ;
wire \timeout_counter[14]~q ;
wire \Equal1~2_combout ;
wire \timeout_counter[14]~16_combout ;
wire \timeout_counter[14]~1_combout ;
wire \timeout_counter[0]~q ;
wire \Add1~2 ;
wire \Add1~5_sumout ;
wire \timeout_counter~3_combout ;
wire \timeout_counter[1]~q ;
wire \Add1~6 ;
wire \Add1~9_sumout ;
wire \timeout_counter~2_combout ;
wire \timeout_counter[2]~q ;
wire \Add1~10 ;
wire \Add1~13_sumout ;
wire \timeout_counter~10_combout ;
wire \timeout_counter[3]~q ;
wire \Equal1~0_combout ;
wire \Selector0~0_combout ;
wire \curr_ctrl.command_ack~q ;
wire \waiting_for_ack~0_combout ;
wire \waiting_for_ack~q ;
wire \flag_ack_timeout~0_combout ;
wire \flag_ack_timeout~q ;
wire \process_10~0_combout ;
wire \state~35_combout ;
wire \state.s_prog_cal_mr~q ;
wire \state~36_combout ;
wire \state.s_write_btp~q ;
wire \last_state.s_write_btp~q ;
wire \last_state.s_cal~q ;
wire \WideNor1~1_combout ;
wire \WideNor1~combout ;
wire \find_cmd~0_combout ;
wire \dll_lock_counter[0]~0_combout ;
wire \dll_lock_counter[0]~q ;
wire \dll_lock_counter[1]~5_combout ;
wire \dll_lock_counter[1]~q ;
wire \dll_lock_counter[3]~6_combout ;
wire \dll_lock_counter[3]~q ;
wire \dll_lock_counter[2]~7_combout ;
wire \dll_lock_counter[2]~q ;
wire \Equal0~1_combout ;
wire \dis_state~0_combout ;
wire \dis_state~q ;
wire \state~29_combout ;
wire \state.s_non_operational~0_combout ;
wire \state.s_non_operational~q ;
wire \Selector40~0_combout ;
wire \int_ctl_init_fail~q ;
wire \Selector39~0_combout ;
wire \int_ctl_init_success~q ;
wire \state~30_combout ;
wire \state~43_combout ;
wire \state~44_combout ;
wire \state~45_combout ;
wire \state~46_combout ;
wire \state~47_combout ;
wire \state~50_combout ;
wire \Selector33~0_combout ;
wire \master_ctrl_op_rec~1_combout ;
wire \master_ctrl_op_rec~2_combout ;
wire \master_ctrl_op_rec~3_combout ;
wire \master_ctrl_op_rec~4_combout ;
wire \master_ctrl_op_rec~5_combout ;
wire \master_ctrl_op_rec~6_combout ;
wire \last_state.s_reset~q ;
wire \last_state.s_init_dram~q ;
wire \last_state.s_phy_initialise~q ;
wire \WideNor1~0_combout ;
wire \WideNor2~0_combout ;
wire \Selector4~0_combout ;
wire \curr_ctrl.command_result[5]~q ;
wire \mtp_almt:dvw_size_a1[0]~0_combout ;
wire \mtp_almt:dvw_size_a1[5]~q ;
wire \Selector6~0_combout ;
wire \curr_ctrl.command_result[3]~q ;
wire \mtp_almt:dvw_size_a0[0]~1_combout ;
wire \mtp_almt:dvw_size_a0[3]~q ;
wire \mtp_almt:dvw_size_a1[3]~q ;
wire \Selector5~0_combout ;
wire \curr_ctrl.command_result[4]~q ;
wire \mtp_almt:dvw_size_a0[4]~q ;
wire \mtp_almt:dvw_size_a1[4]~q ;
wire \LessThan0~1_combout ;
wire \LessThan0~2_combout ;
wire \mtp_correct_almt~q ;


arriaii_lcell_comb \Add0~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dll_lock_counter[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add0~2_cout ),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h000000000000FF00;
defparam \Add0~2 .shared_arith = "off";

arriaii_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dll_lock_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000000000FF00;
defparam \Add0~5 .shared_arith = "off";

arriaii_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dll_lock_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000000000FF00;
defparam \Add0~9 .shared_arith = "off";

arriaii_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dll_lock_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000000000FF00;
defparam \Add0~13 .shared_arith = "off";

arriaii_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dll_lock_counter[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000000000FF00;
defparam \Add0~17 .shared_arith = "off";

arriaii_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dll_lock_counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000000000FF00;
defparam \Add0~21 .shared_arith = "off";

arriaii_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dll_lock_counter[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000000000FF00;
defparam \Add0~25 .shared_arith = "off";

arriaii_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dll_lock_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

arriaii_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dll_lock_counter[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

arriaii_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dll_lock_counter[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000000000FF00;
defparam \Add0~37 .shared_arith = "off";

dffeas \last_state.s_prog_cal_mr (
	.clk(clk),
	.d(\state.s_prog_cal_mr~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\last_state.s_prog_cal_mr~q ),
	.prn(vcc));
defparam \last_state.s_prog_cal_mr .is_wysiwyg = "true";
defparam \last_state.s_prog_cal_mr .power_up = "low";

dffeas \last_state.s_write_mtp (
	.clk(clk),
	.d(\state.s_write_mtp~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\last_state.s_write_mtp~q ),
	.prn(vcc));
defparam \last_state.s_write_mtp .is_wysiwyg = "true";
defparam \last_state.s_write_mtp .power_up = "low";

dffeas \last_state.s_was (
	.clk(clk),
	.d(states_was),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\last_state.s_was~q ),
	.prn(vcc));
defparam \last_state.s_was .is_wysiwyg = "true";
defparam \last_state.s_was .power_up = "low";

dffeas \last_state.s_adv_wr_lat (
	.clk(clk),
	.d(states_adv_wr_lat),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\last_state.s_adv_wr_lat~q ),
	.prn(vcc));
defparam \last_state.s_adv_wr_lat .is_wysiwyg = "true";
defparam \last_state.s_adv_wr_lat .power_up = "low";

dffeas \last_state.s_adv_rd_lat (
	.clk(clk),
	.d(states_adv_rd_lat),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\last_state.s_adv_rd_lat~q ),
	.prn(vcc));
defparam \last_state.s_adv_rd_lat .is_wysiwyg = "true";
defparam \last_state.s_adv_rd_lat .power_up = "low";

arriaii_lcell_comb \WideNor1~4 (
	.dataa(!\last_state.s_was~q ),
	.datab(!states_was),
	.datac(!\last_state.s_adv_wr_lat~q ),
	.datad(!states_adv_wr_lat),
	.datae(!\last_state.s_adv_rd_lat~q ),
	.dataf(!states_adv_rd_lat),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor1~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor1~4 .extended_lut = "off";
defparam \WideNor1~4 .lut_mask = 64'h9009000000009009;
defparam \WideNor1~4 .shared_arith = "off";

dffeas \last_state.s_prep_customer_mr_setup (
	.clk(clk),
	.d(states_prep_customer_mr_setup),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\last_state.s_prep_customer_mr_setup~q ),
	.prn(vcc));
defparam \last_state.s_prep_customer_mr_setup .is_wysiwyg = "true";
defparam \last_state.s_prep_customer_mr_setup .power_up = "low";

dffeas hold_state(
	.clk(clk),
	.d(\hold_state~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\hold_state~q ),
	.prn(vcc));
defparam hold_state.is_wysiwyg = "true";
defparam hold_state.power_up = "low";

arriaii_lcell_comb \hold_state~0 (
	.dataa(!\state.s_operational~q ),
	.datab(!\state.s_non_operational~q ),
	.datac(!\state~29_combout ),
	.datad(!\tracking_update_due~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\hold_state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \hold_state~0 .extended_lut = "off";
defparam \hold_state~0 .lut_mask = 64'h080D080D080D080D;
defparam \hold_state~0 .shared_arith = "off";

dffeas \dll_lock_counter[4] (
	.clk(clk),
	.d(\dll_lock_counter[4]~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal0~1_combout ),
	.q(\dll_lock_counter[4]~q ),
	.prn(vcc));
defparam \dll_lock_counter[4] .is_wysiwyg = "true";
defparam \dll_lock_counter[4] .power_up = "low";

dffeas \dll_lock_counter[5] (
	.clk(clk),
	.d(\dll_lock_counter[5]~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal0~1_combout ),
	.q(\dll_lock_counter[5]~q ),
	.prn(vcc));
defparam \dll_lock_counter[5] .is_wysiwyg = "true";
defparam \dll_lock_counter[5] .power_up = "low";

dffeas \dll_lock_counter[6] (
	.clk(clk),
	.d(\dll_lock_counter[6]~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal0~1_combout ),
	.q(\dll_lock_counter[6]~q ),
	.prn(vcc));
defparam \dll_lock_counter[6] .is_wysiwyg = "true";
defparam \dll_lock_counter[6] .power_up = "low";

dffeas \dll_lock_counter[7] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal0~1_combout ),
	.q(\dll_lock_counter[7]~q ),
	.prn(vcc));
defparam \dll_lock_counter[7] .is_wysiwyg = "true";
defparam \dll_lock_counter[7] .power_up = "low";

dffeas \dll_lock_counter[9] (
	.clk(clk),
	.d(\dll_lock_counter[9]~4_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal0~1_combout ),
	.q(\dll_lock_counter[9]~q ),
	.prn(vcc));
defparam \dll_lock_counter[9] .is_wysiwyg = "true";
defparam \dll_lock_counter[9] .power_up = "low";

dffeas \dll_lock_counter[8] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal0~1_combout ),
	.q(\dll_lock_counter[8]~q ),
	.prn(vcc));
defparam \dll_lock_counter[8] .is_wysiwyg = "true";
defparam \dll_lock_counter[8] .power_up = "low";

arriaii_lcell_comb \Equal0~0 (
	.dataa(!\dll_lock_counter[4]~q ),
	.datab(!\dll_lock_counter[5]~q ),
	.datac(!\dll_lock_counter[6]~q ),
	.datad(!\dll_lock_counter[7]~q ),
	.datae(!\dll_lock_counter[9]~q ),
	.dataf(!\dll_lock_counter[8]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h0000010000000000;
defparam \Equal0~0 .shared_arith = "off";

dffeas \mtp_almt:dvw_size_a0[5] (
	.clk(clk),
	.d(\curr_ctrl.command_result[5]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtp_almt:dvw_size_a0[0]~1_combout ),
	.q(\mtp_almt:dvw_size_a0[5]~q ),
	.prn(vcc));
defparam \mtp_almt:dvw_size_a0[5] .is_wysiwyg = "true";
defparam \mtp_almt:dvw_size_a0[5] .power_up = "low";

dffeas \mtp_almt:dvw_size_a0[2] (
	.clk(clk),
	.d(\curr_ctrl.command_result[2]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtp_almt:dvw_size_a0[0]~1_combout ),
	.q(\mtp_almt:dvw_size_a0[2]~q ),
	.prn(vcc));
defparam \mtp_almt:dvw_size_a0[2] .is_wysiwyg = "true";
defparam \mtp_almt:dvw_size_a0[2] .power_up = "low";

dffeas \mtp_almt:dvw_size_a1[2] (
	.clk(clk),
	.d(\curr_ctrl.command_result[2]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtp_almt:dvw_size_a1[0]~0_combout ),
	.q(\mtp_almt:dvw_size_a1[2]~q ),
	.prn(vcc));
defparam \mtp_almt:dvw_size_a1[2] .is_wysiwyg = "true";
defparam \mtp_almt:dvw_size_a1[2] .power_up = "low";

dffeas \mtp_almt:dvw_size_a0[1] (
	.clk(clk),
	.d(\curr_ctrl.command_result[1]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtp_almt:dvw_size_a0[0]~1_combout ),
	.q(\mtp_almt:dvw_size_a0[1]~q ),
	.prn(vcc));
defparam \mtp_almt:dvw_size_a0[1] .is_wysiwyg = "true";
defparam \mtp_almt:dvw_size_a0[1] .power_up = "low";

dffeas \mtp_almt:dvw_size_a1[1] (
	.clk(clk),
	.d(\curr_ctrl.command_result[1]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtp_almt:dvw_size_a1[0]~0_combout ),
	.q(\mtp_almt:dvw_size_a1[1]~q ),
	.prn(vcc));
defparam \mtp_almt:dvw_size_a1[1] .is_wysiwyg = "true";
defparam \mtp_almt:dvw_size_a1[1] .power_up = "low";

dffeas \mtp_almt:dvw_size_a0[0] (
	.clk(clk),
	.d(\curr_ctrl.command_result[0]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtp_almt:dvw_size_a0[0]~1_combout ),
	.q(\mtp_almt:dvw_size_a0[0]~q ),
	.prn(vcc));
defparam \mtp_almt:dvw_size_a0[0] .is_wysiwyg = "true";
defparam \mtp_almt:dvw_size_a0[0] .power_up = "low";

dffeas \mtp_almt:dvw_size_a1[0] (
	.clk(clk),
	.d(\curr_ctrl.command_result[0]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtp_almt:dvw_size_a1[0]~0_combout ),
	.q(\mtp_almt:dvw_size_a1[0]~q ),
	.prn(vcc));
defparam \mtp_almt:dvw_size_a1[0] .is_wysiwyg = "true";
defparam \mtp_almt:dvw_size_a1[0] .power_up = "low";

arriaii_lcell_comb \LessThan0~0 (
	.dataa(!\mtp_almt:dvw_size_a0[2]~q ),
	.datab(!\mtp_almt:dvw_size_a1[2]~q ),
	.datac(!\mtp_almt:dvw_size_a0[1]~q ),
	.datad(!\mtp_almt:dvw_size_a1[1]~q ),
	.datae(!\mtp_almt:dvw_size_a0[0]~q ),
	.dataf(!\mtp_almt:dvw_size_a1[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h22B222B2B2BB22B2;
defparam \LessThan0~0 .shared_arith = "off";

dffeas \curr_ctrl.command_result[2] (
	.clk(clk),
	.d(\Selector7~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\curr_ctrl.command_result[2]~q ),
	.prn(vcc));
defparam \curr_ctrl.command_result[2] .is_wysiwyg = "true";
defparam \curr_ctrl.command_result[2] .power_up = "low";

dffeas \curr_ctrl.command_result[1] (
	.clk(clk),
	.d(\Selector8~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\curr_ctrl.command_result[1]~q ),
	.prn(vcc));
defparam \curr_ctrl.command_result[1] .is_wysiwyg = "true";
defparam \curr_ctrl.command_result[1] .power_up = "low";

dffeas \curr_ctrl.command_result[0] (
	.clk(clk),
	.d(\Selector9~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\curr_ctrl.command_result[0]~q ),
	.prn(vcc));
defparam \curr_ctrl.command_result[0] .is_wysiwyg = "true";
defparam \curr_ctrl.command_result[0] .power_up = "low";

arriaii_lcell_comb \Selector7~0 (
	.dataa(!curr_ctrlcommand_ack),
	.datab(!curr_cmdcmd_idle),
	.datac(!WideOr0),
	.datad(!dgrb_ctrlcommand_result_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector7~0 .extended_lut = "off";
defparam \Selector7~0 .lut_mask = 64'h0001000100010001;
defparam \Selector7~0 .shared_arith = "off";

arriaii_lcell_comb \Selector8~0 (
	.dataa(!curr_ctrlcommand_ack),
	.datab(!curr_cmdcmd_idle),
	.datac(!WideOr0),
	.datad(!dgrb_ctrlcommand_result_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector8~0 .extended_lut = "off";
defparam \Selector8~0 .lut_mask = 64'h0001000100010001;
defparam \Selector8~0 .shared_arith = "off";

arriaii_lcell_comb \Selector9~0 (
	.dataa(!curr_ctrlcommand_ack),
	.datab(!curr_cmdcmd_idle),
	.datac(!WideOr0),
	.datad(!dgrb_ctrlcommand_result_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector9~0 .extended_lut = "off";
defparam \Selector9~0 .lut_mask = 64'h0001000100010001;
defparam \Selector9~0 .shared_arith = "off";

arriaii_lcell_comb \dll_lock_counter[4]~1 (
	.dataa(!\Add0~17_sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dll_lock_counter[4]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dll_lock_counter[4]~1 .extended_lut = "off";
defparam \dll_lock_counter[4]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dll_lock_counter[4]~1 .shared_arith = "off";

arriaii_lcell_comb \dll_lock_counter[5]~2 (
	.dataa(!\Add0~21_sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dll_lock_counter[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dll_lock_counter[5]~2 .extended_lut = "off";
defparam \dll_lock_counter[5]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dll_lock_counter[5]~2 .shared_arith = "off";

arriaii_lcell_comb \dll_lock_counter[6]~3 (
	.dataa(!\Add0~25_sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dll_lock_counter[6]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dll_lock_counter[6]~3 .extended_lut = "off";
defparam \dll_lock_counter[6]~3 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dll_lock_counter[6]~3 .shared_arith = "off";

arriaii_lcell_comb \dll_lock_counter[9]~4 (
	.dataa(!\Add0~37_sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dll_lock_counter[9]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dll_lock_counter[9]~4 .extended_lut = "off";
defparam \dll_lock_counter[9]~4 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dll_lock_counter[9]~4 .shared_arith = "off";

dffeas ctl_init_fail(
	.clk(clk),
	.d(\int_ctl_init_fail~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ctl_init_fail1),
	.prn(vcc));
defparam ctl_init_fail.is_wysiwyg = "true";
defparam ctl_init_fail.power_up = "low";

dffeas ctl_init_success(
	.clk(clk),
	.d(\int_ctl_init_success~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ctl_init_success1),
	.prn(vcc));
defparam ctl_init_success.is_wysiwyg = "true";
defparam ctl_init_success.power_up = "low";

dffeas \state.s_rrp_sweep (
	.clk(clk),
	.d(\state~30_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(states_rrp_sweep),
	.prn(vcc));
defparam \state.s_rrp_sweep .is_wysiwyg = "true";
defparam \state.s_rrp_sweep .power_up = "low";

dffeas \state.s_rdv (
	.clk(clk),
	.d(\state~43_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(states_rdv),
	.prn(vcc));
defparam \state.s_rdv .is_wysiwyg = "true";
defparam \state.s_rdv .power_up = "low";

dffeas \state.s_rrp_seek (
	.clk(clk),
	.d(\state~44_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(states_rrp_seek),
	.prn(vcc));
defparam \state.s_rrp_seek .is_wysiwyg = "true";
defparam \state.s_rrp_seek .power_up = "low";

dffeas \state.s_was (
	.clk(clk),
	.d(\state~45_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(states_was),
	.prn(vcc));
defparam \state.s_was .is_wysiwyg = "true";
defparam \state.s_was .power_up = "low";

dffeas \state.s_adv_wr_lat (
	.clk(clk),
	.d(\state~46_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(states_adv_wr_lat),
	.prn(vcc));
defparam \state.s_adv_wr_lat .is_wysiwyg = "true";
defparam \state.s_adv_wr_lat .power_up = "low";

dffeas \state.s_adv_rd_lat (
	.clk(clk),
	.d(\state~47_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(states_adv_rd_lat),
	.prn(vcc));
defparam \state.s_adv_rd_lat .is_wysiwyg = "true";
defparam \state.s_adv_rd_lat .power_up = "low";

dffeas \state.s_prep_customer_mr_setup (
	.clk(clk),
	.d(\state~50_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(states_prep_customer_mr_setup),
	.prn(vcc));
defparam \state.s_prep_customer_mr_setup .is_wysiwyg = "true";
defparam \state.s_prep_customer_mr_setup .power_up = "low";

arriaii_lcell_comb \master_ctrl_op_rec~0 (
	.dataa(!\state.s_reset~q ),
	.datab(!\state.s_operational~q ),
	.datac(!\state.s_non_operational~q ),
	.datad(!\WideNor1~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(master_ctrl_op_rec),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_ctrl_op_rec~0 .extended_lut = "off";
defparam \master_ctrl_op_rec~0 .lut_mask = 64'hBF00BF00BF00BF00;
defparam \master_ctrl_op_rec~0 .shared_arith = "off";

dffeas \ac_nt[0] (
	.clk(clk),
	.d(\Selector33~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state~29_combout ),
	.q(ac_nt_0),
	.prn(vcc));
defparam \ac_nt[0] .is_wysiwyg = "true";
defparam \ac_nt[0] .power_up = "low";

arriaii_lcell_comb \Selector61~0 (
	.dataa(!\state.s_reset~q ),
	.datab(!\state.s_operational~q ),
	.datac(!\state.s_non_operational~q ),
	.datad(!\state.s_phy_initialise~q ),
	.datae(!\state.s_cal~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector61),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector61~0 .extended_lut = "off";
defparam \Selector61~0 .lut_mask = 64'h4000000040000000;
defparam \Selector61~0 .shared_arith = "off";

arriaii_lcell_comb \WideOr35~0 (
	.dataa(!\state.s_init_dram~q ),
	.datab(!\state.s_prog_cal_mr~q ),
	.datac(!\state.s_write_btp~q ),
	.datad(!\state.s_write_mtp~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr35),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr35~0 .extended_lut = "off";
defparam \WideOr35~0 .lut_mask = 64'h8000800080008000;
defparam \WideOr35~0 .shared_arith = "off";

dffeas \curr_cmd.cmd_was (
	.clk(clk),
	.d(\master_ctrl_op_rec~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(curr_cmdcmd_was),
	.prn(vcc));
defparam \curr_cmd.cmd_was .is_wysiwyg = "true";
defparam \curr_cmd.cmd_was .power_up = "low";

dffeas \curr_cmd.cmd_write_btp (
	.clk(clk),
	.d(\master_ctrl_op_rec~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(curr_cmdcmd_write_btp),
	.prn(vcc));
defparam \curr_cmd.cmd_write_btp .is_wysiwyg = "true";
defparam \curr_cmd.cmd_write_btp .power_up = "low";

dffeas \curr_cmd.cmd_write_mtp (
	.clk(clk),
	.d(\master_ctrl_op_rec~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(curr_cmdcmd_write_mtp),
	.prn(vcc));
defparam \curr_cmd.cmd_write_mtp .is_wysiwyg = "true";
defparam \curr_cmd.cmd_write_mtp .power_up = "low";

arriaii_lcell_comb \curr_ctrl.command_ack~0 (
	.dataa(!curr_cmdcmd_was),
	.datab(!curr_cmdcmd_write_btp),
	.datac(!curr_cmdcmd_write_mtp),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(curr_ctrlcommand_ack),
	.sumout(),
	.cout(),
	.shareout());
defparam \curr_ctrl.command_ack~0 .extended_lut = "off";
defparam \curr_ctrl.command_ack~0 .lut_mask = 64'h8080808080808080;
defparam \curr_ctrl.command_ack~0 .shared_arith = "off";

dffeas \curr_cmd.cmd_idle (
	.clk(clk),
	.d(Selector61),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(curr_cmdcmd_idle),
	.prn(vcc));
defparam \curr_cmd.cmd_idle .is_wysiwyg = "true";
defparam \curr_cmd.cmd_idle .power_up = "low";

dffeas \curr_cmd.cmd_prep_customer_mr_setup (
	.clk(clk),
	.d(\master_ctrl_op_rec~4_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(curr_cmdcmd_prep_customer_mr_setup),
	.prn(vcc));
defparam \curr_cmd.cmd_prep_customer_mr_setup .is_wysiwyg = "true";
defparam \curr_cmd.cmd_prep_customer_mr_setup .power_up = "low";

dffeas \curr_cmd.cmd_init_dram (
	.clk(clk),
	.d(\master_ctrl_op_rec~5_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(curr_cmdcmd_init_dram),
	.prn(vcc));
defparam \curr_cmd.cmd_init_dram .is_wysiwyg = "true";
defparam \curr_cmd.cmd_init_dram .power_up = "low";

dffeas \curr_cmd.cmd_prog_cal_mr (
	.clk(clk),
	.d(\master_ctrl_op_rec~6_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(curr_cmdcmd_prog_cal_mr),
	.prn(vcc));
defparam \curr_cmd.cmd_prog_cal_mr .is_wysiwyg = "true";
defparam \curr_cmd.cmd_prog_cal_mr .power_up = "low";

arriaii_lcell_comb \WideOr0~0 (
	.dataa(!curr_cmdcmd_prep_customer_mr_setup),
	.datab(!curr_cmdcmd_init_dram),
	.datac(!curr_cmdcmd_prog_cal_mr),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h8080808080808080;
defparam \WideOr0~0 .shared_arith = "off";

arriaii_lcell_comb WideOr2(
	.dataa(!curr_ctrlcommand_ack),
	.datab(!curr_cmdcmd_idle),
	.datac(!WideOr0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr21),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr2.extended_lut = "off";
defparam WideOr2.lut_mask = 64'h0101010101010101;
defparam WideOr2.shared_arith = "off";

arriaii_lcell_comb \Selector61~1 (
	.dataa(!Selector61),
	.datab(!\WideNor1~0_combout ),
	.datac(!\WideNor1~1_combout ),
	.datad(!\WideNor1~2_combout ),
	.datae(!\WideNor1~3_combout ),
	.dataf(!\WideNor1~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector611),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector61~1 .extended_lut = "off";
defparam \Selector61~1 .lut_mask = 64'h5555555555555554;
defparam \Selector61~1 .shared_arith = "off";

arriaii_lcell_comb \master_ctrl_op_rec~7 (
	.dataa(!states_adv_wr_lat),
	.datab(!master_ctrl_op_rec),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(master_ctrl_op_rec1),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_ctrl_op_rec~7 .extended_lut = "off";
defparam \master_ctrl_op_rec~7 .lut_mask = 64'h4444444444444444;
defparam \master_ctrl_op_rec~7 .shared_arith = "off";

arriaii_lcell_comb \master_ctrl_op_rec~8 (
	.dataa(!states_rdv),
	.datab(!master_ctrl_op_rec),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(master_ctrl_op_rec2),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_ctrl_op_rec~8 .extended_lut = "off";
defparam \master_ctrl_op_rec~8 .lut_mask = 64'h4444444444444444;
defparam \master_ctrl_op_rec~8 .shared_arith = "off";

arriaii_lcell_comb \master_ctrl_op_rec~9 (
	.dataa(!\state.s_read_mtp~q ),
	.datab(!master_ctrl_op_rec),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(master_ctrl_op_rec3),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_ctrl_op_rec~9 .extended_lut = "off";
defparam \master_ctrl_op_rec~9 .lut_mask = 64'h4444444444444444;
defparam \master_ctrl_op_rec~9 .shared_arith = "off";

arriaii_lcell_comb \master_ctrl_op_rec~10 (
	.dataa(!states_rrp_seek),
	.datab(!master_ctrl_op_rec),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(master_ctrl_op_rec4),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_ctrl_op_rec~10 .extended_lut = "off";
defparam \master_ctrl_op_rec~10 .lut_mask = 64'h4444444444444444;
defparam \master_ctrl_op_rec~10 .shared_arith = "off";

arriaii_lcell_comb \master_ctrl_op_rec~11 (
	.dataa(!\state.s_rrp_reset~q ),
	.datab(!master_ctrl_op_rec),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(master_ctrl_op_rec5),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_ctrl_op_rec~11 .extended_lut = "off";
defparam \master_ctrl_op_rec~11 .lut_mask = 64'h4444444444444444;
defparam \master_ctrl_op_rec~11 .shared_arith = "off";

arriaii_lcell_comb \master_ctrl_op_rec~12 (
	.dataa(!states_rrp_sweep),
	.datab(!master_ctrl_op_rec),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(master_ctrl_op_rec6),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_ctrl_op_rec~12 .extended_lut = "off";
defparam \master_ctrl_op_rec~12 .lut_mask = 64'h4444444444444444;
defparam \master_ctrl_op_rec~12 .shared_arith = "off";

arriaii_lcell_comb \Selector60~0 (
	.dataa(!\state.s_operational~q ),
	.datab(!\state.s_non_operational~q ),
	.datac(!\state.s_tracking~q ),
	.datad(!\state.s_tracking_setup~q ),
	.datae(!\WideNor2~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector60),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector60~0 .extended_lut = "off";
defparam \Selector60~0 .lut_mask = 64'h07770FFF07770FFF;
defparam \Selector60~0 .shared_arith = "off";

arriaii_lcell_comb \master_ctrl_op_rec~13 (
	.dataa(!\state.s_poa~q ),
	.datab(!master_ctrl_op_rec),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(master_ctrl_op_rec7),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_ctrl_op_rec~13 .extended_lut = "off";
defparam \master_ctrl_op_rec~13 .lut_mask = 64'h4444444444444444;
defparam \master_ctrl_op_rec~13 .shared_arith = "off";

arriaii_lcell_comb \master_ctrl_op_rec~14 (
	.dataa(!states_adv_rd_lat),
	.datab(!master_ctrl_op_rec),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(master_ctrl_op_rec8),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_ctrl_op_rec~14 .extended_lut = "off";
defparam \master_ctrl_op_rec~14 .lut_mask = 64'h4444444444444444;
defparam \master_ctrl_op_rec~14 .shared_arith = "off";

arriaii_lcell_comb \ctrl_op_rec.command_op.mtp_almt~0 (
	.dataa(!states_rrp_sweep),
	.datab(!\state.s_read_mtp~q ),
	.datac(!\state.s_poa~q ),
	.datad(!\mtp_almts_checked[1]~q ),
	.datae(!\mtp_almts_checked[0]~q ),
	.dataf(!\mtp_correct_almt~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ctrl_op_reccommand_opmtp_almt),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_op_rec.command_op.mtp_almt~0 .extended_lut = "off";
defparam \ctrl_op_rec.command_op.mtp_almt~0 .lut_mask = 64'h00007F7F007F7F7F;
defparam \ctrl_op_rec.command_op.mtp_almt~0 .shared_arith = "off";

arriaii_lcell_comb \ctrl_op_rec.command_op.single_bit~0 (
	.dataa(!states_rrp_sweep),
	.datab(!\state.s_read_mtp~q ),
	.datac(!\state.s_poa~q ),
	.datad(!\mtp_almts_checked[1]~q ),
	.datae(!\mtp_almts_checked[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ctrl_op_reccommand_opsingle_bit),
	.sumout(),
	.cout(),
	.shareout());
defparam \ctrl_op_rec.command_op.single_bit~0 .extended_lut = "off";
defparam \ctrl_op_rec.command_op.single_bit~0 .lut_mask = 64'h7F007F7F7F007F7F;
defparam \ctrl_op_rec.command_op.single_bit~0 .shared_arith = "off";

arriaii_lcell_comb \Selector1~0 (
	.dataa(!dgrb_ctrlcommand_done),
	.datab(!curr_ctrlcommand_ack),
	.datac(!curr_cmdcmd_idle),
	.datad(!WideOr0),
	.datae(!dgwb_ctrlcommand_done),
	.dataf(!admin_ctrlcommand_done),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'h0001CCCD3301FFCD;
defparam \Selector1~0 .shared_arith = "off";

dffeas \curr_ctrl.command_done (
	.clk(clk),
	.d(\Selector1~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\curr_ctrl.command_done~q ),
	.prn(vcc));
defparam \curr_ctrl.command_done .is_wysiwyg = "true";
defparam \curr_ctrl.command_done .power_up = "low";

arriaii_lcell_comb \Selector10~0 (
	.dataa(!curr_ctrlcommand_ack),
	.datab(!curr_cmdcmd_idle),
	.datac(!WideOr0),
	.datad(!dgrb_ctrlcommand_err),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector10~0 .extended_lut = "off";
defparam \Selector10~0 .lut_mask = 64'h0001000100010001;
defparam \Selector10~0 .shared_arith = "off";

dffeas \curr_ctrl.command_err (
	.clk(clk),
	.d(\Selector10~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\curr_ctrl.command_err~q ),
	.prn(vcc));
defparam \curr_ctrl.command_err .is_wysiwyg = "true";
defparam \curr_ctrl.command_err .power_up = "low";

arriaii_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\timeout_counter[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(\Add1~2 ),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h000000000000FF00;
defparam \Add1~1 .shared_arith = "off";

arriaii_lcell_comb \timeout_counter~0 (
	.dataa(!\timeout_counter_clear~q ),
	.datab(!\Add1~1_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\timeout_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \timeout_counter~0 .extended_lut = "off";
defparam \timeout_counter~0 .lut_mask = 64'h8888888888888888;
defparam \timeout_counter~0 .shared_arith = "off";

arriaii_lcell_comb \timeout_counter_clear~0 (
	.dataa(!Selector611),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\timeout_counter_clear~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \timeout_counter_clear~0 .extended_lut = "off";
defparam \timeout_counter_clear~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \timeout_counter_clear~0 .shared_arith = "off";

arriaii_lcell_comb \state~34 (
	.dataa(!\state.s_reset~q ),
	.datab(!\state.s_phy_initialise~q ),
	.datac(!\state~29_combout ),
	.datad(!\process_10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~34 .extended_lut = "off";
defparam \state~34 .lut_mask = 64'h003A003A003A003A;
defparam \state~34 .shared_arith = "off";

dffeas \state.s_phy_initialise (
	.clk(clk),
	.d(\state~34_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_phy_initialise~q ),
	.prn(vcc));
defparam \state.s_phy_initialise .is_wysiwyg = "true";
defparam \state.s_phy_initialise .power_up = "low";

arriaii_lcell_comb \state~33 (
	.dataa(!\state.s_init_dram~q ),
	.datab(!\state.s_phy_initialise~q ),
	.datac(!\state~29_combout ),
	.datad(!\process_10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~33 .extended_lut = "off";
defparam \state~33 .lut_mask = 64'h0053005300530053;
defparam \state~33 .shared_arith = "off";

dffeas \state.s_init_dram (
	.clk(clk),
	.d(\state~33_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_init_dram~q ),
	.prn(vcc));
defparam \state.s_init_dram .is_wysiwyg = "true";
defparam \state.s_init_dram .power_up = "low";

arriaii_lcell_comb \flag_done_timeout~0 (
	.dataa(!states_rrp_sweep),
	.datab(!\state.s_init_dram~q ),
	.datac(!\flag_done_timeout~q ),
	.datad(!\Equal1~0_combout ),
	.datae(!\timeout_counter_clear~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\flag_done_timeout~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \flag_done_timeout~0 .extended_lut = "off";
defparam \flag_done_timeout~0 .lut_mask = 64'h0F8F0F0F0F8F0F0F;
defparam \flag_done_timeout~0 .shared_arith = "off";

dffeas flag_done_timeout(
	.clk(clk),
	.d(\flag_done_timeout~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\flag_done_timeout~q ),
	.prn(vcc));
defparam flag_done_timeout.is_wysiwyg = "true";
defparam flag_done_timeout.power_up = "low";

arriaii_lcell_comb \state~48 (
	.dataa(!\state.s_operational~q ),
	.datab(!\flag_done_timeout~q ),
	.datac(!\curr_ctrl.command_err~q ),
	.datad(!\flag_ack_timeout~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~48 .extended_lut = "off";
defparam \state~48 .lut_mask = 64'h4000400040004000;
defparam \state~48 .shared_arith = "off";

arriaii_lcell_comb \Add7~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\milisecond_tick_gen_count[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~1_sumout ),
	.cout(\Add7~2 ),
	.shareout());
defparam \Add7~1 .extended_lut = "off";
defparam \Add7~1 .lut_mask = 64'h00000000000000FF;
defparam \Add7~1 .shared_arith = "off";

arriaii_lcell_comb \milisecond_tick_gen_count[0]~0 (
	.dataa(!\last_state.s_operational~q ),
	.datab(!\Equal4~3_combout ),
	.datac(!\Add7~1_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\milisecond_tick_gen_count[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \milisecond_tick_gen_count[0]~0 .extended_lut = "off";
defparam \milisecond_tick_gen_count[0]~0 .lut_mask = 64'h0404040404040404;
defparam \milisecond_tick_gen_count[0]~0 .shared_arith = "off";

dffeas \milisecond_tick_gen_count[0] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[0]~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state.s_operational~q ),
	.q(\milisecond_tick_gen_count[0]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[0] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[0] .power_up = "low";

arriaii_lcell_comb \Add7~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\milisecond_tick_gen_count[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~5_sumout ),
	.cout(\Add7~6 ),
	.shareout());
defparam \Add7~5 .extended_lut = "off";
defparam \Add7~5 .lut_mask = 64'h000000000000FF00;
defparam \Add7~5 .shared_arith = "off";

arriaii_lcell_comb \milisecond_tick_gen_count[1]~1 (
	.dataa(!\last_state.s_operational~q ),
	.datab(!\tracking_update_due~q ),
	.datac(!\Equal4~3_combout ),
	.datad(!\Add7~5_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\milisecond_tick_gen_count[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \milisecond_tick_gen_count[1]~1 .extended_lut = "off";
defparam \milisecond_tick_gen_count[1]~1 .lut_mask = 64'h5101510151015101;
defparam \milisecond_tick_gen_count[1]~1 .shared_arith = "off";

dffeas \milisecond_tick_gen_count[1] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[1]~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state.s_operational~q ),
	.q(\milisecond_tick_gen_count[1]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[1] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[1] .power_up = "low";

arriaii_lcell_comb \Add7~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\milisecond_tick_gen_count[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~9_sumout ),
	.cout(\Add7~10 ),
	.shareout());
defparam \Add7~9 .extended_lut = "off";
defparam \Add7~9 .lut_mask = 64'h000000000000FF00;
defparam \Add7~9 .shared_arith = "off";

arriaii_lcell_comb \milisecond_tick_gen_count[2]~2 (
	.dataa(!\last_state.s_operational~q ),
	.datab(!\tracking_update_due~q ),
	.datac(!\Equal4~3_combout ),
	.datad(!\Add7~9_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\milisecond_tick_gen_count[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \milisecond_tick_gen_count[2]~2 .extended_lut = "off";
defparam \milisecond_tick_gen_count[2]~2 .lut_mask = 64'h5101510151015101;
defparam \milisecond_tick_gen_count[2]~2 .shared_arith = "off";

dffeas \milisecond_tick_gen_count[2] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[2]~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state.s_operational~q ),
	.q(\milisecond_tick_gen_count[2]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[2] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[2] .power_up = "low";

arriaii_lcell_comb \Add7~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\milisecond_tick_gen_count[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~13_sumout ),
	.cout(\Add7~14 ),
	.shareout());
defparam \Add7~13 .extended_lut = "off";
defparam \Add7~13 .lut_mask = 64'h000000000000FF00;
defparam \Add7~13 .shared_arith = "off";

arriaii_lcell_comb \milisecond_tick_gen_count[3]~3 (
	.dataa(!\last_state.s_operational~q ),
	.datab(!\tracking_update_due~q ),
	.datac(!\Equal4~3_combout ),
	.datad(!\Add7~13_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\milisecond_tick_gen_count[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \milisecond_tick_gen_count[3]~3 .extended_lut = "off";
defparam \milisecond_tick_gen_count[3]~3 .lut_mask = 64'h5101510151015101;
defparam \milisecond_tick_gen_count[3]~3 .shared_arith = "off";

dffeas \milisecond_tick_gen_count[3] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[3]~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state.s_operational~q ),
	.q(\milisecond_tick_gen_count[3]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[3] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[3] .power_up = "low";

arriaii_lcell_comb \Add7~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\milisecond_tick_gen_count[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~17_sumout ),
	.cout(\Add7~18 ),
	.shareout());
defparam \Add7~17 .extended_lut = "off";
defparam \Add7~17 .lut_mask = 64'h000000000000FF00;
defparam \Add7~17 .shared_arith = "off";

arriaii_lcell_comb \milisecond_tick_gen_count[4]~5 (
	.dataa(!\last_state.s_operational~q ),
	.datab(!\tracking_update_due~q ),
	.datac(!\Equal4~3_combout ),
	.datad(!\Add7~17_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\milisecond_tick_gen_count[4]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \milisecond_tick_gen_count[4]~5 .extended_lut = "off";
defparam \milisecond_tick_gen_count[4]~5 .lut_mask = 64'h5101510151015101;
defparam \milisecond_tick_gen_count[4]~5 .shared_arith = "off";

dffeas \milisecond_tick_gen_count[4] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[4]~5_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state.s_operational~q ),
	.q(\milisecond_tick_gen_count[4]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[4] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[4] .power_up = "low";

arriaii_lcell_comb \Add7~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\milisecond_tick_gen_count[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~21_sumout ),
	.cout(\Add7~22 ),
	.shareout());
defparam \Add7~21 .extended_lut = "off";
defparam \Add7~21 .lut_mask = 64'h000000000000FF00;
defparam \Add7~21 .shared_arith = "off";

arriaii_lcell_comb \milisecond_tick_gen_count[5]~4 (
	.dataa(!\last_state.s_operational~q ),
	.datab(!\tracking_update_due~q ),
	.datac(!\Equal4~3_combout ),
	.datad(!\Add7~21_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\milisecond_tick_gen_count[5]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \milisecond_tick_gen_count[5]~4 .extended_lut = "off";
defparam \milisecond_tick_gen_count[5]~4 .lut_mask = 64'h5101510151015101;
defparam \milisecond_tick_gen_count[5]~4 .shared_arith = "off";

dffeas \milisecond_tick_gen_count[5] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[5]~4_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state.s_operational~q ),
	.q(\milisecond_tick_gen_count[5]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[5] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[5] .power_up = "low";

arriaii_lcell_comb \Equal4~0 (
	.dataa(!\milisecond_tick_gen_count[1]~q ),
	.datab(!\milisecond_tick_gen_count[2]~q ),
	.datac(!\milisecond_tick_gen_count[3]~q ),
	.datad(!\milisecond_tick_gen_count[5]~q ),
	.datae(!\milisecond_tick_gen_count[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~0 .extended_lut = "off";
defparam \Equal4~0 .lut_mask = 64'h0000000100000001;
defparam \Equal4~0 .shared_arith = "off";

arriaii_lcell_comb \Add7~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\milisecond_tick_gen_count[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~25_sumout ),
	.cout(\Add7~26 ),
	.shareout());
defparam \Add7~25 .extended_lut = "off";
defparam \Add7~25 .lut_mask = 64'h000000000000FF00;
defparam \Add7~25 .shared_arith = "off";

arriaii_lcell_comb \milisecond_tick_gen_count[6]~12 (
	.dataa(!\last_state.s_operational~q ),
	.datab(!\tracking_update_due~q ),
	.datac(!\Equal4~3_combout ),
	.datad(!\Add7~25_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\milisecond_tick_gen_count[6]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \milisecond_tick_gen_count[6]~12 .extended_lut = "off";
defparam \milisecond_tick_gen_count[6]~12 .lut_mask = 64'h5101510151015101;
defparam \milisecond_tick_gen_count[6]~12 .shared_arith = "off";

dffeas \milisecond_tick_gen_count[6] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[6]~12_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state.s_operational~q ),
	.q(\milisecond_tick_gen_count[6]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[6] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[6] .power_up = "low";

arriaii_lcell_comb \Add7~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\milisecond_tick_gen_count[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~29_sumout ),
	.cout(\Add7~30 ),
	.shareout());
defparam \Add7~29 .extended_lut = "off";
defparam \Add7~29 .lut_mask = 64'h000000000000FF00;
defparam \Add7~29 .shared_arith = "off";

arriaii_lcell_comb \milisecond_tick_gen_count[7]~13 (
	.dataa(!\last_state.s_operational~q ),
	.datab(!\tracking_update_due~q ),
	.datac(!\Equal4~3_combout ),
	.datad(!\Add7~29_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\milisecond_tick_gen_count[7]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \milisecond_tick_gen_count[7]~13 .extended_lut = "off";
defparam \milisecond_tick_gen_count[7]~13 .lut_mask = 64'h5101510151015101;
defparam \milisecond_tick_gen_count[7]~13 .shared_arith = "off";

dffeas \milisecond_tick_gen_count[7] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[7]~13_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state.s_operational~q ),
	.q(\milisecond_tick_gen_count[7]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[7] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[7] .power_up = "low";

arriaii_lcell_comb \Add7~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\milisecond_tick_gen_count[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~33_sumout ),
	.cout(\Add7~34 ),
	.shareout());
defparam \Add7~33 .extended_lut = "off";
defparam \Add7~33 .lut_mask = 64'h000000000000FF00;
defparam \Add7~33 .shared_arith = "off";

arriaii_lcell_comb \milisecond_tick_gen_count[8]~14 (
	.dataa(!\last_state.s_operational~q ),
	.datab(!\tracking_update_due~q ),
	.datac(!\Equal4~3_combout ),
	.datad(!\Add7~33_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\milisecond_tick_gen_count[8]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \milisecond_tick_gen_count[8]~14 .extended_lut = "off";
defparam \milisecond_tick_gen_count[8]~14 .lut_mask = 64'h5101510151015101;
defparam \milisecond_tick_gen_count[8]~14 .shared_arith = "off";

dffeas \milisecond_tick_gen_count[8] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[8]~14_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state.s_operational~q ),
	.q(\milisecond_tick_gen_count[8]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[8] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[8] .power_up = "low";

arriaii_lcell_comb \Add7~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\milisecond_tick_gen_count[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~37_sumout ),
	.cout(\Add7~38 ),
	.shareout());
defparam \Add7~37 .extended_lut = "off";
defparam \Add7~37 .lut_mask = 64'h00000000000000FF;
defparam \Add7~37 .shared_arith = "off";

arriaii_lcell_comb \milisecond_tick_gen_count[9]~15 (
	.dataa(!\last_state.s_operational~q ),
	.datab(!\Equal4~3_combout ),
	.datac(!\Add7~37_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\milisecond_tick_gen_count[9]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \milisecond_tick_gen_count[9]~15 .extended_lut = "off";
defparam \milisecond_tick_gen_count[9]~15 .lut_mask = 64'h0404040404040404;
defparam \milisecond_tick_gen_count[9]~15 .shared_arith = "off";

dffeas \milisecond_tick_gen_count[9] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[9]~15_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state.s_operational~q ),
	.q(\milisecond_tick_gen_count[9]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[9] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[9] .power_up = "low";

arriaii_lcell_comb \Add7~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\milisecond_tick_gen_count[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~41_sumout ),
	.cout(\Add7~42 ),
	.shareout());
defparam \Add7~41 .extended_lut = "off";
defparam \Add7~41 .lut_mask = 64'h00000000000000FF;
defparam \Add7~41 .shared_arith = "off";

arriaii_lcell_comb \milisecond_tick_gen_count[10]~17 (
	.dataa(!\last_state.s_operational~q ),
	.datab(!\Equal4~3_combout ),
	.datac(!\Add7~41_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\milisecond_tick_gen_count[10]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \milisecond_tick_gen_count[10]~17 .extended_lut = "off";
defparam \milisecond_tick_gen_count[10]~17 .lut_mask = 64'h0404040404040404;
defparam \milisecond_tick_gen_count[10]~17 .shared_arith = "off";

dffeas \milisecond_tick_gen_count[10] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[10]~17_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state.s_operational~q ),
	.q(\milisecond_tick_gen_count[10]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[10] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[10] .power_up = "low";

arriaii_lcell_comb \Add7~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\milisecond_tick_gen_count[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~45_sumout ),
	.cout(\Add7~46 ),
	.shareout());
defparam \Add7~45 .extended_lut = "off";
defparam \Add7~45 .lut_mask = 64'h000000000000FF00;
defparam \Add7~45 .shared_arith = "off";

arriaii_lcell_comb \milisecond_tick_gen_count[11]~16 (
	.dataa(!\last_state.s_operational~q ),
	.datab(!\tracking_update_due~q ),
	.datac(!\Equal4~3_combout ),
	.datad(!\Add7~45_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\milisecond_tick_gen_count[11]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \milisecond_tick_gen_count[11]~16 .extended_lut = "off";
defparam \milisecond_tick_gen_count[11]~16 .lut_mask = 64'h5101510151015101;
defparam \milisecond_tick_gen_count[11]~16 .shared_arith = "off";

dffeas \milisecond_tick_gen_count[11] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[11]~16_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state.s_operational~q ),
	.q(\milisecond_tick_gen_count[11]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[11] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[11] .power_up = "low";

arriaii_lcell_comb \Add7~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\milisecond_tick_gen_count[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~49_sumout ),
	.cout(\Add7~50 ),
	.shareout());
defparam \Add7~49 .extended_lut = "off";
defparam \Add7~49 .lut_mask = 64'h00000000000000FF;
defparam \Add7~49 .shared_arith = "off";

arriaii_lcell_comb \milisecond_tick_gen_count[12]~6 (
	.dataa(!\last_state.s_operational~q ),
	.datab(!\Equal4~3_combout ),
	.datac(!\Add7~49_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\milisecond_tick_gen_count[12]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \milisecond_tick_gen_count[12]~6 .extended_lut = "off";
defparam \milisecond_tick_gen_count[12]~6 .lut_mask = 64'h0404040404040404;
defparam \milisecond_tick_gen_count[12]~6 .shared_arith = "off";

dffeas \milisecond_tick_gen_count[12] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[12]~6_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state.s_operational~q ),
	.q(\milisecond_tick_gen_count[12]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[12] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[12] .power_up = "low";

arriaii_lcell_comb \Add7~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\milisecond_tick_gen_count[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~53_sumout ),
	.cout(\Add7~54 ),
	.shareout());
defparam \Add7~53 .extended_lut = "off";
defparam \Add7~53 .lut_mask = 64'h00000000000000FF;
defparam \Add7~53 .shared_arith = "off";

arriaii_lcell_comb \milisecond_tick_gen_count[13]~7 (
	.dataa(!\last_state.s_operational~q ),
	.datab(!\Equal4~3_combout ),
	.datac(!\Add7~53_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\milisecond_tick_gen_count[13]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \milisecond_tick_gen_count[13]~7 .extended_lut = "off";
defparam \milisecond_tick_gen_count[13]~7 .lut_mask = 64'h0404040404040404;
defparam \milisecond_tick_gen_count[13]~7 .shared_arith = "off";

dffeas \milisecond_tick_gen_count[13] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[13]~7_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state.s_operational~q ),
	.q(\milisecond_tick_gen_count[13]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[13] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[13] .power_up = "low";

arriaii_lcell_comb \Add7~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\milisecond_tick_gen_count[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~57_sumout ),
	.cout(\Add7~58 ),
	.shareout());
defparam \Add7~57 .extended_lut = "off";
defparam \Add7~57 .lut_mask = 64'h000000000000FF00;
defparam \Add7~57 .shared_arith = "off";

arriaii_lcell_comb \milisecond_tick_gen_count[14]~8 (
	.dataa(!\last_state.s_operational~q ),
	.datab(!\tracking_update_due~q ),
	.datac(!\Equal4~3_combout ),
	.datad(!\Add7~57_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\milisecond_tick_gen_count[14]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \milisecond_tick_gen_count[14]~8 .extended_lut = "off";
defparam \milisecond_tick_gen_count[14]~8 .lut_mask = 64'h5101510151015101;
defparam \milisecond_tick_gen_count[14]~8 .shared_arith = "off";

dffeas \milisecond_tick_gen_count[14] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[14]~8_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state.s_operational~q ),
	.q(\milisecond_tick_gen_count[14]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[14] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[14] .power_up = "low";

arriaii_lcell_comb \Add7~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\milisecond_tick_gen_count[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~61_sumout ),
	.cout(\Add7~62 ),
	.shareout());
defparam \Add7~61 .extended_lut = "off";
defparam \Add7~61 .lut_mask = 64'h00000000000000FF;
defparam \Add7~61 .shared_arith = "off";

arriaii_lcell_comb \milisecond_tick_gen_count[15]~9 (
	.dataa(!\last_state.s_operational~q ),
	.datab(!\Equal4~3_combout ),
	.datac(!\Add7~61_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\milisecond_tick_gen_count[15]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \milisecond_tick_gen_count[15]~9 .extended_lut = "off";
defparam \milisecond_tick_gen_count[15]~9 .lut_mask = 64'h0404040404040404;
defparam \milisecond_tick_gen_count[15]~9 .shared_arith = "off";

dffeas \milisecond_tick_gen_count[15] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[15]~9_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state.s_operational~q ),
	.q(\milisecond_tick_gen_count[15]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[15] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[15] .power_up = "low";

arriaii_lcell_comb \Add7~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\milisecond_tick_gen_count[16]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~65_sumout ),
	.cout(\Add7~66 ),
	.shareout());
defparam \Add7~65 .extended_lut = "off";
defparam \Add7~65 .lut_mask = 64'h00000000000000FF;
defparam \Add7~65 .shared_arith = "off";

arriaii_lcell_comb \milisecond_tick_gen_count[16]~11 (
	.dataa(!\last_state.s_operational~q ),
	.datab(!\Equal4~3_combout ),
	.datac(!\Add7~65_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\milisecond_tick_gen_count[16]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \milisecond_tick_gen_count[16]~11 .extended_lut = "off";
defparam \milisecond_tick_gen_count[16]~11 .lut_mask = 64'h0404040404040404;
defparam \milisecond_tick_gen_count[16]~11 .shared_arith = "off";

dffeas \milisecond_tick_gen_count[16] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[16]~11_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state.s_operational~q ),
	.q(\milisecond_tick_gen_count[16]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[16] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[16] .power_up = "low";

arriaii_lcell_comb \Add7~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\milisecond_tick_gen_count[17]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~69_sumout ),
	.cout(),
	.shareout());
defparam \Add7~69 .extended_lut = "off";
defparam \Add7~69 .lut_mask = 64'h000000000000FF00;
defparam \Add7~69 .shared_arith = "off";

arriaii_lcell_comb \milisecond_tick_gen_count[17]~10 (
	.dataa(!\last_state.s_operational~q ),
	.datab(!\tracking_update_due~q ),
	.datac(!\Equal4~3_combout ),
	.datad(!\Add7~69_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\milisecond_tick_gen_count[17]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \milisecond_tick_gen_count[17]~10 .extended_lut = "off";
defparam \milisecond_tick_gen_count[17]~10 .lut_mask = 64'h5101510151015101;
defparam \milisecond_tick_gen_count[17]~10 .shared_arith = "off";

dffeas \milisecond_tick_gen_count[17] (
	.clk(clk),
	.d(\milisecond_tick_gen_count[17]~10_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state.s_operational~q ),
	.q(\milisecond_tick_gen_count[17]~q ),
	.prn(vcc));
defparam \milisecond_tick_gen_count[17] .is_wysiwyg = "true";
defparam \milisecond_tick_gen_count[17] .power_up = "low";

arriaii_lcell_comb \Equal4~1 (
	.dataa(!\milisecond_tick_gen_count[13]~q ),
	.datab(!\milisecond_tick_gen_count[14]~q ),
	.datac(!\milisecond_tick_gen_count[15]~q ),
	.datad(!\milisecond_tick_gen_count[17]~q ),
	.datae(!\milisecond_tick_gen_count[16]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~1 .extended_lut = "off";
defparam \Equal4~1 .lut_mask = 64'h0020000000200000;
defparam \Equal4~1 .shared_arith = "off";

arriaii_lcell_comb \Equal4~2 (
	.dataa(!\milisecond_tick_gen_count[7]~q ),
	.datab(!\milisecond_tick_gen_count[8]~q ),
	.datac(!\milisecond_tick_gen_count[9]~q ),
	.datad(!\milisecond_tick_gen_count[11]~q ),
	.datae(!\milisecond_tick_gen_count[10]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~2 .extended_lut = "off";
defparam \Equal4~2 .lut_mask = 64'h0010000000100000;
defparam \Equal4~2 .shared_arith = "off";

arriaii_lcell_comb \Equal4~3 (
	.dataa(!\milisecond_tick_gen_count[0]~q ),
	.datab(!\Equal4~0_combout ),
	.datac(!\milisecond_tick_gen_count[12]~q ),
	.datad(!\Equal4~1_combout ),
	.datae(!\milisecond_tick_gen_count[6]~q ),
	.dataf(!\Equal4~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~3 .extended_lut = "off";
defparam \Equal4~3 .lut_mask = 64'h0000000000000020;
defparam \Equal4~3 .shared_arith = "off";

arriaii_lcell_comb \Add6~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\tracking_ms_counter[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~1_sumout ),
	.cout(\Add6~2 ),
	.shareout());
defparam \Add6~1 .extended_lut = "off";
defparam \Add6~1 .lut_mask = 64'h00000000000000FF;
defparam \Add6~1 .shared_arith = "off";

dffeas \last_state.s_operational (
	.clk(clk),
	.d(\state.s_operational~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\last_state.s_operational~q ),
	.prn(vcc));
defparam \last_state.s_operational .is_wysiwyg = "true";
defparam \last_state.s_operational .power_up = "low";

arriaii_lcell_comb \process_16~0 (
	.dataa(!\state.s_operational~q ),
	.datab(!\last_state.s_operational~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\process_16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \process_16~0 .extended_lut = "off";
defparam \process_16~0 .lut_mask = 64'h4444444444444444;
defparam \process_16~0 .shared_arith = "off";

arriaii_lcell_comb \tracking_ms_counter[0]~0 (
	.dataa(!\state.s_operational~q ),
	.datab(!\last_state.s_operational~q ),
	.datac(!\tracking_update_due~q ),
	.datad(!\Equal4~3_combout ),
	.datae(!\Equal5~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\tracking_ms_counter[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \tracking_ms_counter[0]~0 .extended_lut = "off";
defparam \tracking_ms_counter[0]~0 .lut_mask = 64'h4454444444544444;
defparam \tracking_ms_counter[0]~0 .shared_arith = "off";

dffeas \tracking_ms_counter[0] (
	.clk(clk),
	.d(\Add6~1_sumout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_16~0_combout ),
	.ena(\tracking_ms_counter[0]~0_combout ),
	.q(\tracking_ms_counter[0]~q ),
	.prn(vcc));
defparam \tracking_ms_counter[0] .is_wysiwyg = "true";
defparam \tracking_ms_counter[0] .power_up = "low";

arriaii_lcell_comb \Add6~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\tracking_ms_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~5_sumout ),
	.cout(\Add6~6 ),
	.shareout());
defparam \Add6~5 .extended_lut = "off";
defparam \Add6~5 .lut_mask = 64'h00000000000000FF;
defparam \Add6~5 .shared_arith = "off";

dffeas \tracking_ms_counter[1] (
	.clk(clk),
	.d(\Add6~5_sumout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_16~0_combout ),
	.ena(\tracking_ms_counter[0]~0_combout ),
	.q(\tracking_ms_counter[1]~q ),
	.prn(vcc));
defparam \tracking_ms_counter[1] .is_wysiwyg = "true";
defparam \tracking_ms_counter[1] .power_up = "low";

arriaii_lcell_comb \Add6~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\tracking_ms_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~9_sumout ),
	.cout(\Add6~10 ),
	.shareout());
defparam \Add6~9 .extended_lut = "off";
defparam \Add6~9 .lut_mask = 64'h00000000000000FF;
defparam \Add6~9 .shared_arith = "off";

dffeas \tracking_ms_counter[2] (
	.clk(clk),
	.d(\Add6~9_sumout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_16~0_combout ),
	.ena(\tracking_ms_counter[0]~0_combout ),
	.q(\tracking_ms_counter[2]~q ),
	.prn(vcc));
defparam \tracking_ms_counter[2] .is_wysiwyg = "true";
defparam \tracking_ms_counter[2] .power_up = "low";

arriaii_lcell_comb \Add6~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\tracking_ms_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~13_sumout ),
	.cout(\Add6~14 ),
	.shareout());
defparam \Add6~13 .extended_lut = "off";
defparam \Add6~13 .lut_mask = 64'h00000000000000FF;
defparam \Add6~13 .shared_arith = "off";

dffeas \tracking_ms_counter[3] (
	.clk(clk),
	.d(\Add6~13_sumout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_16~0_combout ),
	.ena(\tracking_ms_counter[0]~0_combout ),
	.q(\tracking_ms_counter[3]~q ),
	.prn(vcc));
defparam \tracking_ms_counter[3] .is_wysiwyg = "true";
defparam \tracking_ms_counter[3] .power_up = "low";

arriaii_lcell_comb \Add6~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\tracking_ms_counter[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~17_sumout ),
	.cout(\Add6~18 ),
	.shareout());
defparam \Add6~17 .extended_lut = "off";
defparam \Add6~17 .lut_mask = 64'h00000000000000FF;
defparam \Add6~17 .shared_arith = "off";

dffeas \tracking_ms_counter[4] (
	.clk(clk),
	.d(\Add6~17_sumout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_16~0_combout ),
	.ena(\tracking_ms_counter[0]~0_combout ),
	.q(\tracking_ms_counter[4]~q ),
	.prn(vcc));
defparam \tracking_ms_counter[4] .is_wysiwyg = "true";
defparam \tracking_ms_counter[4] .power_up = "low";

arriaii_lcell_comb \Add6~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\tracking_ms_counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~21_sumout ),
	.cout(\Add6~22 ),
	.shareout());
defparam \Add6~21 .extended_lut = "off";
defparam \Add6~21 .lut_mask = 64'h00000000000000FF;
defparam \Add6~21 .shared_arith = "off";

dffeas \tracking_ms_counter[5] (
	.clk(clk),
	.d(\Add6~21_sumout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_16~0_combout ),
	.ena(\tracking_ms_counter[0]~0_combout ),
	.q(\tracking_ms_counter[5]~q ),
	.prn(vcc));
defparam \tracking_ms_counter[5] .is_wysiwyg = "true";
defparam \tracking_ms_counter[5] .power_up = "low";

arriaii_lcell_comb \Add6~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\tracking_ms_counter[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~25_sumout ),
	.cout(\Add6~26 ),
	.shareout());
defparam \Add6~25 .extended_lut = "off";
defparam \Add6~25 .lut_mask = 64'h00000000000000FF;
defparam \Add6~25 .shared_arith = "off";

dffeas \tracking_ms_counter[6] (
	.clk(clk),
	.d(\Add6~25_sumout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_16~0_combout ),
	.ena(\tracking_ms_counter[0]~0_combout ),
	.q(\tracking_ms_counter[6]~q ),
	.prn(vcc));
defparam \tracking_ms_counter[6] .is_wysiwyg = "true";
defparam \tracking_ms_counter[6] .power_up = "low";

arriaii_lcell_comb \Add6~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\tracking_ms_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~29_sumout ),
	.cout(),
	.shareout());
defparam \Add6~29 .extended_lut = "off";
defparam \Add6~29 .lut_mask = 64'h00000000000000FF;
defparam \Add6~29 .shared_arith = "off";

arriaii_lcell_comb \tracking_ms_counter~1 (
	.dataa(!\state.s_operational~q ),
	.datab(!\tracking_update_due~q ),
	.datac(!\Equal4~3_combout ),
	.datad(!\tracking_ms_counter[7]~q ),
	.datae(!\Equal5~1_combout ),
	.dataf(!\Add6~29_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\tracking_ms_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \tracking_ms_counter~1 .extended_lut = "off";
defparam \tracking_ms_counter~1 .lut_mask = 64'h00FB00FB04FF00FB;
defparam \tracking_ms_counter~1 .shared_arith = "off";

dffeas \tracking_ms_counter[7] (
	.clk(clk),
	.d(\tracking_ms_counter~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_16~0_combout ),
	.ena(vcc),
	.q(\tracking_ms_counter[7]~q ),
	.prn(vcc));
defparam \tracking_ms_counter[7] .is_wysiwyg = "true";
defparam \tracking_ms_counter[7] .power_up = "low";

arriaii_lcell_comb \Equal5~0 (
	.dataa(!\tracking_ms_counter[4]~q ),
	.datab(!\tracking_ms_counter[5]~q ),
	.datac(!\tracking_ms_counter[7]~q ),
	.datad(!\tracking_ms_counter[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal5~0 .extended_lut = "off";
defparam \Equal5~0 .lut_mask = 64'h8000800080008000;
defparam \Equal5~0 .shared_arith = "off";

arriaii_lcell_comb \Equal5~1 (
	.dataa(!\tracking_ms_counter[2]~q ),
	.datab(!\tracking_ms_counter[3]~q ),
	.datac(!\Equal5~0_combout ),
	.datad(!\tracking_ms_counter[1]~q ),
	.datae(!\tracking_ms_counter[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal5~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal5~1 .extended_lut = "off";
defparam \Equal5~1 .lut_mask = 64'h0800000008000000;
defparam \Equal5~1 .shared_arith = "off";

arriaii_lcell_comb \tracking_update_due~0 (
	.dataa(!\tracking_update_due~q ),
	.datab(!\Equal4~3_combout ),
	.datac(!\Equal5~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\tracking_update_due~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \tracking_update_due~0 .extended_lut = "off";
defparam \tracking_update_due~0 .lut_mask = 64'h5757575757575757;
defparam \tracking_update_due~0 .shared_arith = "off";

dffeas tracking_update_due(
	.clk(clk),
	.d(\tracking_update_due~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\state.s_operational~q ),
	.sload(gnd),
	.ena(!\process_16~0_combout ),
	.q(\tracking_update_due~q ),
	.prn(vcc));
defparam tracking_update_due.is_wysiwyg = "true";
defparam tracking_update_due.power_up = "low";

arriaii_lcell_comb \state~31 (
	.dataa(!\state.s_operational~q ),
	.datab(!\state.s_non_operational~q ),
	.datac(!\state~29_combout ),
	.datad(!\process_10~0_combout ),
	.datae(!\tracking_update_due~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~31 .extended_lut = "off";
defparam \state~31 .lut_mask = 64'hFF08FF0CFF08FF0C;
defparam \state~31 .shared_arith = "off";

dffeas \state.s_tracking (
	.clk(clk),
	.d(\state~48_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state~31_combout ),
	.q(\state.s_tracking~q ),
	.prn(vcc));
defparam \state.s_tracking .is_wysiwyg = "true";
defparam \state.s_tracking .power_up = "low";

arriaii_lcell_comb \state~32 (
	.dataa(!\state.s_operational~q ),
	.datab(!\state.s_tracking~q ),
	.datac(!states_prep_customer_mr_setup),
	.datad(!\state~29_combout ),
	.datae(!\process_10~0_combout ),
	.dataf(!\tracking_update_due~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~32 .extended_lut = "off";
defparam \state~32 .lut_mask = 64'h0000557F0000553F;
defparam \state~32 .shared_arith = "off";

dffeas \state.s_operational (
	.clk(clk),
	.d(\state~32_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_operational~q ),
	.prn(vcc));
defparam \state.s_operational .is_wysiwyg = "true";
defparam \state.s_operational .power_up = "low";

dffeas \last_state.s_tracking (
	.clk(clk),
	.d(\state.s_tracking~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\last_state.s_tracking~q ),
	.prn(vcc));
defparam \last_state.s_tracking .is_wysiwyg = "true";
defparam \last_state.s_tracking .power_up = "low";

dffeas \last_state.s_non_operational (
	.clk(clk),
	.d(\state.s_non_operational~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\last_state.s_non_operational~q ),
	.prn(vcc));
defparam \last_state.s_non_operational .is_wysiwyg = "true";
defparam \last_state.s_non_operational .power_up = "low";

arriaii_lcell_comb \WideNor1~5 (
	.dataa(!\state.s_operational~q ),
	.datab(!\state.s_non_operational~q ),
	.datac(!\last_state.s_tracking~q ),
	.datad(!\state.s_tracking~q ),
	.datae(!\last_state.s_non_operational~q ),
	.dataf(!\last_state.s_operational~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor1~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor1~5 .extended_lut = "off";
defparam \WideNor1~5 .lut_mask = 64'h8008200240041001;
defparam \WideNor1~5 .shared_arith = "off";

arriaii_lcell_comb \state~49 (
	.dataa(!states_adv_wr_lat),
	.datab(!\state.s_poa~q ),
	.datac(!\state~29_combout ),
	.datad(!\process_10~0_combout ),
	.datae(!dgrb_ctrl_ac_nt_good),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~49 .extended_lut = "off";
defparam \state~49 .lut_mask = 64'h0035003000350030;
defparam \state~49 .shared_arith = "off";

dffeas \state.s_poa (
	.clk(clk),
	.d(\state~49_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_poa~q ),
	.prn(vcc));
defparam \state.s_poa .is_wysiwyg = "true";
defparam \state.s_poa .power_up = "low";

dffeas \last_state.s_poa (
	.clk(clk),
	.d(\state.s_poa~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\last_state.s_poa~q ),
	.prn(vcc));
defparam \last_state.s_poa .is_wysiwyg = "true";
defparam \last_state.s_poa .power_up = "low";

arriaii_lcell_comb \state~51 (
	.dataa(!\state.s_poa~q ),
	.datab(!\state.s_tracking_setup~q ),
	.datac(!\state~29_combout ),
	.datad(!\process_10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~51 .extended_lut = "off";
defparam \state~51 .lut_mask = 64'h0035003500350035;
defparam \state~51 .shared_arith = "off";

dffeas \state.s_tracking_setup (
	.clk(clk),
	.d(\state~51_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_tracking_setup~q ),
	.prn(vcc));
defparam \state.s_tracking_setup .is_wysiwyg = "true";
defparam \state.s_tracking_setup .power_up = "low";

dffeas \last_state.s_tracking_setup (
	.clk(clk),
	.d(\state.s_tracking_setup~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\last_state.s_tracking_setup~q ),
	.prn(vcc));
defparam \last_state.s_tracking_setup .is_wysiwyg = "true";
defparam \last_state.s_tracking_setup .power_up = "low";

arriaii_lcell_comb \WideNor1~6 (
	.dataa(!\last_state.s_prep_customer_mr_setup~q ),
	.datab(!states_prep_customer_mr_setup),
	.datac(!\last_state.s_tracking_setup~q ),
	.datad(!\state.s_tracking_setup~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor1~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor1~6 .extended_lut = "off";
defparam \WideNor1~6 .lut_mask = 64'h9009900990099009;
defparam \WideNor1~6 .shared_arith = "off";

arriaii_lcell_comb \WideNor1~7 (
	.dataa(!\WideNor1~4_combout ),
	.datab(!\WideNor1~5_combout ),
	.datac(!\last_state.s_poa~q ),
	.datad(!\state.s_poa~q ),
	.datae(!\WideNor1~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor1~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor1~7 .extended_lut = "off";
defparam \WideNor1~7 .lut_mask = 64'h0000100100001001;
defparam \WideNor1~7 .shared_arith = "off";

arriaii_lcell_comb \state~38 (
	.dataa(!\state.s_write_btp~q ),
	.datab(!\state.s_write_mtp~q ),
	.datac(!\state~29_combout ),
	.datad(!\process_10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~38 .extended_lut = "off";
defparam \state~38 .lut_mask = 64'h0035003500350035;
defparam \state~38 .shared_arith = "off";

dffeas \state.s_write_mtp (
	.clk(clk),
	.d(\state~38_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_write_mtp~q ),
	.prn(vcc));
defparam \state.s_write_mtp .is_wysiwyg = "true";
defparam \state.s_write_mtp .power_up = "low";

arriaii_lcell_comb \Selector34~0 (
	.dataa(!\state.s_read_mtp~q ),
	.datab(!\mtp_almts_checked[1]~q ),
	.datac(!\mtp_almts_checked[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector34~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector34~0 .extended_lut = "off";
defparam \Selector34~0 .lut_mask = 64'h1414141414141414;
defparam \Selector34~0 .shared_arith = "off";

dffeas \state.s_reset (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state~31_combout ),
	.q(\state.s_reset~q ),
	.prn(vcc));
defparam \state.s_reset .is_wysiwyg = "true";
defparam \state.s_reset .power_up = "low";

arriaii_lcell_comb \state~37 (
	.dataa(!\state.s_prog_cal_mr~q ),
	.datab(!\state.s_cal~q ),
	.datac(!\state~29_combout ),
	.datad(!\process_10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~37 .extended_lut = "off";
defparam \state~37 .lut_mask = 64'h0035003500350035;
defparam \state~37 .shared_arith = "off";

dffeas \state.s_cal (
	.clk(clk),
	.d(\state~37_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_cal~q ),
	.prn(vcc));
defparam \state.s_cal .is_wysiwyg = "true";
defparam \state.s_cal .power_up = "low";

arriaii_lcell_comb \Selector36~0 (
	.dataa(!\state.s_reset~q ),
	.datab(!\state.s_cal~q ),
	.datac(!states_adv_wr_lat),
	.datad(!\ac_nt_almts_checked~q ),
	.datae(!dgrb_ctrl_ac_nt_good),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector36~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector36~0 .extended_lut = "off";
defparam \Selector36~0 .lut_mask = 64'h004F0F4F004F0F4F;
defparam \Selector36~0 .shared_arith = "off";

dffeas ac_nt_almts_checked(
	.clk(clk),
	.d(\Selector36~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state~29_combout ),
	.q(\ac_nt_almts_checked~q ),
	.prn(vcc));
defparam ac_nt_almts_checked.is_wysiwyg = "true";
defparam ac_nt_almts_checked.power_up = "low";

arriaii_lcell_comb \mtp_almts_checked[1]~0 (
	.dataa(!\state.s_cal~q ),
	.datab(!\state.s_reset~q ),
	.datac(!dgrb_ctrl_ac_nt_good),
	.datad(!\ac_nt_almts_checked~q ),
	.datae(!states_adv_wr_lat),
	.dataf(!\state~29_combout ),
	.datag(!\state.s_read_mtp~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mtp_almts_checked[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mtp_almts_checked[1]~0 .extended_lut = "on";
defparam \mtp_almts_checked[1]~0 .lut_mask = 64'h00000000DFDF0F00;
defparam \mtp_almts_checked[1]~0 .shared_arith = "off";

dffeas \mtp_almts_checked[1] (
	.clk(clk),
	.d(\Selector34~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtp_almts_checked[1]~0_combout ),
	.q(\mtp_almts_checked[1]~q ),
	.prn(vcc));
defparam \mtp_almts_checked[1] .is_wysiwyg = "true";
defparam \mtp_almts_checked[1] .power_up = "low";

arriaii_lcell_comb \mtp_almt:dvw_size_a0[0]~0 (
	.dataa(!\state.s_read_mtp~q ),
	.datab(!\mtp_almts_checked[1]~q ),
	.datac(!\mtp_almts_checked[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mtp_almt:dvw_size_a0[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mtp_almt:dvw_size_a0[0]~0 .extended_lut = "off";
defparam \mtp_almt:dvw_size_a0[0]~0 .lut_mask = 64'h4040404040404040;
defparam \mtp_almt:dvw_size_a0[0]~0 .shared_arith = "off";

dffeas \mtp_almts_checked[0] (
	.clk(clk),
	.d(\mtp_almt:dvw_size_a0[0]~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtp_almts_checked[1]~0_combout ),
	.q(\mtp_almts_checked[0]~q ),
	.prn(vcc));
defparam \mtp_almts_checked[0] .is_wysiwyg = "true";
defparam \mtp_almts_checked[0] .power_up = "low";

arriaii_lcell_comb \state~41 (
	.dataa(!\mtp_almts_checked[1]~q ),
	.datab(!\mtp_almts_checked[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~41 .extended_lut = "off";
defparam \state~41 .lut_mask = 64'h4444444444444444;
defparam \state~41 .shared_arith = "off";

arriaii_lcell_comb \state~42 (
	.dataa(!states_rrp_sweep),
	.datab(!\state.s_read_mtp~q ),
	.datac(!\state~29_combout ),
	.datad(!\process_10~0_combout ),
	.datae(!\state~41_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~42 .extended_lut = "off";
defparam \state~42 .lut_mask = 64'h0035003000350030;
defparam \state~42 .shared_arith = "off";

dffeas \state.s_read_mtp (
	.clk(clk),
	.d(\state~42_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_read_mtp~q ),
	.prn(vcc));
defparam \state.s_read_mtp .is_wysiwyg = "true";
defparam \state.s_read_mtp .power_up = "low";

arriaii_lcell_comb \state~39 (
	.dataa(!\state.s_write_mtp~q ),
	.datab(!\state.s_read_mtp~q ),
	.datac(!states_adv_wr_lat),
	.datad(!\ac_nt_almts_checked~q ),
	.datae(!dgrb_ctrl_ac_nt_good),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~39 .extended_lut = "off";
defparam \state~39 .lut_mask = 64'h8888808888888088;
defparam \state~39 .shared_arith = "off";

arriaii_lcell_comb \state~40 (
	.dataa(!\state.s_rrp_reset~q ),
	.datab(!\state~29_combout ),
	.datac(!\process_10~0_combout ),
	.datad(!\state~39_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~40 .extended_lut = "off";
defparam \state~40 .lut_mask = 64'h0704070407040704;
defparam \state~40 .shared_arith = "off";

dffeas \state.s_rrp_reset (
	.clk(clk),
	.d(\state~40_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_rrp_reset~q ),
	.prn(vcc));
defparam \state.s_rrp_reset .is_wysiwyg = "true";
defparam \state.s_rrp_reset .power_up = "low";

dffeas \last_state.s_rrp_reset (
	.clk(clk),
	.d(\state.s_rrp_reset~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\last_state.s_rrp_reset~q ),
	.prn(vcc));
defparam \last_state.s_rrp_reset .is_wysiwyg = "true";
defparam \last_state.s_rrp_reset .power_up = "low";

dffeas \last_state.s_read_mtp (
	.clk(clk),
	.d(\state.s_read_mtp~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\last_state.s_read_mtp~q ),
	.prn(vcc));
defparam \last_state.s_read_mtp .is_wysiwyg = "true";
defparam \last_state.s_read_mtp .power_up = "low";

arriaii_lcell_comb \WideNor1~2 (
	.dataa(!\last_state.s_write_mtp~q ),
	.datab(!\state.s_write_mtp~q ),
	.datac(!\last_state.s_rrp_reset~q ),
	.datad(!\state.s_rrp_reset~q ),
	.datae(!\last_state.s_read_mtp~q ),
	.dataf(!\state.s_read_mtp~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor1~2 .extended_lut = "off";
defparam \WideNor1~2 .lut_mask = 64'h9009000000009009;
defparam \WideNor1~2 .shared_arith = "off";

dffeas \last_state.s_rrp_sweep (
	.clk(clk),
	.d(states_rrp_sweep),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\last_state.s_rrp_sweep~q ),
	.prn(vcc));
defparam \last_state.s_rrp_sweep .is_wysiwyg = "true";
defparam \last_state.s_rrp_sweep .power_up = "low";

dffeas \last_state.s_rdv (
	.clk(clk),
	.d(states_rdv),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\last_state.s_rdv~q ),
	.prn(vcc));
defparam \last_state.s_rdv .is_wysiwyg = "true";
defparam \last_state.s_rdv .power_up = "low";

dffeas \last_state.s_rrp_seek (
	.clk(clk),
	.d(states_rrp_seek),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\last_state.s_rrp_seek~q ),
	.prn(vcc));
defparam \last_state.s_rrp_seek .is_wysiwyg = "true";
defparam \last_state.s_rrp_seek .power_up = "low";

arriaii_lcell_comb \WideNor1~3 (
	.dataa(!states_rrp_sweep),
	.datab(!\last_state.s_rrp_sweep~q ),
	.datac(!\last_state.s_rdv~q ),
	.datad(!states_rdv),
	.datae(!\last_state.s_rrp_seek~q ),
	.dataf(!states_rrp_seek),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor1~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor1~3 .extended_lut = "off";
defparam \WideNor1~3 .lut_mask = 64'h9009000000009009;
defparam \WideNor1~3 .shared_arith = "off";

arriaii_lcell_comb \timeout_counter_enable~1 (
	.dataa(!\WideNor1~0_combout ),
	.datab(!\WideNor1~1_combout ),
	.datac(!\WideNor1~2_combout ),
	.datad(!\WideNor1~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\timeout_counter_enable~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \timeout_counter_enable~1 .extended_lut = "off";
defparam \timeout_counter_enable~1 .lut_mask = 64'h0001000100010001;
defparam \timeout_counter_enable~1 .shared_arith = "off";

arriaii_lcell_comb \timeout_counter_enable~2 (
	.dataa(!\state.s_non_operational~q ),
	.datab(!\curr_ctrl.command_done~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\timeout_counter_enable~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \timeout_counter_enable~2 .extended_lut = "off";
defparam \timeout_counter_enable~2 .lut_mask = 64'h8888888888888888;
defparam \timeout_counter_enable~2 .shared_arith = "off";

arriaii_lcell_comb \timeout_counter_enable~0 (
	.dataa(!\state.s_reset~q ),
	.datab(!\state.s_operational~q ),
	.datac(!Selector61),
	.datad(!\WideNor1~7_combout ),
	.datae(!\timeout_counter_enable~1_combout ),
	.dataf(!\timeout_counter_enable~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\timeout_counter_enable~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \timeout_counter_enable~0 .extended_lut = "off";
defparam \timeout_counter_enable~0 .lut_mask = 64'hFFFFFFFFBFBFBFBB;
defparam \timeout_counter_enable~0 .shared_arith = "off";

dffeas timeout_counter_clear(
	.clk(clk),
	.d(\timeout_counter_clear~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\timeout_counter_enable~0_combout ),
	.q(\timeout_counter_clear~q ),
	.prn(vcc));
defparam timeout_counter_clear.is_wysiwyg = "true";
defparam timeout_counter_clear.power_up = "low";

dffeas timeout_counter_enable(
	.clk(clk),
	.d(Selector611),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\timeout_counter_enable~0_combout ),
	.q(\timeout_counter_enable~q ),
	.prn(vcc));
defparam timeout_counter_enable.is_wysiwyg = "true";
defparam timeout_counter_enable.power_up = "low";

arriaii_lcell_comb \Add1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\timeout_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h000000000000FF00;
defparam \Add1~13 .shared_arith = "off";

arriaii_lcell_comb \Add1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\timeout_counter[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h000000000000FF00;
defparam \Add1~17 .shared_arith = "off";

arriaii_lcell_comb \timeout_counter~11 (
	.dataa(!\timeout_counter_clear~q ),
	.datab(!\Add1~17_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\timeout_counter~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \timeout_counter~11 .extended_lut = "off";
defparam \timeout_counter~11 .lut_mask = 64'h8888888888888888;
defparam \timeout_counter~11 .shared_arith = "off";

dffeas \timeout_counter[4] (
	.clk(clk),
	.d(\timeout_counter~11_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\timeout_counter[14]~1_combout ),
	.q(\timeout_counter[4]~q ),
	.prn(vcc));
defparam \timeout_counter[4] .is_wysiwyg = "true";
defparam \timeout_counter[4] .power_up = "low";

arriaii_lcell_comb \Add1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\timeout_counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~21_sumout ),
	.cout(\Add1~22 ),
	.shareout());
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h000000000000FF00;
defparam \Add1~21 .shared_arith = "off";

arriaii_lcell_comb \timeout_counter~12 (
	.dataa(!\timeout_counter_clear~q ),
	.datab(!\Add1~21_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\timeout_counter~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \timeout_counter~12 .extended_lut = "off";
defparam \timeout_counter~12 .lut_mask = 64'h8888888888888888;
defparam \timeout_counter~12 .shared_arith = "off";

dffeas \timeout_counter[5] (
	.clk(clk),
	.d(\timeout_counter~12_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\timeout_counter[14]~1_combout ),
	.q(\timeout_counter[5]~q ),
	.prn(vcc));
defparam \timeout_counter[5] .is_wysiwyg = "true";
defparam \timeout_counter[5] .power_up = "low";

arriaii_lcell_comb \Add1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\timeout_counter[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~25_sumout ),
	.cout(\Add1~26 ),
	.shareout());
defparam \Add1~25 .extended_lut = "off";
defparam \Add1~25 .lut_mask = 64'h000000000000FF00;
defparam \Add1~25 .shared_arith = "off";

arriaii_lcell_comb \timeout_counter~13 (
	.dataa(!\timeout_counter_clear~q ),
	.datab(!\Add1~25_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\timeout_counter~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \timeout_counter~13 .extended_lut = "off";
defparam \timeout_counter~13 .lut_mask = 64'h8888888888888888;
defparam \timeout_counter~13 .shared_arith = "off";

dffeas \timeout_counter[6] (
	.clk(clk),
	.d(\timeout_counter~13_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\timeout_counter[14]~1_combout ),
	.q(\timeout_counter[6]~q ),
	.prn(vcc));
defparam \timeout_counter[6] .is_wysiwyg = "true";
defparam \timeout_counter[6] .power_up = "low";

arriaii_lcell_comb \Add1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\timeout_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~29_sumout ),
	.cout(\Add1~30 ),
	.shareout());
defparam \Add1~29 .extended_lut = "off";
defparam \Add1~29 .lut_mask = 64'h000000000000FF00;
defparam \Add1~29 .shared_arith = "off";

arriaii_lcell_comb \timeout_counter~15 (
	.dataa(!\timeout_counter_clear~q ),
	.datab(!\Add1~29_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\timeout_counter~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \timeout_counter~15 .extended_lut = "off";
defparam \timeout_counter~15 .lut_mask = 64'h8888888888888888;
defparam \timeout_counter~15 .shared_arith = "off";

dffeas \timeout_counter[7] (
	.clk(clk),
	.d(\timeout_counter~15_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\timeout_counter[14]~1_combout ),
	.q(\timeout_counter[7]~q ),
	.prn(vcc));
defparam \timeout_counter[7] .is_wysiwyg = "true";
defparam \timeout_counter[7] .power_up = "low";

arriaii_lcell_comb \Add1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\timeout_counter[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~33_sumout ),
	.cout(\Add1~34 ),
	.shareout());
defparam \Add1~33 .extended_lut = "off";
defparam \Add1~33 .lut_mask = 64'h000000000000FF00;
defparam \Add1~33 .shared_arith = "off";

arriaii_lcell_comb \timeout_counter~14 (
	.dataa(!\timeout_counter_clear~q ),
	.datab(!\Add1~33_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\timeout_counter~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \timeout_counter~14 .extended_lut = "off";
defparam \timeout_counter~14 .lut_mask = 64'h8888888888888888;
defparam \timeout_counter~14 .shared_arith = "off";

dffeas \timeout_counter[8] (
	.clk(clk),
	.d(\timeout_counter~14_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\timeout_counter[14]~1_combout ),
	.q(\timeout_counter[8]~q ),
	.prn(vcc));
defparam \timeout_counter[8] .is_wysiwyg = "true";
defparam \timeout_counter[8] .power_up = "low";

arriaii_lcell_comb \Equal1~1 (
	.dataa(!\timeout_counter[13]~q ),
	.datab(!\timeout_counter[4]~q ),
	.datac(!\timeout_counter[5]~q ),
	.datad(!\timeout_counter[6]~q ),
	.datae(!\timeout_counter[8]~q ),
	.dataf(!\timeout_counter[7]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~1 .extended_lut = "off";
defparam \Equal1~1 .lut_mask = 64'h0000000000000001;
defparam \Equal1~1 .shared_arith = "off";

arriaii_lcell_comb \Add1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\timeout_counter[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~37_sumout ),
	.cout(\Add1~38 ),
	.shareout());
defparam \Add1~37 .extended_lut = "off";
defparam \Add1~37 .lut_mask = 64'h000000000000FF00;
defparam \Add1~37 .shared_arith = "off";

arriaii_lcell_comb \timeout_counter~4 (
	.dataa(!\timeout_counter_clear~q ),
	.datab(!\Add1~37_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\timeout_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \timeout_counter~4 .extended_lut = "off";
defparam \timeout_counter~4 .lut_mask = 64'h8888888888888888;
defparam \timeout_counter~4 .shared_arith = "off";

dffeas \timeout_counter[9] (
	.clk(clk),
	.d(\timeout_counter~4_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\timeout_counter[14]~1_combout ),
	.q(\timeout_counter[9]~q ),
	.prn(vcc));
defparam \timeout_counter[9] .is_wysiwyg = "true";
defparam \timeout_counter[9] .power_up = "low";

arriaii_lcell_comb \Add1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\timeout_counter[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~41_sumout ),
	.cout(\Add1~42 ),
	.shareout());
defparam \Add1~41 .extended_lut = "off";
defparam \Add1~41 .lut_mask = 64'h000000000000FF00;
defparam \Add1~41 .shared_arith = "off";

arriaii_lcell_comb \timeout_counter~5 (
	.dataa(!\timeout_counter_clear~q ),
	.datab(!\Add1~41_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\timeout_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \timeout_counter~5 .extended_lut = "off";
defparam \timeout_counter~5 .lut_mask = 64'h8888888888888888;
defparam \timeout_counter~5 .shared_arith = "off";

dffeas \timeout_counter[10] (
	.clk(clk),
	.d(\timeout_counter~5_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\timeout_counter[14]~1_combout ),
	.q(\timeout_counter[10]~q ),
	.prn(vcc));
defparam \timeout_counter[10] .is_wysiwyg = "true";
defparam \timeout_counter[10] .power_up = "low";

arriaii_lcell_comb \Add1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\timeout_counter[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~45_sumout ),
	.cout(\Add1~46 ),
	.shareout());
defparam \Add1~45 .extended_lut = "off";
defparam \Add1~45 .lut_mask = 64'h000000000000FF00;
defparam \Add1~45 .shared_arith = "off";

arriaii_lcell_comb \timeout_counter~6 (
	.dataa(!\timeout_counter_clear~q ),
	.datab(!\Add1~45_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\timeout_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \timeout_counter~6 .extended_lut = "off";
defparam \timeout_counter~6 .lut_mask = 64'h8888888888888888;
defparam \timeout_counter~6 .shared_arith = "off";

dffeas \timeout_counter[11] (
	.clk(clk),
	.d(\timeout_counter~6_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\timeout_counter[14]~1_combout ),
	.q(\timeout_counter[11]~q ),
	.prn(vcc));
defparam \timeout_counter[11] .is_wysiwyg = "true";
defparam \timeout_counter[11] .power_up = "low";

arriaii_lcell_comb \Add1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\timeout_counter[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~49_sumout ),
	.cout(\Add1~50 ),
	.shareout());
defparam \Add1~49 .extended_lut = "off";
defparam \Add1~49 .lut_mask = 64'h000000000000FF00;
defparam \Add1~49 .shared_arith = "off";

arriaii_lcell_comb \timeout_counter~7 (
	.dataa(!\timeout_counter_clear~q ),
	.datab(!\Add1~49_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\timeout_counter~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \timeout_counter~7 .extended_lut = "off";
defparam \timeout_counter~7 .lut_mask = 64'h8888888888888888;
defparam \timeout_counter~7 .shared_arith = "off";

dffeas \timeout_counter[12] (
	.clk(clk),
	.d(\timeout_counter~7_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\timeout_counter[14]~1_combout ),
	.q(\timeout_counter[12]~q ),
	.prn(vcc));
defparam \timeout_counter[12] .is_wysiwyg = "true";
defparam \timeout_counter[12] .power_up = "low";

arriaii_lcell_comb \Add1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\timeout_counter[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~53_sumout ),
	.cout(\Add1~54 ),
	.shareout());
defparam \Add1~53 .extended_lut = "off";
defparam \Add1~53 .lut_mask = 64'h000000000000FF00;
defparam \Add1~53 .shared_arith = "off";

arriaii_lcell_comb \timeout_counter~9 (
	.dataa(!\timeout_counter_clear~q ),
	.datab(!\Add1~53_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\timeout_counter~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \timeout_counter~9 .extended_lut = "off";
defparam \timeout_counter~9 .lut_mask = 64'h8888888888888888;
defparam \timeout_counter~9 .shared_arith = "off";

dffeas \timeout_counter[13] (
	.clk(clk),
	.d(\timeout_counter~9_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\timeout_counter[14]~1_combout ),
	.q(\timeout_counter[13]~q ),
	.prn(vcc));
defparam \timeout_counter[13] .is_wysiwyg = "true";
defparam \timeout_counter[13] .power_up = "low";

arriaii_lcell_comb \Add1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\timeout_counter[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~57_sumout ),
	.cout(),
	.shareout());
defparam \Add1~57 .extended_lut = "off";
defparam \Add1~57 .lut_mask = 64'h000000000000FF00;
defparam \Add1~57 .shared_arith = "off";

arriaii_lcell_comb \timeout_counter~8 (
	.dataa(!\timeout_counter_clear~q ),
	.datab(!\Add1~57_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\timeout_counter~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \timeout_counter~8 .extended_lut = "off";
defparam \timeout_counter~8 .lut_mask = 64'h8888888888888888;
defparam \timeout_counter~8 .shared_arith = "off";

dffeas \timeout_counter[14] (
	.clk(clk),
	.d(\timeout_counter~8_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\timeout_counter[14]~1_combout ),
	.q(\timeout_counter[14]~q ),
	.prn(vcc));
defparam \timeout_counter[14] .is_wysiwyg = "true";
defparam \timeout_counter[14] .power_up = "low";

arriaii_lcell_comb \Equal1~2 (
	.dataa(!\timeout_counter[1]~q ),
	.datab(!\timeout_counter[10]~q ),
	.datac(!\timeout_counter[11]~q ),
	.datad(!\timeout_counter[12]~q ),
	.datae(!\timeout_counter[14]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~2 .extended_lut = "off";
defparam \Equal1~2 .lut_mask = 64'h0000000100000001;
defparam \Equal1~2 .shared_arith = "off";

arriaii_lcell_comb \timeout_counter[14]~16 (
	.dataa(!\timeout_counter[9]~q ),
	.datab(!\timeout_counter[3]~q ),
	.datac(!\timeout_counter[0]~q ),
	.datad(!\timeout_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\timeout_counter[14]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \timeout_counter[14]~16 .extended_lut = "off";
defparam \timeout_counter[14]~16 .lut_mask = 64'h0001000100010001;
defparam \timeout_counter[14]~16 .shared_arith = "off";

arriaii_lcell_comb \timeout_counter[14]~1 (
	.dataa(!\state.s_init_dram~q ),
	.datab(!\timeout_counter_clear~q ),
	.datac(!\timeout_counter_enable~q ),
	.datad(!\Equal1~1_combout ),
	.datae(!\Equal1~2_combout ),
	.dataf(!\timeout_counter[14]~16_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\timeout_counter[14]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \timeout_counter[14]~1 .extended_lut = "off";
defparam \timeout_counter[14]~1 .lut_mask = 64'h3B3B3B3B3B3B3B33;
defparam \timeout_counter[14]~1 .shared_arith = "off";

dffeas \timeout_counter[0] (
	.clk(clk),
	.d(\timeout_counter~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\timeout_counter[14]~1_combout ),
	.q(\timeout_counter[0]~q ),
	.prn(vcc));
defparam \timeout_counter[0] .is_wysiwyg = "true";
defparam \timeout_counter[0] .power_up = "low";

arriaii_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\timeout_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h000000000000FF00;
defparam \Add1~5 .shared_arith = "off";

arriaii_lcell_comb \timeout_counter~3 (
	.dataa(!\timeout_counter_clear~q ),
	.datab(!\Add1~5_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\timeout_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \timeout_counter~3 .extended_lut = "off";
defparam \timeout_counter~3 .lut_mask = 64'h8888888888888888;
defparam \timeout_counter~3 .shared_arith = "off";

dffeas \timeout_counter[1] (
	.clk(clk),
	.d(\timeout_counter~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\timeout_counter[14]~1_combout ),
	.q(\timeout_counter[1]~q ),
	.prn(vcc));
defparam \timeout_counter[1] .is_wysiwyg = "true";
defparam \timeout_counter[1] .power_up = "low";

arriaii_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\timeout_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h000000000000FF00;
defparam \Add1~9 .shared_arith = "off";

arriaii_lcell_comb \timeout_counter~2 (
	.dataa(!\timeout_counter_clear~q ),
	.datab(!\Add1~9_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\timeout_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \timeout_counter~2 .extended_lut = "off";
defparam \timeout_counter~2 .lut_mask = 64'h8888888888888888;
defparam \timeout_counter~2 .shared_arith = "off";

dffeas \timeout_counter[2] (
	.clk(clk),
	.d(\timeout_counter~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\timeout_counter[14]~1_combout ),
	.q(\timeout_counter[2]~q ),
	.prn(vcc));
defparam \timeout_counter[2] .is_wysiwyg = "true";
defparam \timeout_counter[2] .power_up = "low";

arriaii_lcell_comb \timeout_counter~10 (
	.dataa(!\timeout_counter_clear~q ),
	.datab(!\Add1~13_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\timeout_counter~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \timeout_counter~10 .extended_lut = "off";
defparam \timeout_counter~10 .lut_mask = 64'h8888888888888888;
defparam \timeout_counter~10 .shared_arith = "off";

dffeas \timeout_counter[3] (
	.clk(clk),
	.d(\timeout_counter~10_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\timeout_counter[14]~1_combout ),
	.q(\timeout_counter[3]~q ),
	.prn(vcc));
defparam \timeout_counter[3] .is_wysiwyg = "true";
defparam \timeout_counter[3] .power_up = "low";

arriaii_lcell_comb \Equal1~0 (
	.dataa(!\timeout_counter[9]~q ),
	.datab(!\timeout_counter[3]~q ),
	.datac(!\timeout_counter[0]~q ),
	.datad(!\timeout_counter[2]~q ),
	.datae(!\Equal1~1_combout ),
	.dataf(!\Equal1~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'h0000000000000001;
defparam \Equal1~0 .shared_arith = "off";

arriaii_lcell_comb \Selector0~0 (
	.dataa(!curr_ctrlcommand_ack),
	.datab(!curr_cmdcmd_idle),
	.datac(!WideOr0),
	.datad(!dgrb_ctrlcommand_ack),
	.datae(!dgwb_ctrlcommand_ack),
	.dataf(!admin_ctrlcommand_ack),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'h0001AAAB5051FAFB;
defparam \Selector0~0 .shared_arith = "off";

dffeas \curr_ctrl.command_ack (
	.clk(clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\curr_ctrl.command_ack~q ),
	.prn(vcc));
defparam \curr_ctrl.command_ack .is_wysiwyg = "true";
defparam \curr_ctrl.command_ack .power_up = "low";

arriaii_lcell_comb \waiting_for_ack~0 (
	.dataa(!\WideNor1~combout ),
	.datab(!Selector61),
	.datac(!\waiting_for_ack~q ),
	.datad(!\curr_ctrl.command_ack~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\waiting_for_ack~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \waiting_for_ack~0 .extended_lut = "off";
defparam \waiting_for_ack~0 .lut_mask = 64'h2F222F222F222F22;
defparam \waiting_for_ack~0 .shared_arith = "off";

dffeas waiting_for_ack(
	.clk(clk),
	.d(\waiting_for_ack~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\waiting_for_ack~q ),
	.prn(vcc));
defparam waiting_for_ack.is_wysiwyg = "true";
defparam waiting_for_ack.power_up = "low";

arriaii_lcell_comb \flag_ack_timeout~0 (
	.dataa(!\flag_ack_timeout~q ),
	.datab(!\Equal1~0_combout ),
	.datac(!\waiting_for_ack~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\flag_ack_timeout~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \flag_ack_timeout~0 .extended_lut = "off";
defparam \flag_ack_timeout~0 .lut_mask = 64'h5757575757575757;
defparam \flag_ack_timeout~0 .shared_arith = "off";

dffeas flag_ack_timeout(
	.clk(clk),
	.d(\flag_ack_timeout~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\flag_ack_timeout~q ),
	.prn(vcc));
defparam flag_ack_timeout.is_wysiwyg = "true";
defparam flag_ack_timeout.power_up = "low";

arriaii_lcell_comb \process_10~0 (
	.dataa(!\flag_done_timeout~q ),
	.datab(!\curr_ctrl.command_err~q ),
	.datac(!\flag_ack_timeout~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\process_10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \process_10~0 .extended_lut = "off";
defparam \process_10~0 .lut_mask = 64'h8080808080808080;
defparam \process_10~0 .shared_arith = "off";

arriaii_lcell_comb \state~35 (
	.dataa(!\state.s_init_dram~q ),
	.datab(!\state.s_prog_cal_mr~q ),
	.datac(!\state~29_combout ),
	.datad(!\process_10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~35 .extended_lut = "off";
defparam \state~35 .lut_mask = 64'h0035003500350035;
defparam \state~35 .shared_arith = "off";

dffeas \state.s_prog_cal_mr (
	.clk(clk),
	.d(\state~35_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_prog_cal_mr~q ),
	.prn(vcc));
defparam \state.s_prog_cal_mr .is_wysiwyg = "true";
defparam \state.s_prog_cal_mr .power_up = "low";

arriaii_lcell_comb \state~36 (
	.dataa(!\state.s_write_btp~q ),
	.datab(!\state.s_cal~q ),
	.datac(!\state~29_combout ),
	.datad(!\process_10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~36 .extended_lut = "off";
defparam \state~36 .lut_mask = 64'h0053005300530053;
defparam \state~36 .shared_arith = "off";

dffeas \state.s_write_btp (
	.clk(clk),
	.d(\state~36_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_write_btp~q ),
	.prn(vcc));
defparam \state.s_write_btp .is_wysiwyg = "true";
defparam \state.s_write_btp .power_up = "low";

dffeas \last_state.s_write_btp (
	.clk(clk),
	.d(\state.s_write_btp~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\last_state.s_write_btp~q ),
	.prn(vcc));
defparam \last_state.s_write_btp .is_wysiwyg = "true";
defparam \last_state.s_write_btp .power_up = "low";

dffeas \last_state.s_cal (
	.clk(clk),
	.d(\state.s_cal~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\last_state.s_cal~q ),
	.prn(vcc));
defparam \last_state.s_cal .is_wysiwyg = "true";
defparam \last_state.s_cal .power_up = "low";

arriaii_lcell_comb \WideNor1~1 (
	.dataa(!\last_state.s_prog_cal_mr~q ),
	.datab(!\state.s_prog_cal_mr~q ),
	.datac(!\last_state.s_write_btp~q ),
	.datad(!\state.s_write_btp~q ),
	.datae(!\last_state.s_cal~q ),
	.dataf(!\state.s_cal~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor1~1 .extended_lut = "off";
defparam \WideNor1~1 .lut_mask = 64'h9009000000009009;
defparam \WideNor1~1 .shared_arith = "off";

arriaii_lcell_comb WideNor1(
	.dataa(!\WideNor1~0_combout ),
	.datab(!\WideNor1~1_combout ),
	.datac(!\WideNor1~2_combout ),
	.datad(!\WideNor1~3_combout ),
	.datae(!\WideNor1~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideNor1.extended_lut = "off";
defparam WideNor1.lut_mask = 64'h0000000100000001;
defparam WideNor1.shared_arith = "off";

arriaii_lcell_comb \find_cmd~0 (
	.dataa(!\state.s_reset~q ),
	.datab(!\state.s_operational~q ),
	.datac(!\state.s_non_operational~q ),
	.datad(!\state.s_cal~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\find_cmd~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \find_cmd~0 .extended_lut = "off";
defparam \find_cmd~0 .lut_mask = 64'h4000400040004000;
defparam \find_cmd~0 .shared_arith = "off";

arriaii_lcell_comb \dll_lock_counter[0]~0 (
	.dataa(!\dll_lock_counter[0]~q ),
	.datab(!\Equal0~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dll_lock_counter[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dll_lock_counter[0]~0 .extended_lut = "off";
defparam \dll_lock_counter[0]~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \dll_lock_counter[0]~0 .shared_arith = "off";

dffeas \dll_lock_counter[0] (
	.clk(clk),
	.d(\dll_lock_counter[0]~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dll_lock_counter[0]~q ),
	.prn(vcc));
defparam \dll_lock_counter[0] .is_wysiwyg = "true";
defparam \dll_lock_counter[0] .power_up = "low";

arriaii_lcell_comb \dll_lock_counter[1]~5 (
	.dataa(!\Add0~5_sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dll_lock_counter[1]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dll_lock_counter[1]~5 .extended_lut = "off";
defparam \dll_lock_counter[1]~5 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dll_lock_counter[1]~5 .shared_arith = "off";

dffeas \dll_lock_counter[1] (
	.clk(clk),
	.d(\dll_lock_counter[1]~5_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal0~1_combout ),
	.q(\dll_lock_counter[1]~q ),
	.prn(vcc));
defparam \dll_lock_counter[1] .is_wysiwyg = "true";
defparam \dll_lock_counter[1] .power_up = "low";

arriaii_lcell_comb \dll_lock_counter[3]~6 (
	.dataa(!\Add0~13_sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dll_lock_counter[3]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dll_lock_counter[3]~6 .extended_lut = "off";
defparam \dll_lock_counter[3]~6 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dll_lock_counter[3]~6 .shared_arith = "off";

dffeas \dll_lock_counter[3] (
	.clk(clk),
	.d(\dll_lock_counter[3]~6_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal0~1_combout ),
	.q(\dll_lock_counter[3]~q ),
	.prn(vcc));
defparam \dll_lock_counter[3] .is_wysiwyg = "true";
defparam \dll_lock_counter[3] .power_up = "low";

arriaii_lcell_comb \dll_lock_counter[2]~7 (
	.dataa(!\Add0~9_sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dll_lock_counter[2]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dll_lock_counter[2]~7 .extended_lut = "off";
defparam \dll_lock_counter[2]~7 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dll_lock_counter[2]~7 .shared_arith = "off";

dffeas \dll_lock_counter[2] (
	.clk(clk),
	.d(\dll_lock_counter[2]~7_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal0~1_combout ),
	.q(\dll_lock_counter[2]~q ),
	.prn(vcc));
defparam \dll_lock_counter[2] .is_wysiwyg = "true";
defparam \dll_lock_counter[2] .power_up = "low";

arriaii_lcell_comb \Equal0~1 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\dll_lock_counter[0]~q ),
	.datac(!\dll_lock_counter[1]~q ),
	.datad(!\dll_lock_counter[3]~q ),
	.datae(!\dll_lock_counter[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~1 .extended_lut = "off";
defparam \Equal0~1 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \Equal0~1 .shared_arith = "off";

arriaii_lcell_comb \dis_state~0 (
	.dataa(!\state.s_phy_initialise~q ),
	.datab(!\WideNor1~combout ),
	.datac(!\dis_state~q ),
	.datad(!\find_cmd~0_combout ),
	.datae(!\Equal0~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dis_state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dis_state~0 .extended_lut = "off";
defparam \dis_state~0 .lut_mask = 64'hFF57AA02FF57AA02;
defparam \dis_state~0 .shared_arith = "off";

dffeas dis_state(
	.clk(clk),
	.d(\dis_state~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dis_state~q ),
	.prn(vcc));
defparam dis_state.is_wysiwyg = "true";
defparam dis_state.power_up = "low";

arriaii_lcell_comb \state~29 (
	.dataa(!\hold_state~q ),
	.datab(!\curr_ctrl.command_done~q ),
	.datac(!\dis_state~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~29 .extended_lut = "off";
defparam \state~29 .lut_mask = 64'h2A2A2A2A2A2A2A2A;
defparam \state~29 .shared_arith = "off";

arriaii_lcell_comb \state.s_non_operational~0 (
	.dataa(!\state.s_non_operational~q ),
	.datab(!states_adv_wr_lat),
	.datac(!\state~29_combout ),
	.datad(!\process_10~0_combout ),
	.datae(!\ac_nt_almts_checked~q ),
	.dataf(!dgrb_ctrl_ac_nt_good),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state.s_non_operational~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state.s_non_operational~0 .extended_lut = "off";
defparam \state.s_non_operational~0 .lut_mask = 64'hFF55FF55FF55FF57;
defparam \state.s_non_operational~0 .shared_arith = "off";

dffeas \state.s_non_operational (
	.clk(clk),
	.d(\state.s_non_operational~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.s_non_operational~q ),
	.prn(vcc));
defparam \state.s_non_operational .is_wysiwyg = "true";
defparam \state.s_non_operational .power_up = "low";

arriaii_lcell_comb \Selector40~0 (
	.dataa(!\int_ctl_init_fail~q ),
	.datab(!\state.s_non_operational~q ),
	.datac(!\state.s_tracking~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector40~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector40~0 .extended_lut = "off";
defparam \Selector40~0 .lut_mask = 64'h3737373737373737;
defparam \Selector40~0 .shared_arith = "off";

dffeas int_ctl_init_fail(
	.clk(clk),
	.d(\Selector40~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state~29_combout ),
	.q(\int_ctl_init_fail~q ),
	.prn(vcc));
defparam int_ctl_init_fail.is_wysiwyg = "true";
defparam int_ctl_init_fail.power_up = "low";

arriaii_lcell_comb \Selector39~0 (
	.dataa(!\int_ctl_init_success~q ),
	.datab(!\state.s_operational~q ),
	.datac(!\state.s_tracking~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector39~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector39~0 .extended_lut = "off";
defparam \Selector39~0 .lut_mask = 64'h3737373737373737;
defparam \Selector39~0 .shared_arith = "off";

dffeas int_ctl_init_success(
	.clk(clk),
	.d(\Selector39~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\state~29_combout ),
	.q(\int_ctl_init_success~q ),
	.prn(vcc));
defparam int_ctl_init_success.is_wysiwyg = "true";
defparam int_ctl_init_success.power_up = "low";

arriaii_lcell_comb \state~30 (
	.dataa(!states_rrp_sweep),
	.datab(!\state.s_rrp_reset~q ),
	.datac(!\state~29_combout ),
	.datad(!\process_10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~30 .extended_lut = "off";
defparam \state~30 .lut_mask = 64'h0053005300530053;
defparam \state~30 .shared_arith = "off";

arriaii_lcell_comb \state~43 (
	.dataa(!states_rdv),
	.datab(!states_rrp_seek),
	.datac(!\state~29_combout ),
	.datad(!\process_10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~43 .extended_lut = "off";
defparam \state~43 .lut_mask = 64'h0053005300530053;
defparam \state~43 .shared_arith = "off";

arriaii_lcell_comb \state~44 (
	.dataa(!states_rrp_sweep),
	.datab(!states_rrp_seek),
	.datac(!\state~29_combout ),
	.datad(!\process_10~0_combout ),
	.datae(!\state~41_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~44 .extended_lut = "off";
defparam \state~44 .lut_mask = 64'h0030003500300035;
defparam \state~44 .shared_arith = "off";

arriaii_lcell_comb \state~45 (
	.dataa(!states_rdv),
	.datab(!states_was),
	.datac(!\state~29_combout ),
	.datad(!\process_10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~45 .extended_lut = "off";
defparam \state~45 .lut_mask = 64'h0035003500350035;
defparam \state~45 .shared_arith = "off";

arriaii_lcell_comb \state~46 (
	.dataa(!states_adv_wr_lat),
	.datab(!states_adv_rd_lat),
	.datac(!\state~29_combout ),
	.datad(!\process_10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~46 .extended_lut = "off";
defparam \state~46 .lut_mask = 64'h0053005300530053;
defparam \state~46 .shared_arith = "off";

arriaii_lcell_comb \state~47 (
	.dataa(!states_was),
	.datab(!states_adv_rd_lat),
	.datac(!\state~29_combout ),
	.datad(!\process_10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~47 .extended_lut = "off";
defparam \state~47 .lut_mask = 64'h0035003500350035;
defparam \state~47 .shared_arith = "off";

arriaii_lcell_comb \state~50 (
	.dataa(!states_prep_customer_mr_setup),
	.datab(!\state.s_tracking_setup~q ),
	.datac(!\state~29_combout ),
	.datad(!\process_10~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~50_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~50 .extended_lut = "off";
defparam \state~50 .lut_mask = 64'h0053005300530053;
defparam \state~50 .shared_arith = "off";

arriaii_lcell_comb \Selector33~0 (
	.dataa(!\state.s_reset~q ),
	.datab(!states_adv_wr_lat),
	.datac(!ac_nt_0),
	.datad(!\ac_nt_almts_checked~q ),
	.datae(!dgrb_ctrl_ac_nt_good),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector33~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector33~0 .extended_lut = "off";
defparam \Selector33~0 .lut_mask = 64'h0707340707073407;
defparam \Selector33~0 .shared_arith = "off";

arriaii_lcell_comb \master_ctrl_op_rec~1 (
	.dataa(!states_was),
	.datab(!master_ctrl_op_rec),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_ctrl_op_rec~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_ctrl_op_rec~1 .extended_lut = "off";
defparam \master_ctrl_op_rec~1 .lut_mask = 64'h4444444444444444;
defparam \master_ctrl_op_rec~1 .shared_arith = "off";

arriaii_lcell_comb \master_ctrl_op_rec~2 (
	.dataa(!\state.s_write_btp~q ),
	.datab(!master_ctrl_op_rec),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_ctrl_op_rec~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_ctrl_op_rec~2 .extended_lut = "off";
defparam \master_ctrl_op_rec~2 .lut_mask = 64'h4444444444444444;
defparam \master_ctrl_op_rec~2 .shared_arith = "off";

arriaii_lcell_comb \master_ctrl_op_rec~3 (
	.dataa(!\state.s_write_mtp~q ),
	.datab(!master_ctrl_op_rec),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_ctrl_op_rec~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_ctrl_op_rec~3 .extended_lut = "off";
defparam \master_ctrl_op_rec~3 .lut_mask = 64'h4444444444444444;
defparam \master_ctrl_op_rec~3 .shared_arith = "off";

arriaii_lcell_comb \master_ctrl_op_rec~4 (
	.dataa(!states_prep_customer_mr_setup),
	.datab(!master_ctrl_op_rec),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_ctrl_op_rec~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_ctrl_op_rec~4 .extended_lut = "off";
defparam \master_ctrl_op_rec~4 .lut_mask = 64'h4444444444444444;
defparam \master_ctrl_op_rec~4 .shared_arith = "off";

arriaii_lcell_comb \master_ctrl_op_rec~5 (
	.dataa(!\state.s_init_dram~q ),
	.datab(!master_ctrl_op_rec),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_ctrl_op_rec~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_ctrl_op_rec~5 .extended_lut = "off";
defparam \master_ctrl_op_rec~5 .lut_mask = 64'h4444444444444444;
defparam \master_ctrl_op_rec~5 .shared_arith = "off";

arriaii_lcell_comb \master_ctrl_op_rec~6 (
	.dataa(!\state.s_prog_cal_mr~q ),
	.datab(!master_ctrl_op_rec),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\master_ctrl_op_rec~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \master_ctrl_op_rec~6 .extended_lut = "off";
defparam \master_ctrl_op_rec~6 .lut_mask = 64'h4444444444444444;
defparam \master_ctrl_op_rec~6 .shared_arith = "off";

dffeas \last_state.s_reset (
	.clk(clk),
	.d(\state.s_reset~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\last_state.s_reset~q ),
	.prn(vcc));
defparam \last_state.s_reset .is_wysiwyg = "true";
defparam \last_state.s_reset .power_up = "low";

dffeas \last_state.s_init_dram (
	.clk(clk),
	.d(\state.s_init_dram~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\last_state.s_init_dram~q ),
	.prn(vcc));
defparam \last_state.s_init_dram .is_wysiwyg = "true";
defparam \last_state.s_init_dram .power_up = "low";

dffeas \last_state.s_phy_initialise (
	.clk(clk),
	.d(\state.s_phy_initialise~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\last_state.s_phy_initialise~q ),
	.prn(vcc));
defparam \last_state.s_phy_initialise .is_wysiwyg = "true";
defparam \last_state.s_phy_initialise .power_up = "low";

arriaii_lcell_comb \WideNor1~0 (
	.dataa(!\state.s_reset~q ),
	.datab(!\last_state.s_reset~q ),
	.datac(!\last_state.s_init_dram~q ),
	.datad(!\state.s_init_dram~q ),
	.datae(!\last_state.s_phy_initialise~q ),
	.dataf(!\state.s_phy_initialise~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor1~0 .extended_lut = "off";
defparam \WideNor1~0 .lut_mask = 64'h9009000000009009;
defparam \WideNor1~0 .shared_arith = "off";

arriaii_lcell_comb \WideNor2~0 (
	.dataa(!\state.s_reset~q ),
	.datab(!\state.s_phy_initialise~q ),
	.datac(!\state.s_cal~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideNor2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideNor2~0 .extended_lut = "off";
defparam \WideNor2~0 .lut_mask = 64'h4040404040404040;
defparam \WideNor2~0 .shared_arith = "off";

arriaii_lcell_comb \Selector4~0 (
	.dataa(!curr_ctrlcommand_ack),
	.datab(!curr_cmdcmd_idle),
	.datac(!WideOr0),
	.datad(!dgrb_ctrlcommand_result_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~0 .extended_lut = "off";
defparam \Selector4~0 .lut_mask = 64'h0001000100010001;
defparam \Selector4~0 .shared_arith = "off";

dffeas \curr_ctrl.command_result[5] (
	.clk(clk),
	.d(\Selector4~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\curr_ctrl.command_result[5]~q ),
	.prn(vcc));
defparam \curr_ctrl.command_result[5] .is_wysiwyg = "true";
defparam \curr_ctrl.command_result[5] .power_up = "low";

arriaii_lcell_comb \mtp_almt:dvw_size_a1[0]~0 (
	.dataa(!\state.s_read_mtp~q ),
	.datab(!\curr_ctrl.command_done~q ),
	.datac(!\mtp_almts_checked[1]~q ),
	.datad(!\mtp_almts_checked[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mtp_almt:dvw_size_a1[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mtp_almt:dvw_size_a1[0]~0 .extended_lut = "off";
defparam \mtp_almt:dvw_size_a1[0]~0 .lut_mask = 64'h0111011101110111;
defparam \mtp_almt:dvw_size_a1[0]~0 .shared_arith = "off";

dffeas \mtp_almt:dvw_size_a1[5] (
	.clk(clk),
	.d(\curr_ctrl.command_result[5]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtp_almt:dvw_size_a1[0]~0_combout ),
	.q(\mtp_almt:dvw_size_a1[5]~q ),
	.prn(vcc));
defparam \mtp_almt:dvw_size_a1[5] .is_wysiwyg = "true";
defparam \mtp_almt:dvw_size_a1[5] .power_up = "low";

arriaii_lcell_comb \Selector6~0 (
	.dataa(!curr_ctrlcommand_ack),
	.datab(!curr_cmdcmd_idle),
	.datac(!WideOr0),
	.datad(!dgrb_ctrlcommand_result_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~0 .extended_lut = "off";
defparam \Selector6~0 .lut_mask = 64'h0001000100010001;
defparam \Selector6~0 .shared_arith = "off";

dffeas \curr_ctrl.command_result[3] (
	.clk(clk),
	.d(\Selector6~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\curr_ctrl.command_result[3]~q ),
	.prn(vcc));
defparam \curr_ctrl.command_result[3] .is_wysiwyg = "true";
defparam \curr_ctrl.command_result[3] .power_up = "low";

arriaii_lcell_comb \mtp_almt:dvw_size_a0[0]~1 (
	.dataa(!\state.s_read_mtp~q ),
	.datab(!\curr_ctrl.command_done~q ),
	.datac(!\mtp_almts_checked[1]~q ),
	.datad(!\mtp_almts_checked[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mtp_almt:dvw_size_a0[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mtp_almt:dvw_size_a0[0]~1 .extended_lut = "off";
defparam \mtp_almt:dvw_size_a0[0]~1 .lut_mask = 64'h1000100010001000;
defparam \mtp_almt:dvw_size_a0[0]~1 .shared_arith = "off";

dffeas \mtp_almt:dvw_size_a0[3] (
	.clk(clk),
	.d(\curr_ctrl.command_result[3]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtp_almt:dvw_size_a0[0]~1_combout ),
	.q(\mtp_almt:dvw_size_a0[3]~q ),
	.prn(vcc));
defparam \mtp_almt:dvw_size_a0[3] .is_wysiwyg = "true";
defparam \mtp_almt:dvw_size_a0[3] .power_up = "low";

dffeas \mtp_almt:dvw_size_a1[3] (
	.clk(clk),
	.d(\curr_ctrl.command_result[3]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtp_almt:dvw_size_a1[0]~0_combout ),
	.q(\mtp_almt:dvw_size_a1[3]~q ),
	.prn(vcc));
defparam \mtp_almt:dvw_size_a1[3] .is_wysiwyg = "true";
defparam \mtp_almt:dvw_size_a1[3] .power_up = "low";

arriaii_lcell_comb \Selector5~0 (
	.dataa(!curr_ctrlcommand_ack),
	.datab(!curr_cmdcmd_idle),
	.datac(!WideOr0),
	.datad(!dgrb_ctrlcommand_result_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~0 .extended_lut = "off";
defparam \Selector5~0 .lut_mask = 64'h0001000100010001;
defparam \Selector5~0 .shared_arith = "off";

dffeas \curr_ctrl.command_result[4] (
	.clk(clk),
	.d(\Selector5~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\curr_ctrl.command_result[4]~q ),
	.prn(vcc));
defparam \curr_ctrl.command_result[4] .is_wysiwyg = "true";
defparam \curr_ctrl.command_result[4] .power_up = "low";

dffeas \mtp_almt:dvw_size_a0[4] (
	.clk(clk),
	.d(\curr_ctrl.command_result[4]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtp_almt:dvw_size_a0[0]~1_combout ),
	.q(\mtp_almt:dvw_size_a0[4]~q ),
	.prn(vcc));
defparam \mtp_almt:dvw_size_a0[4] .is_wysiwyg = "true";
defparam \mtp_almt:dvw_size_a0[4] .power_up = "low";

dffeas \mtp_almt:dvw_size_a1[4] (
	.clk(clk),
	.d(\curr_ctrl.command_result[4]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mtp_almt:dvw_size_a1[0]~0_combout ),
	.q(\mtp_almt:dvw_size_a1[4]~q ),
	.prn(vcc));
defparam \mtp_almt:dvw_size_a1[4] .is_wysiwyg = "true";
defparam \mtp_almt:dvw_size_a1[4] .power_up = "low";

arriaii_lcell_comb \LessThan0~1 (
	.dataa(!\LessThan0~0_combout ),
	.datab(!\mtp_almt:dvw_size_a0[3]~q ),
	.datac(!\mtp_almt:dvw_size_a1[3]~q ),
	.datad(!\mtp_almt:dvw_size_a0[4]~q ),
	.datae(!\mtp_almt:dvw_size_a1[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~1 .extended_lut = "off";
defparam \LessThan0~1 .lut_mask = 64'h4D00FF4D4D00FF4D;
defparam \LessThan0~1 .shared_arith = "off";

arriaii_lcell_comb \LessThan0~2 (
	.dataa(!\mtp_almt:dvw_size_a0[5]~q ),
	.datab(!\mtp_almt:dvw_size_a1[5]~q ),
	.datac(!\LessThan0~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~2 .extended_lut = "off";
defparam \LessThan0~2 .lut_mask = 64'h2B2B2B2B2B2B2B2B;
defparam \LessThan0~2 .shared_arith = "off";

dffeas mtp_correct_almt(
	.clk(clk),
	.d(\LessThan0~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mtp_correct_almt~q ),
	.prn(vcc));
defparam mtp_correct_almt.is_wysiwyg = "true";
defparam mtp_correct_almt.power_up = "low";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_dgrb (
	q_b_0,
	q_b_64,
	q_b_1,
	q_b_65,
	q_b_2,
	q_b_66,
	q_b_3,
	q_b_67,
	q_b_4,
	q_b_68,
	q_b_5,
	q_b_69,
	q_b_6,
	q_b_70,
	q_b_7,
	q_b_71,
	q_b_16,
	q_b_80,
	q_b_17,
	q_b_81,
	q_b_18,
	q_b_82,
	q_b_19,
	q_b_83,
	q_b_20,
	q_b_84,
	q_b_21,
	q_b_85,
	q_b_22,
	q_b_86,
	q_b_23,
	q_b_87,
	q_b_32,
	q_b_96,
	q_b_33,
	q_b_97,
	q_b_34,
	q_b_98,
	q_b_35,
	q_b_99,
	q_b_36,
	q_b_100,
	q_b_37,
	q_b_101,
	q_b_38,
	q_b_102,
	q_b_39,
	q_b_103,
	q_b_48,
	q_b_112,
	q_b_49,
	q_b_113,
	q_b_50,
	q_b_114,
	q_b_51,
	q_b_115,
	q_b_52,
	q_b_116,
	q_b_53,
	q_b_117,
	q_b_54,
	q_b_118,
	q_b_55,
	q_b_119,
	q_b_8,
	q_b_72,
	q_b_9,
	q_b_73,
	q_b_10,
	q_b_74,
	q_b_11,
	q_b_75,
	q_b_12,
	q_b_76,
	q_b_13,
	q_b_77,
	q_b_14,
	q_b_78,
	q_b_15,
	q_b_79,
	q_b_24,
	q_b_88,
	q_b_25,
	q_b_89,
	q_b_26,
	q_b_90,
	q_b_27,
	q_b_91,
	q_b_28,
	q_b_92,
	q_b_29,
	q_b_93,
	q_b_30,
	q_b_94,
	q_b_31,
	q_b_95,
	q_b_40,
	q_b_104,
	q_b_41,
	q_b_105,
	q_b_42,
	q_b_106,
	q_b_43,
	q_b_107,
	q_b_44,
	q_b_108,
	q_b_45,
	q_b_109,
	q_b_46,
	q_b_110,
	q_b_47,
	q_b_111,
	q_b_56,
	q_b_120,
	q_b_57,
	q_b_121,
	q_b_58,
	q_b_122,
	q_b_59,
	q_b_123,
	q_b_60,
	q_b_124,
	q_b_61,
	q_b_125,
	q_b_62,
	q_b_126,
	q_b_63,
	q_b_127,
	clk,
	rst_n,
	wd_lat_2,
	wd_lat_1,
	wd_lat_0,
	wd_lat_3,
	wd_lat_4,
	sig_doing_rd_0,
	seq_rdata_valid_lat_dec1,
	sig_doing_rd_4,
	dgb_ac_access_gnt_r,
	dgrb_ctrl_ac_nt_good1,
	seq_pll_inc_dec_n1,
	seq_pll_start_reconfig1,
	dgrb_ctrlcommand_done,
	curr_ctrlcommand_ack,
	curr_cmdcmd_idle,
	WideOr0,
	rdata_valid,
	seq_rdata_valid_1,
	dgrb_ctrlcommand_err,
	seq_pll_select_0,
	seq_pll_select_1,
	WideOr2,
	ac_muxctrl_broadcast_rcommand_req,
	sig_addr_cmd0cke0,
	dgrb_ac_access_req1,
	sig_addr_cmd1cs_n0,
	sig_addr_cmd0addr3,
	sig_addr_cmd0addr4,
	sig_addr_cmd0addr5,
	sig_addr_cmd0addr12,
	\ctrl_dgrb.command.cmd_prep_adv_wr_lat ,
	\ctrl_dgrb.command.cmd_rdv ,
	\ctrl_dgrb.command.cmd_read_mtp ,
	dgrb_ctrlcommand_ack,
	\ctrl_dgrb.command.cmd_rrp_seek ,
	\ctrl_dgrb.command.cmd_rrp_reset ,
	\ctrl_dgrb.command.cmd_rrp_sweep ,
	\ctrl_dgrb.command.cmd_tr_due ,
	\ctrl_dgrb.command.cmd_poa ,
	\ctrl_dgrb.command.cmd_prep_adv_rd_lat ,
	phs_shft_busy,
	\ctrl_dgrb.command_op.mtp_almt ,
	mmc_seq_done,
	seq_poa_lat_dec_1x_0,
	\ctrl_dgrb.command_op.single_bit ,
	dgrb_ctrlcommand_result_5,
	dgrb_ctrlcommand_result_2,
	dgrb_ctrlcommand_result_1,
	dgrb_ctrlcommand_result_0,
	dgrb_ctrlcommand_result_3,
	dgrb_ctrlcommand_result_4,
	seq_mmc_start1,
	mmc_seq_value,
	GND_port)/* synthesis synthesis_greybox=0 */;
input 	q_b_0;
input 	q_b_64;
input 	q_b_1;
input 	q_b_65;
input 	q_b_2;
input 	q_b_66;
input 	q_b_3;
input 	q_b_67;
input 	q_b_4;
input 	q_b_68;
input 	q_b_5;
input 	q_b_69;
input 	q_b_6;
input 	q_b_70;
input 	q_b_7;
input 	q_b_71;
input 	q_b_16;
input 	q_b_80;
input 	q_b_17;
input 	q_b_81;
input 	q_b_18;
input 	q_b_82;
input 	q_b_19;
input 	q_b_83;
input 	q_b_20;
input 	q_b_84;
input 	q_b_21;
input 	q_b_85;
input 	q_b_22;
input 	q_b_86;
input 	q_b_23;
input 	q_b_87;
input 	q_b_32;
input 	q_b_96;
input 	q_b_33;
input 	q_b_97;
input 	q_b_34;
input 	q_b_98;
input 	q_b_35;
input 	q_b_99;
input 	q_b_36;
input 	q_b_100;
input 	q_b_37;
input 	q_b_101;
input 	q_b_38;
input 	q_b_102;
input 	q_b_39;
input 	q_b_103;
input 	q_b_48;
input 	q_b_112;
input 	q_b_49;
input 	q_b_113;
input 	q_b_50;
input 	q_b_114;
input 	q_b_51;
input 	q_b_115;
input 	q_b_52;
input 	q_b_116;
input 	q_b_53;
input 	q_b_117;
input 	q_b_54;
input 	q_b_118;
input 	q_b_55;
input 	q_b_119;
input 	q_b_8;
input 	q_b_72;
input 	q_b_9;
input 	q_b_73;
input 	q_b_10;
input 	q_b_74;
input 	q_b_11;
input 	q_b_75;
input 	q_b_12;
input 	q_b_76;
input 	q_b_13;
input 	q_b_77;
input 	q_b_14;
input 	q_b_78;
input 	q_b_15;
input 	q_b_79;
input 	q_b_24;
input 	q_b_88;
input 	q_b_25;
input 	q_b_89;
input 	q_b_26;
input 	q_b_90;
input 	q_b_27;
input 	q_b_91;
input 	q_b_28;
input 	q_b_92;
input 	q_b_29;
input 	q_b_93;
input 	q_b_30;
input 	q_b_94;
input 	q_b_31;
input 	q_b_95;
input 	q_b_40;
input 	q_b_104;
input 	q_b_41;
input 	q_b_105;
input 	q_b_42;
input 	q_b_106;
input 	q_b_43;
input 	q_b_107;
input 	q_b_44;
input 	q_b_108;
input 	q_b_45;
input 	q_b_109;
input 	q_b_46;
input 	q_b_110;
input 	q_b_47;
input 	q_b_111;
input 	q_b_56;
input 	q_b_120;
input 	q_b_57;
input 	q_b_121;
input 	q_b_58;
input 	q_b_122;
input 	q_b_59;
input 	q_b_123;
input 	q_b_60;
input 	q_b_124;
input 	q_b_61;
input 	q_b_125;
input 	q_b_62;
input 	q_b_126;
input 	q_b_63;
input 	q_b_127;
input 	clk;
input 	rst_n;
output 	wd_lat_2;
output 	wd_lat_1;
output 	wd_lat_0;
output 	wd_lat_3;
output 	wd_lat_4;
output 	sig_doing_rd_0;
output 	seq_rdata_valid_lat_dec1;
output 	sig_doing_rd_4;
input 	dgb_ac_access_gnt_r;
output 	dgrb_ctrl_ac_nt_good1;
output 	seq_pll_inc_dec_n1;
output 	seq_pll_start_reconfig1;
output 	dgrb_ctrlcommand_done;
input 	curr_ctrlcommand_ack;
input 	curr_cmdcmd_idle;
input 	WideOr0;
input 	[1:0] rdata_valid;
input 	seq_rdata_valid_1;
output 	dgrb_ctrlcommand_err;
output 	seq_pll_select_0;
output 	seq_pll_select_1;
input 	WideOr2;
input 	ac_muxctrl_broadcast_rcommand_req;
input 	sig_addr_cmd0cke0;
output 	dgrb_ac_access_req1;
output 	sig_addr_cmd1cs_n0;
output 	sig_addr_cmd0addr3;
output 	sig_addr_cmd0addr4;
output 	sig_addr_cmd0addr5;
output 	sig_addr_cmd0addr12;
input 	\ctrl_dgrb.command.cmd_prep_adv_wr_lat ;
input 	\ctrl_dgrb.command.cmd_rdv ;
input 	\ctrl_dgrb.command.cmd_read_mtp ;
output 	dgrb_ctrlcommand_ack;
input 	\ctrl_dgrb.command.cmd_rrp_seek ;
input 	\ctrl_dgrb.command.cmd_rrp_reset ;
input 	\ctrl_dgrb.command.cmd_rrp_sweep ;
input 	\ctrl_dgrb.command.cmd_tr_due ;
input 	\ctrl_dgrb.command.cmd_poa ;
input 	\ctrl_dgrb.command.cmd_prep_adv_rd_lat ;
input 	phs_shft_busy;
input 	\ctrl_dgrb.command_op.mtp_almt ;
input 	mmc_seq_done;
output 	seq_poa_lat_dec_1x_0;
input 	\ctrl_dgrb.command_op.single_bit ;
output 	dgrb_ctrlcommand_result_5;
output 	dgrb_ctrlcommand_result_2;
output 	dgrb_ctrlcommand_result_1;
output 	dgrb_ctrlcommand_result_0;
output 	dgrb_ctrlcommand_result_3;
output 	dgrb_ctrlcommand_result_4;
output 	seq_mmc_start1;
input 	mmc_seq_value;
input 	GND_port;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add24~1_sumout ;
wire \trk_block:sig_trk_state.s_trk_complete~q ;
wire \Add5~3_sumout ;
wire \Add15~5_sumout ;
wire \Add15~9_sumout ;
wire \Add15~13_sumout ;
wire \Add15~17_sumout ;
wire \Add18~21_sumout ;
wire \Add12~1_sumout ;
wire \Add12~13_sumout ;
wire \rsc_block:sig_rewind_direction~q ;
wire \rsc_block:sig_num_phase_shifts[0]~q ;
wire \sig_cmd_err~2_combout ;
wire \sig_rewind_direction~0_combout ;
wire \rsc_block:sig_num_phase_shifts[0]~0_combout ;
wire \sig_trk_state~20_combout ;
wire \sig_trk_state~23_combout ;
wire \sig_cdvw_state.invalid_phase_seen~q ;
wire \Equal15~0_combout ;
wire \tp_match_block:sig_rdata_current_pin[1]~q ;
wire \LessThan3~0_combout ;
wire \v_cdvw_state~7_combout ;
wire \single_bit_cal~q ;
wire \Mux6~1_combout ;
wire \Mux5~1_combout ;
wire \Mux8~1_combout ;
wire \Mux7~1_combout ;
wire \ctrl_dgrb_r.command_op.single_bit~q ;
wire \ac_block:sig_addr_cmd_last_state.s_ac_relax~q ;
wire \ctrl_dgrb_r.command.cmd_rdv~q ;
wire \sig_dgrb_state~47_combout ;
wire \sig_dgrb_state.s_rdata_valid_align~q ;
wire \ctrl_dgrb_r.command.cmd_prep_adv_rd_lat~q ;
wire \sig_dgrb_state~57_combout ;
wire \sig_dgrb_state.s_adv_rd_lat_setup~q ;
wire \v_aligned~0_combout ;
wire \ctrl_dgrb_r.command.cmd_tr_due~q ;
wire \sig_dgrb_state~51_combout ;
wire \sig_dgrb_state.s_track~q ;
wire \Add4~1_sumout ;
wire \ctrl_dgrb_r.command.cmd_read_mtp~q ;
wire \sig_dgrb_state~61_combout ;
wire \sig_dgrb_state.s_read_mtp~q ;
wire \cdvw_block:sig_cdvw_calc_1t~q ;
wire \v_cdvw_state~2_combout ;
wire \sig_dgrb_last_state.s_track~q ;
wire \cdvw_proc~2_combout ;
wire \trk_block:mmc_seq_req_sync:v_mmc_seq_done_1r~q ;
wire \trk_block:mmc_seq_req_sync:v_mmc_seq_done_2r~q ;
wire \trk_block:mmc_seq_req_sync:v_mmc_seq_done_3r~q ;
wire \trk_block:sig_mmc_seq_done_1t~q ;
wire \shift_in_mmc_seq_value~0_combout ;
wire \sig_trk_cdvw_shift_in~q ;
wire \Add7~1_sumout ;
wire \single_bit_cal~_wirecell_combout ;
wire \phs_shft_busy_reg:phs_shft_busy_1r~q ;
wire \phs_shft_busy_reg:phs_shft_busy_2r~q ;
wire \sig_phs_shft_end~0_combout ;
wire \sig_phs_shft_end~q ;
wire \Selector23~0_combout ;
wire \sig_rsc_req.s_rsc_test_phase~q ;
wire \Selector51~0_combout ;
wire \rsc_block:sig_rsc_state.s_rsc_test_phase~q ;
wire \sig_dq_pin_ctr[0]~0_combout ;
wire \rsc_block:sig_rsc_last_state.s_rsc_test_dq~q ;
wire \rsc_block:sig_rsc_last_state.s_rsc_seek_cdvw~q ;
wire \rsc_block:sig_rsc_last_state.s_rsc_cdvw_calc~q ;
wire \Selector58~2_combout ;
wire \rsc_block:sig_rsc_state.s_rsc_cdvw_wait~q ;
wire \Selector59~0_combout ;
wire \rsc_block:sig_rsc_state.s_rsc_seek_cdvw~q ;
wire \rsc_block:sig_count[6]~0_combout ;
wire \Add2~1_sumout ;
wire \cdvw_proc~1_combout ;
wire \Add2~6 ;
wire \Add2~9_sumout ;
wire \Add4~6 ;
wire \Add4~9_sumout ;
wire \sig_cdvw_state.current_bit[5]~0_combout ;
wire \sig_cdvw_state.current_bit[2]~q ;
wire \v_cdvw_state~21_combout ;
wire \sig_cdvw_state.last_bit_value~q ;
wire \find_centre_of_largest_data_valid_window~2_combout ;
wire \v_cdvw_state~6_combout ;
wire \sig_cdvw_state.found_a_good_edge~q ;
wire \v_cdvw_state~22_combout ;
wire \sig_cdvw_state.window_centre_update~q ;
wire \sig_cdvw_state.current_window_centre[4]~4_combout ;
wire \sig_cdvw_state.current_window_centre[4]~1_combout ;
wire \sig_cdvw_state.current_window_centre[2]~q ;
wire \Add2~10 ;
wire \Add2~13_sumout ;
wire \Add4~10 ;
wire \Add4~13_sumout ;
wire \sig_cdvw_state.current_bit[3]~q ;
wire \sig_cdvw_state.current_window_centre[3]~q ;
wire \Add2~14 ;
wire \Add2~17_sumout ;
wire \Add4~14 ;
wire \Add4~17_sumout ;
wire \sig_cdvw_state.current_bit[4]~q ;
wire \sig_cdvw_state.current_window_centre[4]~q ;
wire \Add2~18 ;
wire \Add2~21_sumout ;
wire \Add4~18 ;
wire \Add4~21_sumout ;
wire \sig_cdvw_state.current_bit[5]~q ;
wire \sig_cdvw_state.current_window_centre[5]~q ;
wire \sig_cdvw_state.current_window_centre[4]~2_combout ;
wire \sig_cdvw_state.current_window_centre[4]~3_combout ;
wire \sig_cdvw_state.current_window_centre[4]~0_combout ;
wire \sig_cdvw_state.current_window_centre[0]~q ;
wire \Add2~2 ;
wire \Add2~5_sumout ;
wire \sig_cdvw_state.current_window_centre[1]~q ;
wire \v_cdvw_state~5_combout ;
wire \Add3~1_sumout ;
wire \sig_cdvw_state.current_window_size[0]~0_combout ;
wire \sig_cdvw_state.current_window_size[0]~2_combout ;
wire \sig_cdvw_state.current_window_size[0]~1_combout ;
wire \sig_cdvw_state.current_window_size[0]~q ;
wire \Add3~2 ;
wire \Add3~5_sumout ;
wire \sig_cdvw_state.current_window_size[1]~q ;
wire \Add3~6 ;
wire \Add3~9_sumout ;
wire \sig_cdvw_state.current_window_size[2]~q ;
wire \Add3~10 ;
wire \Add3~13_sumout ;
wire \sig_cdvw_state.current_window_size[3]~q ;
wire \sig_cdvw_state.largest_window_size[3]~q ;
wire \Add3~14 ;
wire \Add3~17_sumout ;
wire \sig_cdvw_state.current_window_size[4]~q ;
wire \Add3~18 ;
wire \Add3~21_sumout ;
wire \sig_cdvw_state.current_window_size[5]~q ;
wire \sig_cdvw_state.largest_window_size[5]~q ;
wire \LessThan3~1_combout ;
wire \LessThan3~2_combout ;
wire \LessThan3~3_combout ;
wire \sig_cdvw_state.largest_window_centre[1]~0_combout ;
wire \sig_cdvw_state.largest_window_centre[1]~q ;
wire \sig_cdvw_state.largest_window_centre[2]~q ;
wire \rsc_block:sig_count[2]~0_combout ;
wire \Add6~1_sumout ;
wire \sig_cdvw_state.largest_window_centre[0]~q ;
wire \Selector48~0_combout ;
wire \sig_cdvw_state.largest_window_centre[4]~q ;
wire \sig_cdvw_state.largest_window_centre[3]~q ;
wire \Add6~10 ;
wire \Add6~13_sumout ;
wire \Selector45~0_combout ;
wire \rsc_block:sig_count[3]~q ;
wire \Add6~14 ;
wire \Add6~17_sumout ;
wire \Selector44~0_combout ;
wire \Selector44~1_combout ;
wire \rsc_block:sig_count[4]~q ;
wire \Add6~18 ;
wire \Add6~21_sumout ;
wire \sig_cdvw_state.largest_window_centre[5]~q ;
wire \Selector43~0_combout ;
wire \rsc_block:sig_count[5]~q ;
wire \Add6~22 ;
wire \Add6~25_sumout ;
wire \Selector58~1_combout ;
wire \Selector42~0_combout ;
wire \rsc_block:sig_count[2]~3_combout ;
wire \rsc_block:sig_count[2]~4_combout ;
wire \rsc_block:sig_count[2]~1_combout ;
wire \rsc_block:sig_count[6]~2_combout ;
wire \rsc_block:sig_count[6]~q ;
wire \Add6~26 ;
wire \Add6~29_sumout ;
wire \Selector41~0_combout ;
wire \rsc_block:sig_count[7]~q ;
wire \Equal14~0_combout ;
wire \rsc_block:sig_curr_byte_ln_dis~q ;
wire \Add7~6 ;
wire \Add7~9_sumout ;
wire \sig_dq_pin_ctr[0]~1_combout ;
wire \sig_dq_pin_ctr[2]~q ;
wire \tp_match_block:sig_rdata_current_pin[15]~0_combout ;
wire \Add7~10 ;
wire \Add7~13_sumout ;
wire \sig_dq_pin_ctr[3]~q ;
wire \Add7~14 ;
wire \Add7~17_sumout ;
wire \sig_dq_pin_ctr[4]~q ;
wire \Mux7~0_combout ;
wire \Mux7~2_combout ;
wire \Mux7~3_combout ;
wire \Mux7~4_combout ;
wire \Mux7~5_combout ;
wire \Mux7~6_combout ;
wire \Mux7~7_combout ;
wire \Mux7~8_combout ;
wire \Mux7~9_combout ;
wire \Mux7~10_combout ;
wire \tp_match_block:sig_rdata_current_pin[14]~q ;
wire \tp_match_block:sig_rdata_current_pin[10]~q ;
wire \tp_match_block:sig_rdata_current_pin[6]~q ;
wire \Mux8~0_combout ;
wire \Mux8~2_combout ;
wire \Mux8~3_combout ;
wire \Mux8~4_combout ;
wire \Mux8~5_combout ;
wire \Mux8~6_combout ;
wire \Mux8~7_combout ;
wire \Mux8~8_combout ;
wire \Mux8~9_combout ;
wire \Mux8~10_combout ;
wire \tp_match_block:sig_rdata_current_pin[15]~q ;
wire \tp_match_block:sig_rdata_current_pin[11]~q ;
wire \Equal15~1_combout ;
wire \Mux5~0_combout ;
wire \Mux5~2_combout ;
wire \Mux5~3_combout ;
wire \Mux5~4_combout ;
wire \Mux5~5_combout ;
wire \Mux5~6_combout ;
wire \Mux5~7_combout ;
wire \Mux5~8_combout ;
wire \Mux5~9_combout ;
wire \Mux5~10_combout ;
wire \tp_match_block:sig_rdata_current_pin[12]~q ;
wire \tp_match_block:sig_rdata_current_pin[8]~q ;
wire \tp_match_block:sig_rdata_current_pin[4]~q ;
wire \tp_match_block:sig_rdata_current_pin[0]~q ;
wire \tp_match_block:sig_rdata_current_pin[2]~q ;
wire \tp_match_block:sig_rdata_current_pin[7]~q ;
wire \tp_match_block:sig_rdata_current_pin[3]~q ;
wire \Mux6~0_combout ;
wire \Mux6~2_combout ;
wire \Mux6~3_combout ;
wire \Mux6~4_combout ;
wire \Mux6~5_combout ;
wire \Mux6~6_combout ;
wire \Mux6~7_combout ;
wire \Mux6~8_combout ;
wire \Mux6~9_combout ;
wire \Mux6~10_combout ;
wire \tp_match_block:sig_rdata_current_pin[13]~q ;
wire \tp_match_block:sig_rdata_current_pin[9]~q ;
wire \tp_match_block:sig_rdata_current_pin[5]~q ;
wire \Equal15~2_combout ;
wire \Equal15~3_combout ;
wire \sig_mtp_match~q ;
wire \rsc_block:sig_count[6]~3_combout ;
wire \rsc_block:sig_count[6]~1_combout ;
wire \rsc_block:sig_count[2]~2_combout ;
wire \rsc_block:sig_count[0]~q ;
wire \Add6~2 ;
wire \Add6~6 ;
wire \Add6~9_sumout ;
wire \Selector46~0_combout ;
wire \Selector46~1_combout ;
wire \rsc_block:sig_count[2]~q ;
wire \sig_test_dq_expired~0_combout ;
wire \sig_test_dq_expired~1_combout ;
wire \rsc_block:sig_test_dq_expired~q ;
wire \Selector53~0_combout ;
wire \Selector52~0_combout ;
wire \rsc_block:sig_rsc_state.s_rsc_wait_for_idle_dimm~q ;
wire \Selector53~1_combout ;
wire \Selector53~2_combout ;
wire \rsc_block:sig_rsc_state.s_rsc_flush_datapath~q ;
wire \rsc_block:sig_rsc_last_state.s_rsc_flush_datapath~q ;
wire \Add6~5_sumout ;
wire \Selector47~0_combout ;
wire \Selector47~1_combout ;
wire \rsc_block:sig_count[1]~q ;
wire \Equal14~1_combout ;
wire \Selector54~0_combout ;
wire \rsc_block:sig_rsc_state.s_rsc_test_dq~q ;
wire \sig_dq_pin_ctr[0]~q ;
wire \Add7~2 ;
wire \Add7~5_sumout ;
wire \sig_dq_pin_ctr[1]~q ;
wire \Equal11~0_combout ;
wire \rsc_block:sig_chkd_all_dq_pins~q ;
wire \sig_rsc_cdvw_shift_in~0_combout ;
wire \sig_rsc_cdvw_shift_in~q ;
wire \v_cdvw_state~20_combout ;
wire \sig_cdvw_state.working_window[23]~0_combout ;
wire \Selector35~0_combout ;
wire \Selector68~0_combout ;
wire \Selector68~1_combout ;
wire \rsc_block:rsc_proc:v_phase_works~q ;
wire \sig_rsc_cdvw_phase~0_combout ;
wire \sig_rsc_cdvw_phase~q ;
wire \working_window~0_combout ;
wire \trk_block:mmc_seq_value_r~q ;
wire \sig_trk_cdvw_phase~0_combout ;
wire \sig_trk_cdvw_phase~q ;
wire \v_cdvw_state~56_combout ;
wire \ctrl_dgrb_r.command.cmd_rrp_seek~q ;
wire \sig_dgrb_state~48_combout ;
wire \sig_dgrb_state.s_seek_cdvw~q ;
wire \sig_cdvw_state.working_window[32]~2_combout ;
wire \v_cdvw_state~90_combout ;
wire \v_cdvw_state~91_combout ;
wire \sig_cdvw_state.working_window[63]~q ;
wire \v_cdvw_state~89_combout ;
wire \sig_cdvw_state.working_window[32]~3_combout ;
wire \sig_cdvw_state.working_window[62]~q ;
wire \v_cdvw_state~88_combout ;
wire \sig_cdvw_state.working_window[61]~q ;
wire \v_cdvw_state~87_combout ;
wire \sig_cdvw_state.working_window[60]~q ;
wire \v_cdvw_state~86_combout ;
wire \sig_cdvw_state.working_window[59]~q ;
wire \v_cdvw_state~85_combout ;
wire \sig_cdvw_state.working_window[58]~q ;
wire \v_cdvw_state~84_combout ;
wire \sig_cdvw_state.working_window[57]~q ;
wire \v_cdvw_state~83_combout ;
wire \sig_cdvw_state.working_window[56]~q ;
wire \v_cdvw_state~82_combout ;
wire \sig_cdvw_state.working_window[55]~q ;
wire \v_cdvw_state~81_combout ;
wire \sig_cdvw_state.working_window[54]~q ;
wire \v_cdvw_state~80_combout ;
wire \sig_cdvw_state.working_window[53]~q ;
wire \v_cdvw_state~79_combout ;
wire \sig_cdvw_state.working_window[52]~q ;
wire \v_cdvw_state~78_combout ;
wire \sig_cdvw_state.working_window[51]~q ;
wire \v_cdvw_state~77_combout ;
wire \sig_cdvw_state.working_window[50]~q ;
wire \v_cdvw_state~76_combout ;
wire \sig_cdvw_state.working_window[49]~q ;
wire \v_cdvw_state~75_combout ;
wire \sig_cdvw_state.working_window[48]~q ;
wire \v_cdvw_state~74_combout ;
wire \sig_cdvw_state.working_window[47]~q ;
wire \v_cdvw_state~73_combout ;
wire \sig_cdvw_state.working_window[46]~q ;
wire \v_cdvw_state~72_combout ;
wire \sig_cdvw_state.working_window[45]~q ;
wire \v_cdvw_state~71_combout ;
wire \sig_cdvw_state.working_window[44]~q ;
wire \v_cdvw_state~70_combout ;
wire \sig_cdvw_state.working_window[43]~q ;
wire \v_cdvw_state~69_combout ;
wire \sig_cdvw_state.working_window[42]~q ;
wire \v_cdvw_state~68_combout ;
wire \sig_cdvw_state.working_window[41]~q ;
wire \v_cdvw_state~67_combout ;
wire \sig_cdvw_state.working_window[40]~q ;
wire \v_cdvw_state~66_combout ;
wire \sig_cdvw_state.working_window[39]~q ;
wire \v_cdvw_state~65_combout ;
wire \sig_cdvw_state.working_window[38]~q ;
wire \v_cdvw_state~64_combout ;
wire \sig_cdvw_state.working_window[37]~q ;
wire \v_cdvw_state~63_combout ;
wire \sig_cdvw_state.working_window[36]~q ;
wire \v_cdvw_state~62_combout ;
wire \sig_cdvw_state.working_window[35]~q ;
wire \v_cdvw_state~61_combout ;
wire \sig_cdvw_state.working_window[34]~q ;
wire \v_cdvw_state~60_combout ;
wire \sig_cdvw_state.working_window[33]~q ;
wire \v_cdvw_state~59_combout ;
wire \sig_cdvw_state.working_window[32]~q ;
wire \v_cdvw_state~57_combout ;
wire \v_cdvw_state~58_combout ;
wire \sig_cdvw_state.working_window[31]~q ;
wire \v_cdvw_state~55_combout ;
wire \sig_cdvw_state.working_window[23]~4_combout ;
wire \sig_cdvw_state.working_window[23]~1_combout ;
wire \sig_cdvw_state.working_window[30]~q ;
wire \v_cdvw_state~54_combout ;
wire \sig_cdvw_state.working_window[29]~q ;
wire \v_cdvw_state~53_combout ;
wire \sig_cdvw_state.working_window[28]~q ;
wire \v_cdvw_state~52_combout ;
wire \sig_cdvw_state.working_window[27]~q ;
wire \v_cdvw_state~51_combout ;
wire \sig_cdvw_state.working_window[26]~q ;
wire \v_cdvw_state~50_combout ;
wire \sig_cdvw_state.working_window[25]~q ;
wire \v_cdvw_state~49_combout ;
wire \sig_cdvw_state.working_window[24]~q ;
wire \v_cdvw_state~48_combout ;
wire \sig_cdvw_state.working_window[23]~q ;
wire \v_cdvw_state~47_combout ;
wire \sig_cdvw_state.working_window[22]~q ;
wire \v_cdvw_state~46_combout ;
wire \sig_cdvw_state.working_window[21]~q ;
wire \v_cdvw_state~45_combout ;
wire \sig_cdvw_state.working_window[20]~q ;
wire \v_cdvw_state~44_combout ;
wire \sig_cdvw_state.working_window[19]~q ;
wire \v_cdvw_state~43_combout ;
wire \sig_cdvw_state.working_window[18]~q ;
wire \v_cdvw_state~42_combout ;
wire \sig_cdvw_state.working_window[17]~q ;
wire \v_cdvw_state~41_combout ;
wire \sig_cdvw_state.working_window[16]~q ;
wire \v_cdvw_state~40_combout ;
wire \sig_cdvw_state.working_window[15]~q ;
wire \v_cdvw_state~39_combout ;
wire \sig_cdvw_state.working_window[14]~q ;
wire \v_cdvw_state~38_combout ;
wire \sig_cdvw_state.working_window[13]~q ;
wire \v_cdvw_state~37_combout ;
wire \sig_cdvw_state.working_window[12]~q ;
wire \v_cdvw_state~36_combout ;
wire \sig_cdvw_state.working_window[11]~q ;
wire \v_cdvw_state~35_combout ;
wire \sig_cdvw_state.working_window[10]~q ;
wire \v_cdvw_state~34_combout ;
wire \sig_cdvw_state.working_window[9]~q ;
wire \v_cdvw_state~33_combout ;
wire \sig_cdvw_state.working_window[8]~q ;
wire \v_cdvw_state~32_combout ;
wire \sig_cdvw_state.working_window[7]~q ;
wire \v_cdvw_state~28_combout ;
wire \sig_cdvw_state.working_window[6]~q ;
wire \v_cdvw_state~27_combout ;
wire \sig_cdvw_state.working_window[5]~q ;
wire \v_cdvw_state~26_combout ;
wire \sig_cdvw_state.working_window[4]~q ;
wire \v_cdvw_state~25_combout ;
wire \sig_cdvw_state.working_window[3]~q ;
wire \v_cdvw_state~24_combout ;
wire \sig_cdvw_state.working_window[2]~q ;
wire \v_cdvw_state~23_combout ;
wire \sig_cdvw_state.working_window[1]~q ;
wire \v_cdvw_state~19_combout ;
wire \sig_cdvw_state.working_window[0]~q ;
wire \v_cdvw_state~8_combout ;
wire \sig_cdvw_state.valid_phase_seen~q ;
wire \v_cdvw_state~9_combout ;
wire \sig_cdvw_state.first_cycle~q ;
wire \v_cdvw_state~10_combout ;
wire \sig_cdvw_state.first_good_edge[0]~0_combout ;
wire \sig_cdvw_state.first_good_edge[2]~q ;
wire \v_cdvw_state~11_combout ;
wire \sig_cdvw_state.first_good_edge[0]~q ;
wire \v_cdvw_state~12_combout ;
wire \sig_cdvw_state.first_good_edge[1]~q ;
wire \Equal9~0_combout ;
wire \v_cdvw_state~13_combout ;
wire \sig_cdvw_state.first_good_edge[5]~q ;
wire \v_cdvw_state~14_combout ;
wire \sig_cdvw_state.first_good_edge[3]~q ;
wire \v_cdvw_state~15_combout ;
wire \sig_cdvw_state.first_good_edge[4]~q ;
wire \Equal9~1_combout ;
wire \Equal9~2_combout ;
wire \v_cdvw_state~0_combout ;
wire \v_cdvw_state~4_combout ;
wire \sig_cdvw_state.status.calculating~q ;
wire \Selector128~1_combout ;
wire \sig_trk_state~27_combout ;
wire \trk_block:sig_trk_state.s_trk_idle~q ;
wire \Selector121~0_combout ;
wire \Add10~1_sumout ;
wire \Selector126~0_combout ;
wire \trk_block:sig_remaining_samples[0]~q ;
wire \Add10~2 ;
wire \Add10~5_sumout ;
wire \Selector125~0_combout ;
wire \trk_block:sig_remaining_samples[1]~q ;
wire \Add10~6 ;
wire \Add10~9_sumout ;
wire \Selector124~0_combout ;
wire \trk_block:sig_remaining_samples[2]~q ;
wire \Add10~10 ;
wire \Add10~13_sumout ;
wire \Selector123~0_combout ;
wire \trk_block:sig_remaining_samples[3]~q ;
wire \Add10~14 ;
wire \Add10~17_sumout ;
wire \Selector122~0_combout ;
wire \trk_block:sig_remaining_samples[4]~q ;
wire \Add10~18 ;
wire \Add10~21_sumout ;
wire \Selector121~1_combout ;
wire \trk_block:sig_remaining_samples[5]~q ;
wire \Add10~22 ;
wire \Add10~25_sumout ;
wire \Selector120~0_combout ;
wire \trk_block:sig_remaining_samples[6]~q ;
wire \Add10~26 ;
wire \Add10~29_sumout ;
wire \Selector119~0_combout ;
wire \trk_block:sig_remaining_samples[7]~q ;
wire \Equal17~0_combout ;
wire \Equal17~1_combout ;
wire \sig_trk_state~14_combout ;
wire \sig_trk_state~15_combout ;
wire \Selector88~0_combout ;
wire \sig_trk_state~16_combout ;
wire \Selector95~0_combout ;
wire \trk_block:sig_mimic_cdv_found~q ;
wire \Selector128~2_combout ;
wire \Selector88~1_combout ;
wire \trk_block:sig_trk_state.s_trk_mimic_sample~q ;
wire \sig_trk_state~21_combout ;
wire \sig_trk_state~22_combout ;
wire \sig_trk_state~25_combout ;
wire \trk_block:sig_trk_state.s_trk_cdvw_drift~q ;
wire \sig_trk_last_state~0_combout ;
wire \trk_block:sig_trk_last_state.s_trk_cdvw_drift~q ;
wire \trk_block:sig_req_rsc_shift[5]~0_combout ;
wire \sig_req_rsc_shift~2_combout ;
wire \trk_block:sig_mimic_cdv[5]~0_combout ;
wire \trk_block:sig_mimic_cdv[0]~q ;
wire \Add11~1_sumout ;
wire \sig_mimic_delta~7_combout ;
wire \sig_mimic_delta~1_combout ;
wire \trk_block:sig_mimic_delta[0]~q ;
wire \Add15~1_sumout ;
wire \sig_trk_state~12_combout ;
wire \Add18~2 ;
wire \Add18~5_sumout ;
wire \Add16~2 ;
wire \Add16~5_sumout ;
wire \trk_block:sig_req_rsc_shift[5]~1_combout ;
wire \trk_block:sig_req_rsc_shift[5]~2_combout ;
wire \trk_block:sig_req_rsc_shift[5]~3_combout ;
wire \sig_req_rsc_shift~5_combout ;
wire \Add18~6 ;
wire \Add18~9_sumout ;
wire \Add16~6 ;
wire \Add16~9_sumout ;
wire \sig_req_rsc_shift~6_combout ;
wire \trk_block:sig_req_rsc_shift[2]~q ;
wire \Add18~10 ;
wire \Add18~13_sumout ;
wire \Add16~10 ;
wire \Add16~13_sumout ;
wire \sig_req_rsc_shift~7_combout ;
wire \trk_block:sig_req_rsc_shift[3]~q ;
wire \Add18~14 ;
wire \Add18~17_sumout ;
wire \Add16~14 ;
wire \Add16~17_sumout ;
wire \sig_req_rsc_shift~8_combout ;
wire \trk_block:sig_req_rsc_shift[4]~q ;
wire \trk_block:sig_req_rsc_shift[5]~5_combout ;
wire \trk_block:sig_mimic_cdv[4]~q ;
wire \trk_block:sig_mimic_cdv[3]~q ;
wire \trk_block:sig_mimic_cdv[2]~q ;
wire \trk_block:sig_mimic_cdv[1]~q ;
wire \Add11~2 ;
wire \Add11~3 ;
wire \Add11~6 ;
wire \Add11~7 ;
wire \Add11~10 ;
wire \Add11~11 ;
wire \Add11~14 ;
wire \Add11~15 ;
wire \Add11~17_sumout ;
wire \sig_mimic_delta~3_combout ;
wire \trk_block:sig_mimic_delta[4]~q ;
wire \Add11~13_sumout ;
wire \sig_mimic_delta~4_combout ;
wire \trk_block:sig_mimic_delta[3]~q ;
wire \Add11~9_sumout ;
wire \sig_mimic_delta~5_combout ;
wire \trk_block:sig_mimic_delta[2]~q ;
wire \Add11~5_sumout ;
wire \sig_mimic_delta~6_combout ;
wire \trk_block:sig_mimic_delta[1]~q ;
wire \Add12~2 ;
wire \Add12~6 ;
wire \Add12~10 ;
wire \Add12~14 ;
wire \Add12~17_sumout ;
wire \trk_block:sig_mimic_cdv[5]~q ;
wire \Add11~18 ;
wire \Add11~19 ;
wire \Add11~21_sumout ;
wire \sig_mimic_delta~2_combout ;
wire \trk_block:sig_mimic_delta[5]~q ;
wire \Add12~18 ;
wire \Add12~21_sumout ;
wire \Add12~22 ;
wire \Add12~25_sumout ;
wire \Add12~5_sumout ;
wire \Add12~9_sumout ;
wire \LessThan8~0_combout ;
wire \LessThan8~1_combout ;
wire \trk_block:sig_large_drift_seen~q ;
wire \trk_block:sig_req_rsc_shift[5]~6_combout ;
wire \Add15~2 ;
wire \Add15~6 ;
wire \Add15~10 ;
wire \Add15~14 ;
wire \Add15~18 ;
wire \Add15~21_sumout ;
wire \Add16~18 ;
wire \Add16~21_sumout ;
wire \sig_req_rsc_shift~12_combout ;
wire \trk_block:sig_req_rsc_shift[5]~q ;
wire \Add16~22 ;
wire \Add16~25_sumout ;
wire \Add15~22 ;
wire \Add15~25_sumout ;
wire \Add18~18 ;
wire \Add18~22 ;
wire \Add18~25_sumout ;
wire \sig_req_rsc_shift~9_combout ;
wire \sig_req_rsc_shift~10_combout ;
wire \trk_block:sig_req_rsc_shift[6]~q ;
wire \LessThan11~0_combout ;
wire \trk_block:sig_req_rsc_shift[5]~7_combout ;
wire \trk_block:sig_req_rsc_shift[5]~4_combout ;
wire \trk_block:sig_req_rsc_shift[1]~q ;
wire \LessThan11~1_combout ;
wire \Add18~1_sumout ;
wire \Add16~1_sumout ;
wire \sig_req_rsc_shift~11_combout ;
wire \sig_req_rsc_shift~4_combout ;
wire \trk_block:sig_req_rsc_shift[0]~q ;
wire \sig_trk_state~11_combout ;
wire \sig_trk_state~13_combout ;
wire \trk_block:sig_trk_state.s_trk_adjust_resync~q ;
wire \sig_trk_pll_inc_dec_n~1_combout ;
wire \trk_block:sig_trk_last_state.s_trk_adjust_resync~q ;
wire \sig_trk_state~17_combout ;
wire \sig_trk_state~18_combout ;
wire \sig_trk_state~26_combout ;
wire \trk_block:sig_trk_state.s_trk_cdvw_calc~q ;
wire \sig_trk_last_state~1_combout ;
wire \trk_block:sig_trk_last_state.s_trk_cdvw_calc~q ;
wire \sig_trk_state~24_combout ;
wire \trk_block:sig_trk_state.s_trk_cdvw_wait~q ;
wire \Add11~22 ;
wire \Add11~23 ;
wire \Add11~25_sumout ;
wire \sig_mimic_delta~0_combout ;
wire \trk_block:sig_mimic_delta[6]~q ;
wire \Add15~26 ;
wire \Add15~29_sumout ;
wire \sig_req_rsc_shift~1_combout ;
wire \Add16~26 ;
wire \Add16~29_sumout ;
wire \Add18~26 ;
wire \Add18~29_sumout ;
wire \sig_req_rsc_shift~16_combout ;
wire \sig_req_rsc_shift~3_combout ;
wire \trk_block:sig_req_rsc_shift[7]~q ;
wire \Add17~2_sumout ;
wire \sig_rsc_drift~0_combout ;
wire \sig_rsc_drift~1_combout ;
wire \sig_rsc_drift~7_combout ;
wire \trk_block:sig_rsc_drift[0]~q ;
wire \Add17~3 ;
wire \Add17~6_sumout ;
wire \sig_rsc_drift~6_combout ;
wire \trk_block:sig_rsc_drift[1]~q ;
wire \Selector75~0_combout ;
wire \Selector55~0_combout ;
wire \rsc_block:sig_rsc_state.s_rsc_reset_cdvw~q ;
wire \Selector71~3_combout ;
wire \Selector71~2_combout ;
wire \cal_codvw_phase[1]~q ;
wire \Selector76~0_combout ;
wire \cal_codvw_phase[0]~q ;
wire \Add9~2 ;
wire \Add9~5_sumout ;
wire \Add17~7 ;
wire \Add17~10_sumout ;
wire \sig_rsc_drift~5_combout ;
wire \trk_block:sig_rsc_drift[2]~q ;
wire \Add17~11 ;
wire \Add17~14_sumout ;
wire \sig_rsc_drift~4_combout ;
wire \trk_block:sig_rsc_drift[3]~q ;
wire \Add17~15 ;
wire \Add17~18_sumout ;
wire \sig_rsc_drift~3_combout ;
wire \trk_block:sig_rsc_drift[4]~q ;
wire \Add17~19 ;
wire \Add17~22_sumout ;
wire \sig_rsc_drift~8_combout ;
wire \trk_block:sig_rsc_drift[5]~q ;
wire \Add17~23 ;
wire \Add17~26_sumout ;
wire \sig_rsc_drift~9_combout ;
wire \trk_block:sig_rsc_drift[6]~q ;
wire \Add17~27 ;
wire \Add17~30_sumout ;
wire \sig_rsc_drift~2_combout ;
wire \trk_block:sig_rsc_drift[7]~q ;
wire \Selector71~1_combout ;
wire \cal_codvw_phase[5]~q ;
wire \Selector72~0_combout ;
wire \cal_codvw_phase[4]~q ;
wire \Selector73~0_combout ;
wire \cal_codvw_phase[3]~q ;
wire \Selector74~0_combout ;
wire \cal_codvw_phase[2]~q ;
wire \Add9~6 ;
wire \Add9~10 ;
wire \Add9~14 ;
wire \Add9~18 ;
wire \Add9~22 ;
wire \Add9~26_cout ;
wire \Add9~30_cout ;
wire \Add9~33_sumout ;
wire \rsc_block:sig_num_phase_shifts[2]~0_combout ;
wire \sig_phs_shft_busy~q ;
wire \Selector50~0_combout ;
wire \rsc_block:sig_rsc_state.s_rsc_next_phase~q ;
wire \WideOr17~0_combout ;
wire \Selector56~0_combout ;
wire \rsc_block:sig_rsc_state.s_rsc_rewind_phase~q ;
wire \rsc_block:sig_num_phase_shifts[2]~3_combout ;
wire \rsc_block:sig_num_phase_shifts[2]~1_combout ;
wire \rsc_block:sig_num_phase_shifts[5]~0_combout ;
wire \Add5~6_combout ;
wire \Add9~1_sumout ;
wire \Add5~1_combout ;
wire \Add5~4 ;
wire \Add5~8_sumout ;
wire \rsc_block:sig_num_phase_shifts[1]~0_combout ;
wire \rsc_block:sig_num_phase_shifts[1]~q ;
wire \Add9~9_sumout ;
wire \Add5~11_combout ;
wire \Add5~9 ;
wire \Add5~13_sumout ;
wire \rsc_block:sig_num_phase_shifts[2]~2_combout ;
wire \rsc_block:sig_num_phase_shifts[2]~q ;
wire \Add9~13_sumout ;
wire \Add5~16_combout ;
wire \Add5~14 ;
wire \Add5~18_sumout ;
wire \rsc_block:sig_num_phase_shifts[3]~0_combout ;
wire \rsc_block:sig_num_phase_shifts[3]~q ;
wire \Add9~21_sumout ;
wire \Add5~21_combout ;
wire \Add9~17_sumout ;
wire \Add5~22_combout ;
wire \Add5~19 ;
wire \Add5~25 ;
wire \Add5~28_sumout ;
wire \rsc_block:sig_num_phase_shifts[5]~1_combout ;
wire \rsc_block:sig_num_phase_shifts[5]~q ;
wire \Add5~24_sumout ;
wire \rsc_block:sig_num_phase_shifts[4]~0_combout ;
wire \rsc_block:sig_num_phase_shifts[4]~q ;
wire \Equal13~0_combout ;
wire \Selector71~0_combout ;
wire \Selector85~0_combout ;
wire \Selector85~1_combout ;
wire \sig_rsc_ack~q ;
wire \sig_rsc_req~16_combout ;
wire \sig_rsc_req.s_rsc_reset_cdvw~q ;
wire \sig_rsc_req~17_combout ;
wire \sig_rsc_req.s_rsc_cdvw_calc~q ;
wire \Selector49~0_combout ;
wire \rsc_block:sig_rsc_state.s_rsc_idle~q ;
wire \rsc_block:sig_rsc_last_state.s_rsc_idle~q ;
wire \Selector57~0_combout ;
wire \rsc_block:sig_rsc_state.s_rsc_cdvw_calc~q ;
wire \sig_rsc_cdvw_calc~0_combout ;
wire \sig_rsc_cdvw_calc~q ;
wire \sig_trk_cdvw_calc~0_combout ;
wire \sig_trk_cdvw_calc~q ;
wire \Selector33~0_combout ;
wire \sig_cdvw_state.current_bit[5]~1_combout ;
wire \sig_cdvw_state.current_bit[5]~2_combout ;
wire \sig_cdvw_state.current_bit[0]~q ;
wire \Add4~2 ;
wire \Add4~5_sumout ;
wire \sig_cdvw_state.current_bit[1]~q ;
wire \find_centre_of_largest_data_valid_window~0_combout ;
wire \find_centre_of_largest_data_valid_window~1_combout ;
wire \v_cdvw_state~1_combout ;
wire \sig_cdvw_state.largest_window_size[1]~q ;
wire \v_cdvw_state~16_combout ;
wire \v_cdvw_state~17_combout ;
wire \v_cdvw_state~18_combout ;
wire \sig_cdvw_state.multiple_eq_windows~q ;
wire \v_cdvw_state~3_combout ;
wire \sig_cdvw_state.status.valid_result~q ;
wire \Selector128~0_combout ;
wire \sig_trk_ack~q ;
wire \tp_match_block:sig_rdata_valid_1t~q ;
wire \tp_match_block:sig_rdata_valid_2t~q ;
wire \poa_match_proc~0_combout ;
wire \sig_poa_match_en~q ;
wire \Equal16~0_combout ;
wire \sig_poa_match~q ;
wire \sig_poa_state~0_combout ;
wire \poa_block:sig_poa_state~q ;
wire \sig_poa_ack~0_combout ;
wire \sig_poa_ack~q ;
wire \sig_dgrb_state~34_combout ;
wire \sig_dgrb_state~35_combout ;
wire \ctrl_dgrb_r.command.cmd_poa~q ;
wire \sig_dgrb_state~60_combout ;
wire \sig_dgrb_state.s_poa_cal~q ;
wire \sig_dgrb_state~36_combout ;
wire \sig_dgrb_state~37_combout ;
wire \sig_dgrb_state~67_combout ;
wire \sig_dgrb_state~39_combout ;
wire \sig_dgrb_state~40_combout ;
wire \sig_dgrb_last_state.s_adv_rd_lat_setup~q ;
wire \sig_dgrb_state~41_combout ;
wire \sig_dgrb_state~42_combout ;
wire \sig_dgrb_state~43_combout ;
wire \sig_dgrb_state~44_combout ;
wire \sig_dgrb_state~45_combout ;
wire \ctrl_dgrb_r.command.cmd_rrp_sweep~q ;
wire \sig_dgrb_state~50_combout ;
wire \sig_dgrb_state.s_test_phases~q ;
wire \Selector25~0_combout ;
wire \Selector25~1_combout ;
wire \sig_rsc_ac_access_req~0_combout ;
wire \sig_rsc_ac_access_req~q ;
wire \Selector21~0_combout ;
wire \sig_ac_req.s_ac_idle~q ;
wire \sig_addr_cmd_state~5_combout ;
wire \ac_block:sig_addr_cmd_state.s_ac_idle~q ;
wire \Selector25~2_combout ;
wire \sig_ac_req.s_ac_read_poa_mtp~q ;
wire \Selector26~0_combout ;
wire \sig_ac_req.s_ac_read_wd_lat~q ;
wire \ac_proc~0_combout ;
wire \sig_addr_cmd_state~0_combout ;
wire \sig_addr_cmd_state~4_combout ;
wire \ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ;
wire \Selector24~0_combout ;
wire \sig_ac_req.s_ac_read_rdv~q ;
wire \Selector23~1_combout ;
wire \sig_ac_req.s_ac_read_mtp~q ;
wire \ac_proc~1_combout ;
wire \ac_proc~2_combout ;
wire \sig_addr_cmd_state~6_combout ;
wire \ac_block:sig_addr_cmd_state.s_ac_relax~q ;
wire \Add22~1_sumout ;
wire \sig_setup~0_combout ;
wire \ac_block:sig_setup[4]~0_combout ;
wire \ac_block:sig_setup[0]~q ;
wire \Add22~2 ;
wire \Add22~5_sumout ;
wire \sig_setup~1_combout ;
wire \ac_block:sig_setup[1]~q ;
wire \Add22~6 ;
wire \Add22~9_sumout ;
wire \sig_setup~2_combout ;
wire \ac_block:sig_setup[2]~q ;
wire \Add22~10 ;
wire \Add22~13_sumout ;
wire \sig_setup~3_combout ;
wire \ac_block:sig_setup[3]~q ;
wire \Add22~14 ;
wire \Add22~17_sumout ;
wire \sig_setup~4_combout ;
wire \ac_block:sig_setup[4]~q ;
wire \Selector141~0_combout ;
wire \Selector141~1_combout ;
wire \sig_dimm_driving_dq~q ;
wire \sig_dgrb_state~58_combout ;
wire \sig_dgrb_state~59_combout ;
wire \sig_dgrb_state.s_adv_rd_lat~q ;
wire \ctrl_dgrb_r.command.cmd_rrp_reset~q ;
wire \sig_dgrb_state~49_combout ;
wire \sig_dgrb_state.s_reset_cdvw~q ;
wire \sig_dgrb_state~38_combout ;
wire \sig_dgrb_state~62_combout ;
wire \sig_dgrb_state~63_combout ;
wire \sig_dgrb_state~64_combout ;
wire \sig_dgrb_state~65_combout ;
wire \sig_dgrb_state~66_combout ;
wire \sig_dgrb_state.s_release_admin~q ;
wire \dgrb_state_proc~0_combout ;
wire \sig_dgrb_state~52_combout ;
wire \sig_dgrb_state~53_combout ;
wire \sig_dgrb_state~54_combout ;
wire \sig_dgrb_state~55_combout ;
wire \sig_dgrb_state.s_idle~q ;
wire \sig_dgrb_state~56_combout ;
wire \sig_dgrb_state.s_wait_admin~q ;
wire \ctrl_dgrb_r.command.cmd_prep_adv_wr_lat~q ;
wire \sig_dgrb_state~46_combout ;
wire \sig_dgrb_state.s_adv_wd_lat~q ;
wire \sig_dgrb_last_state.s_adv_wd_lat~q ;
wire \sig_wd_lat~1_combout ;
wire \dgrb_main_block:sig_wd_lat[1]~0_combout ;
wire \dgrb_main_block:sig_wd_lat[2]~q ;
wire \wd_lat[2]~0_combout ;
wire \sig_wd_lat~2_combout ;
wire \dgrb_main_block:sig_wd_lat[1]~q ;
wire \sig_wd_lat~3_combout ;
wire \dgrb_main_block:sig_wd_lat[0]~q ;
wire \wd_lat[0]~1_combout ;
wire \sig_wd_lat~4_combout ;
wire \dgrb_main_block:sig_wd_lat[3]~q ;
wire \sig_wd_lat~5_combout ;
wire \dgrb_main_block:sig_wd_lat[4]~q ;
wire \sig_burst_count~0_combout ;
wire \ac_block:sig_burst_count[0]~q ;
wire \sig_addr_cmd_state~1_combout ;
wire \ac_block:sig_addr_cmd_state.s_ac_read_wd_lat~q ;
wire \ac_block:sig_addr_cmd_last_state.s_ac_read_wd_lat~q ;
wire \Selector188~0_combout ;
wire \sig_addr_cmd_state~2_combout ;
wire \ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ;
wire \ac_block:sig_count[7]~0_combout ;
wire \Selector153~0_combout ;
wire \sig_addr_cmd_state~3_combout ;
wire \ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ;
wire \ac_block:sig_addr_cmd_last_state.s_ac_read_mtp~q ;
wire \ac_block:sig_addr_cmd_last_state.s_ac_read_rdv~q ;
wire \ac_block:sig_count[7]~1_combout ;
wire \Selector182~0_combout ;
wire \Selector186~0_combout ;
wire \Add24~14 ;
wire \Add24~17_sumout ;
wire \ac_block:sig_addr_cmd_last_state.s_ac_read_poa_mtp~q ;
wire \Selector153~1_combout ;
wire \Selector183~0_combout ;
wire \Selector183~1_combout ;
wire \Selector183~2_combout ;
wire \Selector183~3_combout ;
wire \Selector183~4_combout ;
wire \Selector183~5_combout ;
wire \ac_block:sig_count[4]~q ;
wire \Add24~18 ;
wire \Add24~21_sumout ;
wire \Selector182~1_combout ;
wire \ac_block:sig_count[5]~3_combout ;
wire \ac_block:sig_count[5]~4_combout ;
wire \ac_block:sig_count[5]~5_combout ;
wire \ac_block:sig_count[5]~0_combout ;
wire \Selector187~0_combout ;
wire \ac_block:sig_count[0]~q ;
wire \ac_block:sig_count[7]~4_combout ;
wire \ac_block:sig_count[5]~1_combout ;
wire \ac_block:sig_count[5]~q ;
wire \Equal21~1_combout ;
wire \ac_block:sig_count[5]~2_combout ;
wire \Add24~2 ;
wire \Add24~5_sumout ;
wire \Selector186~1_combout ;
wire \ac_block:sig_count[1]~q ;
wire \Add24~6 ;
wire \Add24~9_sumout ;
wire \Selector185~0_combout ;
wire \ac_block:sig_count[7]~3_combout ;
wire \ac_block:sig_count[7]~2_combout ;
wire \ac_block:sig_count[2]~q ;
wire \Add24~10 ;
wire \Add24~13_sumout ;
wire \Selector184~0_combout ;
wire \ac_block:sig_count[3]~q ;
wire \Add24~22 ;
wire \Add24~25_sumout ;
wire \Selector181~0_combout ;
wire \ac_block:sig_count[6]~q ;
wire \Add24~26 ;
wire \Add24~29_sumout ;
wire \Selector180~0_combout ;
wire \ac_block:sig_count[7]~q ;
wire \Selector189~0_combout ;
wire \Equal21~0_combout ;
wire \sig_doing_rd_count~0_combout ;
wire \ac_block:sig_doing_rd_count~q ;
wire \Selector188~1_combout ;
wire \dimm_driving_dq_proc~0_combout ;
wire \Selector188~2_combout ;
wire \Selector188~3_combout ;
wire \seq_rdata_valid_lat_dec~0_combout ;
wire \Selector189~1_combout ;
wire \Selector189~2_combout ;
wire \dgrb_ctrl_ac_nt_good~0_combout ;
wire \dgrb_ctrl_ac_nt_good~1_combout ;
wire \dgrb_ctrl_ac_nt_good~2_combout ;
wire \dgrb_ctrl_ac_nt_good~3_combout ;
wire \dgrb_ctrl_ac_nt_good~4_combout ;
wire \dgrb_ctrl_ac_nt_good~5_combout ;
wire \dgrb_ctrl_ac_nt_good~6_combout ;
wire \Selector32~0_combout ;
wire \dgrb_ctrl_ac_nt_good~7_combout ;
wire \pll_reconf_mux~0_combout ;
wire \sig_rsc_pll_inc_dec_n~0_combout ;
wire \sig_rsc_pll_inc_dec_n~q ;
wire \sig_trk_pll_inc_dec_n~2_combout ;
wire \sig_trk_pll_inc_dec_n~q ;
wire \seq_pll_inc_dec_n~0_combout ;
wire \sig_phs_shft_busy_1t~q ;
wire \Selector61~0_combout ;
wire \Selector61~1_combout ;
wire \sig_rsc_pll_start_reconfig~q ;
wire \sig_phs_shft_start~0_combout ;
wire \sig_phs_shft_start~q ;
wire \sig_trk_state~19_combout ;
wire \trk_block:sig_trk_state.s_trk_next_phase~q ;
wire \Selector127~0_combout ;
wire \sig_trk_pll_start_reconfig~q ;
wire \seq_pll_start_reconfig~0_combout ;
wire \sig_dgrb_last_state.s_release_admin~q ;
wire \ac_handshake_proc~2_combout ;
wire \sig_rsc_result[0]~0_combout ;
wire \sig_rsc_err~0_combout ;
wire \sig_rsc_err~q ;
wire \Add20~2 ;
wire \Add20~6 ;
wire \Add20~10 ;
wire \Add20~14 ;
wire \Add20~17_sumout ;
wire \Add20~1_sumout ;
wire \Add20~5_sumout ;
wire \Add20~9_sumout ;
wire \Add20~13_sumout ;
wire \Selector129~0_combout ;
wire \Add20~18 ;
wire \Add20~21_sumout ;
wire \Add20~22 ;
wire \Add20~25_sumout ;
wire \Add20~26 ;
wire \Add20~29_sumout ;
wire \Selector129~2_combout ;
wire \sig_trk_err~q ;
wire \sig_cmd_err~0_combout ;
wire \sig_cmd_err~1_combout ;
wire \sig_cmd_err~3_combout ;
wire \sig_cmd_err~4_combout ;
wire \sig_cmd_err~6_combout ;
wire \sig_cmd_err~7_combout ;
wire \sig_cmd_err~5_combout ;
wire \Selector32~2_combout ;
wire \Selector32~3_combout ;
wire \sig_cmd_err~q ;
wire \dgrb_ctrl~0_combout ;
wire \seq_pll_select~0_combout ;
wire \sig_trk_pll_select[1]~0_combout ;
wire \sig_trk_pll_select[1]~q ;
wire \seq_pll_select~1_combout ;
wire \Selector179~0_combout ;
wire \Selector179~1_combout ;
wire \btp_addr_array~0_combout ;
wire \ac_block:btp_addr_array[0][4]~q ;
wire \ctrl_dgrb_r.command_op.mtp_almt~q ;
wire \current_mtp_almt~q ;
wire \ac_block:btp_addr_array[0][3]~q ;
wire \Selector153~2_combout ;
wire \Selector153~3_combout ;
wire \sig_addr_cmd~0_combout ;
wire \Selector152~0_combout ;
wire \Selector152~1_combout ;
wire \Selector152~2_combout ;
wire \Selector153~4_combout ;
wire \Selector153~5_combout ;
wire \Selector152~3_combout ;
wire \Selector152~4_combout ;
wire \Selector152~5_combout ;
wire \Selector151~0_combout ;
wire \Selector151~1_combout ;
wire \sig_addr_cmd[0].addr[12]~0_combout ;
wire \sig_addr_cmd[0].addr[12]~1_combout ;
wire \sig_addr_cmd[0].addr[12]~2_combout ;
wire \sig_addr_cmd[0].addr[12]~3_combout ;
wire \sig_dgrb_last_state.s_idle~q ;
wire \ac_handshake_proc~3_combout ;
wire \seq_poa_lat_dec_1x~0_combout ;
wire \dgrb_ctrl~1_combout ;
wire \sig_cmd_result[2]~q ;
wire \sig_cdvw_state.largest_window_size[2]~q ;
wire \sig_trk_result[2]~q ;
wire \sig_rsc_result[2]~3_combout ;
wire \sig_rsc_result[2]~q ;
wire \dgrb_ctrl.command_result[3]~0_combout ;
wire \dgrb_ctrl.command_result[3]~1_combout ;
wire \dgrb_ctrl~2_combout ;
wire \v_cdvw_state~29_combout ;
wire \sig_cdvw_state.status.no_valid_phases~q ;
wire \Selector131~1_combout ;
wire \Selector131~0_combout ;
wire \sig_trk_result[1]~q ;
wire \v_cdvw_state~30_combout ;
wire \sig_cdvw_state.status.no_invalid_phases~q ;
wire \sig_rsc_result~1_combout ;
wire \sig_rsc_result[1]~q ;
wire \dgrb_ctrl~3_combout ;
wire \Add0~1_sumout ;
wire \dgrb_main_block:sig_count[0]~0_combout ;
wire \dgrb_main_block:sig_count[0]~q ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \dgrb_main_block:sig_count[1]~q ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \dgrb_main_block:sig_count[2]~q ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \dgrb_main_block:sig_count[3]~q ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \dgrb_main_block:sig_count[4]~q ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \dgrb_main_block:sig_count[5]~q ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \dgrb_main_block:sig_count[6]~q ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \dgrb_main_block:sig_count[7]~q ;
wire \Selector32~1_combout ;
wire \sig_cmd_result[3]~q ;
wire \sig_cdvw_state.largest_window_size[0]~q ;
wire \v_cdvw_state~31_combout ;
wire \sig_cdvw_state.status.multiple_equal_windows~q ;
wire \sig_trk_result~0_combout ;
wire \sig_trk_result[0]~q ;
wire \sig_rsc_result~2_combout ;
wire \sig_rsc_result[0]~q ;
wire \dgrb_ctrl~4_combout ;
wire \Selector129~1_combout ;
wire \sig_trk_result[4]~q ;
wire \dgrb_ctrl~5_combout ;
wire \sig_cdvw_state.largest_window_size[4]~q ;
wire \dgrb_ctrl~6_combout ;
wire \sig_trk_last_state~2_combout ;
wire \trk_block:sig_trk_last_state.s_trk_mimic_sample~q ;
wire \sig_mmc_start~1_combout ;
wire \trk_block:sig_mmc_start~q ;
wire \trk_block:mimic_sample_req:seq_mmc_start_r[0]~q ;
wire \trk_block:mimic_sample_req:seq_mmc_start_r[1]~q ;
wire \trk_block:mimic_sample_req:seq_mmc_start_r[2]~q ;
wire \seq_mmc_start~0_combout ;


arriaii_lcell_comb \Add24~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\ac_block:sig_count[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~1_sumout ),
	.cout(\Add24~2 ),
	.shareout());
defparam \Add24~1 .extended_lut = "off";
defparam \Add24~1 .lut_mask = 64'h00000000000000FF;
defparam \Add24~1 .shared_arith = "off";

dffeas \trk_block:sig_trk_state.s_trk_complete (
	.clk(clk),
	.d(\sig_trk_state~23_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_track~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_trk_state.s_trk_complete~q ),
	.prn(vcc));
defparam \trk_block:sig_trk_state.s_trk_complete .is_wysiwyg = "true";
defparam \trk_block:sig_trk_state.s_trk_complete .power_up = "low";

arriaii_lcell_comb \Add5~3 (
	.dataa(!\WideOr17~0_combout ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datac(gnd),
	.datad(!\Add5~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~3_sumout ),
	.cout(\Add5~4 ),
	.shareout());
defparam \Add5~3 .extended_lut = "off";
defparam \Add5~3 .lut_mask = 64'h0000BBBB00004400;
defparam \Add5~3 .shared_arith = "off";

arriaii_lcell_comb \Add15~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_mimic_delta[1]~q ),
	.datae(gnd),
	.dataf(!\trk_block:sig_req_rsc_shift[1]~q ),
	.datag(gnd),
	.cin(\Add15~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add15~5_sumout ),
	.cout(\Add15~6 ),
	.shareout());
defparam \Add15~5 .extended_lut = "off";
defparam \Add15~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add15~5 .shared_arith = "off";

arriaii_lcell_comb \Add15~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_mimic_delta[2]~q ),
	.datae(gnd),
	.dataf(!\trk_block:sig_req_rsc_shift[2]~q ),
	.datag(gnd),
	.cin(\Add15~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add15~9_sumout ),
	.cout(\Add15~10 ),
	.shareout());
defparam \Add15~9 .extended_lut = "off";
defparam \Add15~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add15~9 .shared_arith = "off";

arriaii_lcell_comb \Add15~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_mimic_delta[3]~q ),
	.datae(gnd),
	.dataf(!\trk_block:sig_req_rsc_shift[3]~q ),
	.datag(gnd),
	.cin(\Add15~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add15~13_sumout ),
	.cout(\Add15~14 ),
	.shareout());
defparam \Add15~13 .extended_lut = "off";
defparam \Add15~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add15~13 .shared_arith = "off";

arriaii_lcell_comb \Add15~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_mimic_delta[4]~q ),
	.datae(gnd),
	.dataf(!\trk_block:sig_req_rsc_shift[4]~q ),
	.datag(gnd),
	.cin(\Add15~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add15~17_sumout ),
	.cout(\Add15~18 ),
	.shareout());
defparam \Add15~17 .extended_lut = "off";
defparam \Add15~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add15~17 .shared_arith = "off";

arriaii_lcell_comb \Add18~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_req_rsc_shift[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add18~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add18~21_sumout ),
	.cout(\Add18~22 ),
	.shareout());
defparam \Add18~21 .extended_lut = "off";
defparam \Add18~21 .lut_mask = 64'h00000000000000FF;
defparam \Add18~21 .shared_arith = "off";

arriaii_lcell_comb \Add12~1 (
	.dataa(!\trk_block:sig_mimic_delta[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(!\trk_block:sig_mimic_delta[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~1_sumout ),
	.cout(\Add12~2 ),
	.shareout());
defparam \Add12~1 .extended_lut = "off";
defparam \Add12~1 .lut_mask = 64'h000055AA0000AAAA;
defparam \Add12~1 .shared_arith = "off";

arriaii_lcell_comb \Add12~13 (
	.dataa(!\trk_block:sig_mimic_delta[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_mimic_delta[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add12~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~13_sumout ),
	.cout(\Add12~14 ),
	.shareout());
defparam \Add12~13 .extended_lut = "off";
defparam \Add12~13 .lut_mask = 64'h0000FFFF0000AA55;
defparam \Add12~13 .shared_arith = "off";

dffeas \rsc_block:sig_rewind_direction (
	.clk(clk),
	.d(\sig_rewind_direction~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rewind_direction~q ),
	.prn(vcc));
defparam \rsc_block:sig_rewind_direction .is_wysiwyg = "true";
defparam \rsc_block:sig_rewind_direction .power_up = "low";

dffeas \rsc_block:sig_num_phase_shifts[0] (
	.clk(clk),
	.d(\rsc_block:sig_num_phase_shifts[0]~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_num_phase_shifts[0]~q ),
	.prn(vcc));
defparam \rsc_block:sig_num_phase_shifts[0] .is_wysiwyg = "true";
defparam \rsc_block:sig_num_phase_shifts[0] .power_up = "low";

arriaii_lcell_comb \sig_cmd_err~2 (
	.dataa(!q_b_4),
	.datab(!q_b_20),
	.datac(!q_b_36),
	.datad(!q_b_52),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_cmd_err~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_cmd_err~2 .extended_lut = "off";
defparam \sig_cmd_err~2 .lut_mask = 64'h8001800180018001;
defparam \sig_cmd_err~2 .shared_arith = "off";

arriaii_lcell_comb \sig_rewind_direction~0 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_reset_cdvw~q ),
	.datab(!\Add9~33_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_rewind_direction~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_rewind_direction~0 .extended_lut = "off";
defparam \sig_rewind_direction~0 .lut_mask = 64'h1111111111111111;
defparam \sig_rewind_direction~0 .shared_arith = "off";

arriaii_lcell_comb \rsc_block:sig_num_phase_shifts[0]~0 (
	.dataa(!\rsc_block:sig_num_phase_shifts[0]~q ),
	.datab(!\Add9~1_sumout ),
	.datac(!\Add5~3_sumout ),
	.datad(!\rsc_block:sig_num_phase_shifts[2]~0_combout ),
	.datae(!\rsc_block:sig_num_phase_shifts[2]~1_combout ),
	.dataf(!\rsc_block:sig_num_phase_shifts[5]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rsc_block:sig_num_phase_shifts[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rsc_block:sig_num_phase_shifts[0]~0 .extended_lut = "off";
defparam \rsc_block:sig_num_phase_shifts[0]~0 .lut_mask = 64'h555500005555F0CC;
defparam \rsc_block:sig_num_phase_shifts[0]~0 .shared_arith = "off";

arriaii_lcell_comb \sig_trk_state~20 (
	.dataa(!\trk_block:sig_trk_last_state.s_trk_adjust_resync~q ),
	.datab(!\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.datac(!\sig_trk_state~11_combout ),
	.datad(!\sig_phs_shft_end~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_trk_state~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_trk_state~20 .extended_lut = "off";
defparam \sig_trk_state~20 .lut_mask = 64'h0233023302330233;
defparam \sig_trk_state~20 .shared_arith = "off";

arriaii_lcell_comb \sig_trk_state~23 (
	.dataa(!\trk_block:sig_trk_state.s_trk_complete~q ),
	.datab(!\Selector128~2_combout ),
	.datac(!\trk_block:sig_mimic_cdv_found~q ),
	.datad(!\sig_trk_state~20_combout ),
	.datae(!\sig_trk_state~22_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_trk_state~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_trk_state~23 .extended_lut = "off";
defparam \sig_trk_state~23 .lut_mask = 64'h00FF74FF00FF74FF;
defparam \sig_trk_state~23 .shared_arith = "off";

dffeas \sig_cdvw_state.invalid_phase_seen (
	.clk(clk),
	.d(\v_cdvw_state~7_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_cdvw_state.invalid_phase_seen~q ),
	.prn(vcc));
defparam \sig_cdvw_state.invalid_phase_seen .is_wysiwyg = "true";
defparam \sig_cdvw_state.invalid_phase_seen .power_up = "low";

arriaii_lcell_comb \Equal15~0 (
	.dataa(!\tp_match_block:sig_rdata_current_pin[8]~q ),
	.datab(!\tp_match_block:sig_rdata_current_pin[9]~q ),
	.datac(!\tp_match_block:sig_rdata_current_pin[13]~q ),
	.datad(!\tp_match_block:sig_rdata_current_pin[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal15~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal15~0 .extended_lut = "off";
defparam \Equal15~0 .lut_mask = 64'h0008000800080008;
defparam \Equal15~0 .shared_arith = "off";

dffeas \tp_match_block:sig_rdata_current_pin[1] (
	.clk(clk),
	.d(\tp_match_block:sig_rdata_current_pin[5]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_current_pin[1]~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_current_pin[1] .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_current_pin[1] .power_up = "low";

arriaii_lcell_comb \LessThan3~0 (
	.dataa(!\sig_cdvw_state.largest_window_size[2]~q ),
	.datab(!\sig_cdvw_state.current_window_size[2]~q ),
	.datac(!\sig_cdvw_state.largest_window_size[1]~q ),
	.datad(!\sig_cdvw_state.current_window_size[1]~q ),
	.datae(!\sig_cdvw_state.largest_window_size[0]~q ),
	.dataf(!\sig_cdvw_state.current_window_size[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan3~0 .extended_lut = "off";
defparam \LessThan3~0 .lut_mask = 64'h22B222B2B2BB22B2;
defparam \LessThan3~0 .shared_arith = "off";

arriaii_lcell_comb \v_cdvw_state~7 (
	.dataa(!\sig_cdvw_state.status.calculating~q ),
	.datab(!\sig_cdvw_state.invalid_phase_seen~q ),
	.datac(!\v_cdvw_state~2_combout ),
	.datad(!\sig_cdvw_state.working_window[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~7 .extended_lut = "off";
defparam \v_cdvw_state~7 .lut_mask = 64'h3070307030703070;
defparam \v_cdvw_state~7 .shared_arith = "off";

dffeas single_bit_cal(
	.clk(clk),
	.d(\ctrl_dgrb_r.command_op.single_bit~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ac_muxctrl_broadcast_rcommand_req),
	.q(\single_bit_cal~q ),
	.prn(vcc));
defparam single_bit_cal.is_wysiwyg = "true";
defparam single_bit_cal.power_up = "low";

arriaii_lcell_comb \Mux6~1 (
	.dataa(!q_b_9),
	.datab(!q_b_13),
	.datac(!q_b_11),
	.datad(!q_b_15),
	.datae(!\sig_dq_pin_ctr[2]~q ),
	.dataf(!\sig_dq_pin_ctr[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux6~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux6~1 .extended_lut = "off";
defparam \Mux6~1 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux6~1 .shared_arith = "off";

arriaii_lcell_comb \Mux5~1 (
	.dataa(!q_b_1),
	.datab(!q_b_5),
	.datac(!q_b_3),
	.datad(!q_b_7),
	.datae(!\sig_dq_pin_ctr[2]~q ),
	.dataf(!\sig_dq_pin_ctr[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux5~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux5~1 .extended_lut = "off";
defparam \Mux5~1 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux5~1 .shared_arith = "off";

arriaii_lcell_comb \Mux8~1 (
	.dataa(!q_b_73),
	.datab(!q_b_77),
	.datac(!q_b_75),
	.datad(!q_b_79),
	.datae(!\sig_dq_pin_ctr[2]~q ),
	.dataf(!\sig_dq_pin_ctr[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux8~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux8~1 .extended_lut = "off";
defparam \Mux8~1 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux8~1 .shared_arith = "off";

arriaii_lcell_comb \Mux7~1 (
	.dataa(!q_b_65),
	.datab(!q_b_69),
	.datac(!q_b_67),
	.datad(!q_b_71),
	.datae(!\sig_dq_pin_ctr[2]~q ),
	.dataf(!\sig_dq_pin_ctr[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux7~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux7~1 .extended_lut = "off";
defparam \Mux7~1 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux7~1 .shared_arith = "off";

dffeas \ctrl_dgrb_r.command_op.single_bit (
	.clk(clk),
	.d(\ctrl_dgrb.command_op.single_bit ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_dgrb_r.command_op.single_bit~q ),
	.prn(vcc));
defparam \ctrl_dgrb_r.command_op.single_bit .is_wysiwyg = "true";
defparam \ctrl_dgrb_r.command_op.single_bit .power_up = "low";

dffeas \wd_lat[2] (
	.clk(clk),
	.d(\wd_lat[2]~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wd_lat_2),
	.prn(vcc));
defparam \wd_lat[2] .is_wysiwyg = "true";
defparam \wd_lat[2] .power_up = "low";

dffeas \wd_lat[1] (
	.clk(clk),
	.d(\dgrb_main_block:sig_wd_lat[1]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wd_lat_1),
	.prn(vcc));
defparam \wd_lat[1] .is_wysiwyg = "true";
defparam \wd_lat[1] .power_up = "low";

dffeas \wd_lat[0] (
	.clk(clk),
	.d(\wd_lat[0]~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wd_lat_0),
	.prn(vcc));
defparam \wd_lat[0] .is_wysiwyg = "true";
defparam \wd_lat[0] .power_up = "low";

dffeas \wd_lat[3] (
	.clk(clk),
	.d(\dgrb_main_block:sig_wd_lat[3]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wd_lat_3),
	.prn(vcc));
defparam \wd_lat[3] .is_wysiwyg = "true";
defparam \wd_lat[3] .power_up = "low";

dffeas \wd_lat[4] (
	.clk(clk),
	.d(\dgrb_main_block:sig_wd_lat[4]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wd_lat_4),
	.prn(vcc));
defparam \wd_lat[4] .is_wysiwyg = "true";
defparam \wd_lat[4] .power_up = "low";

dffeas \sig_doing_rd[0] (
	.clk(clk),
	.d(\Selector188~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sig_doing_rd_0),
	.prn(vcc));
defparam \sig_doing_rd[0] .is_wysiwyg = "true";
defparam \sig_doing_rd[0] .power_up = "low";

dffeas seq_rdata_valid_lat_dec(
	.clk(clk),
	.d(\seq_rdata_valid_lat_dec~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_rdata_valid_lat_dec1),
	.prn(vcc));
defparam seq_rdata_valid_lat_dec.is_wysiwyg = "true";
defparam seq_rdata_valid_lat_dec.power_up = "low";

dffeas \sig_doing_rd[4] (
	.clk(clk),
	.d(\Selector189~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sig_doing_rd_4),
	.prn(vcc));
defparam \sig_doing_rd[4] .is_wysiwyg = "true";
defparam \sig_doing_rd[4] .power_up = "low";

dffeas dgrb_ctrl_ac_nt_good(
	.clk(clk),
	.d(\dgrb_ctrl_ac_nt_good~7_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgrb_ctrl_ac_nt_good1),
	.prn(vcc));
defparam dgrb_ctrl_ac_nt_good.is_wysiwyg = "true";
defparam dgrb_ctrl_ac_nt_good.power_up = "low";

dffeas seq_pll_inc_dec_n(
	.clk(clk),
	.d(\seq_pll_inc_dec_n~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_pll_inc_dec_n1),
	.prn(vcc));
defparam seq_pll_inc_dec_n.is_wysiwyg = "true";
defparam seq_pll_inc_dec_n.power_up = "low";

dffeas seq_pll_start_reconfig(
	.clk(clk),
	.d(\seq_pll_start_reconfig~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_pll_start_reconfig1),
	.prn(vcc));
defparam seq_pll_start_reconfig.is_wysiwyg = "true";
defparam seq_pll_start_reconfig.power_up = "low";

dffeas \dgrb_ctrl.command_done (
	.clk(clk),
	.d(\ac_handshake_proc~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgrb_ctrlcommand_done),
	.prn(vcc));
defparam \dgrb_ctrl.command_done .is_wysiwyg = "true";
defparam \dgrb_ctrl.command_done .power_up = "low";

dffeas \dgrb_ctrl.command_err (
	.clk(clk),
	.d(\dgrb_ctrl~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgrb_ctrlcommand_err),
	.prn(vcc));
defparam \dgrb_ctrl.command_err .is_wysiwyg = "true";
defparam \dgrb_ctrl.command_err .power_up = "low";

dffeas \seq_pll_select[0] (
	.clk(clk),
	.d(\seq_pll_select~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_pll_select_0),
	.prn(vcc));
defparam \seq_pll_select[0] .is_wysiwyg = "true";
defparam \seq_pll_select[0] .power_up = "low";

dffeas \seq_pll_select[1] (
	.clk(clk),
	.d(\seq_pll_select~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_pll_select_1),
	.prn(vcc));
defparam \seq_pll_select[1] .is_wysiwyg = "true";
defparam \seq_pll_select[1] .power_up = "low";

dffeas dgrb_ac_access_req(
	.clk(clk),
	.d(\dimm_driving_dq_proc~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgrb_ac_access_req1),
	.prn(vcc));
defparam dgrb_ac_access_req.is_wysiwyg = "true";
defparam dgrb_ac_access_req.power_up = "low";

dffeas \sig_addr_cmd[1].cs_n[0] (
	.clk(clk),
	.d(\Selector179~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sig_addr_cmd1cs_n0),
	.prn(vcc));
defparam \sig_addr_cmd[1].cs_n[0] .is_wysiwyg = "true";
defparam \sig_addr_cmd[1].cs_n[0] .power_up = "low";

dffeas \sig_addr_cmd[0].addr[3] (
	.clk(clk),
	.d(\Selector153~5_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sig_addr_cmd0addr3),
	.prn(vcc));
defparam \sig_addr_cmd[0].addr[3] .is_wysiwyg = "true";
defparam \sig_addr_cmd[0].addr[3] .power_up = "low";

dffeas \sig_addr_cmd[0].addr[4] (
	.clk(clk),
	.d(\Selector152~5_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sig_addr_cmd0addr4),
	.prn(vcc));
defparam \sig_addr_cmd[0].addr[4] .is_wysiwyg = "true";
defparam \sig_addr_cmd[0].addr[4] .power_up = "low";

dffeas \sig_addr_cmd[0].addr[5] (
	.clk(clk),
	.d(\Selector151~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sig_addr_cmd0addr5),
	.prn(vcc));
defparam \sig_addr_cmd[0].addr[5] .is_wysiwyg = "true";
defparam \sig_addr_cmd[0].addr[5] .power_up = "low";

dffeas \sig_addr_cmd[0].addr[12] (
	.clk(clk),
	.d(\sig_addr_cmd[0].addr[12]~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sig_addr_cmd0addr12),
	.prn(vcc));
defparam \sig_addr_cmd[0].addr[12] .is_wysiwyg = "true";
defparam \sig_addr_cmd[0].addr[12] .power_up = "low";

dffeas \dgrb_ctrl.command_ack (
	.clk(clk),
	.d(\ac_handshake_proc~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgrb_ctrlcommand_ack),
	.prn(vcc));
defparam \dgrb_ctrl.command_ack .is_wysiwyg = "true";
defparam \dgrb_ctrl.command_ack .power_up = "low";

dffeas \seq_poa_lat_dec_1x[0] (
	.clk(clk),
	.d(\seq_poa_lat_dec_1x~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_poa_lat_dec_1x_0),
	.prn(vcc));
defparam \seq_poa_lat_dec_1x[0] .is_wysiwyg = "true";
defparam \seq_poa_lat_dec_1x[0] .power_up = "low";

dffeas \dgrb_ctrl.command_result[5] (
	.clk(clk),
	.d(\dgrb_ctrl~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgrb_ctrlcommand_result_5),
	.prn(vcc));
defparam \dgrb_ctrl.command_result[5] .is_wysiwyg = "true";
defparam \dgrb_ctrl.command_result[5] .power_up = "low";

dffeas \dgrb_ctrl.command_result[2] (
	.clk(clk),
	.d(\dgrb_ctrl~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgrb_ctrlcommand_result_2),
	.prn(vcc));
defparam \dgrb_ctrl.command_result[2] .is_wysiwyg = "true";
defparam \dgrb_ctrl.command_result[2] .power_up = "low";

dffeas \dgrb_ctrl.command_result[1] (
	.clk(clk),
	.d(\dgrb_ctrl~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgrb_ctrlcommand_result_1),
	.prn(vcc));
defparam \dgrb_ctrl.command_result[1] .is_wysiwyg = "true";
defparam \dgrb_ctrl.command_result[1] .power_up = "low";

dffeas \dgrb_ctrl.command_result[0] (
	.clk(clk),
	.d(\dgrb_ctrl~4_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgrb_ctrlcommand_result_0),
	.prn(vcc));
defparam \dgrb_ctrl.command_result[0] .is_wysiwyg = "true";
defparam \dgrb_ctrl.command_result[0] .power_up = "low";

dffeas \dgrb_ctrl.command_result[3] (
	.clk(clk),
	.d(\dgrb_ctrl~5_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgrb_ctrlcommand_result_3),
	.prn(vcc));
defparam \dgrb_ctrl.command_result[3] .is_wysiwyg = "true";
defparam \dgrb_ctrl.command_result[3] .power_up = "low";

dffeas \dgrb_ctrl.command_result[4] (
	.clk(clk),
	.d(\dgrb_ctrl~6_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgrb_ctrlcommand_result_4),
	.prn(vcc));
defparam \dgrb_ctrl.command_result[4] .is_wysiwyg = "true";
defparam \dgrb_ctrl.command_result[4] .power_up = "low";

dffeas seq_mmc_start(
	.clk(clk),
	.d(\seq_mmc_start~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(seq_mmc_start1),
	.prn(vcc));
defparam seq_mmc_start.is_wysiwyg = "true";
defparam seq_mmc_start.power_up = "low";

dffeas \ac_block:sig_addr_cmd_last_state.s_ac_relax (
	.clk(clk),
	.d(\ac_block:sig_addr_cmd_state.s_ac_relax~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_block:sig_addr_cmd_last_state.s_ac_relax~q ),
	.prn(vcc));
defparam \ac_block:sig_addr_cmd_last_state.s_ac_relax .is_wysiwyg = "true";
defparam \ac_block:sig_addr_cmd_last_state.s_ac_relax .power_up = "low";

dffeas \ctrl_dgrb_r.command.cmd_rdv (
	.clk(clk),
	.d(\ctrl_dgrb.command.cmd_rdv ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_dgrb_r.command.cmd_rdv~q ),
	.prn(vcc));
defparam \ctrl_dgrb_r.command.cmd_rdv .is_wysiwyg = "true";
defparam \ctrl_dgrb_r.command.cmd_rdv .power_up = "low";

arriaii_lcell_comb \sig_dgrb_state~47 (
	.dataa(!\sig_dgrb_state.s_rdata_valid_align~q ),
	.datab(!\sig_dgrb_state.s_wait_admin~q ),
	.datac(!\sig_dgrb_state~45_combout ),
	.datad(!\ctrl_dgrb_r.command.cmd_rdv~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~47 .extended_lut = "off";
defparam \sig_dgrb_state~47 .lut_mask = 64'h0407040704070407;
defparam \sig_dgrb_state~47 .shared_arith = "off";

dffeas \sig_dgrb_state.s_rdata_valid_align (
	.clk(clk),
	.d(\sig_dgrb_state~47_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgrb_state.s_rdata_valid_align~q ),
	.prn(vcc));
defparam \sig_dgrb_state.s_rdata_valid_align .is_wysiwyg = "true";
defparam \sig_dgrb_state.s_rdata_valid_align .power_up = "low";

dffeas \ctrl_dgrb_r.command.cmd_prep_adv_rd_lat (
	.clk(clk),
	.d(\ctrl_dgrb.command.cmd_prep_adv_rd_lat ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_dgrb_r.command.cmd_prep_adv_rd_lat~q ),
	.prn(vcc));
defparam \ctrl_dgrb_r.command.cmd_prep_adv_rd_lat .is_wysiwyg = "true";
defparam \ctrl_dgrb_r.command.cmd_prep_adv_rd_lat .power_up = "low";

arriaii_lcell_comb \sig_dgrb_state~57 (
	.dataa(!\sig_dgrb_state.s_wait_admin~q ),
	.datab(!\sig_dgrb_state.s_adv_rd_lat_setup~q ),
	.datac(!\sig_dgrb_state~45_combout ),
	.datad(!\ctrl_dgrb_r.command.cmd_prep_adv_rd_lat~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~57_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~57 .extended_lut = "off";
defparam \sig_dgrb_state~57 .lut_mask = 64'h0207020702070207;
defparam \sig_dgrb_state~57 .shared_arith = "off";

dffeas \sig_dgrb_state.s_adv_rd_lat_setup (
	.clk(clk),
	.d(\sig_dgrb_state~57_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgrb_state.s_adv_rd_lat_setup~q ),
	.prn(vcc));
defparam \sig_dgrb_state.s_adv_rd_lat_setup .is_wysiwyg = "true";
defparam \sig_dgrb_state.s_adv_rd_lat_setup .power_up = "low";

arriaii_lcell_comb \v_aligned~0 (
	.dataa(!q_b_0),
	.datab(!q_b_64),
	.datac(!q_b_8),
	.datad(!q_b_72),
	.datae(!rdata_valid[0]),
	.dataf(!seq_rdata_valid_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_aligned~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_aligned~0 .extended_lut = "off";
defparam \v_aligned~0 .lut_mask = 64'h0000A0A0CC00ECA0;
defparam \v_aligned~0 .shared_arith = "off";

dffeas \ctrl_dgrb_r.command.cmd_tr_due (
	.clk(clk),
	.d(\ctrl_dgrb.command.cmd_tr_due ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_dgrb_r.command.cmd_tr_due~q ),
	.prn(vcc));
defparam \ctrl_dgrb_r.command.cmd_tr_due .is_wysiwyg = "true";
defparam \ctrl_dgrb_r.command.cmd_tr_due .power_up = "low";

arriaii_lcell_comb \sig_dgrb_state~51 (
	.dataa(!\sig_dgrb_state.s_track~q ),
	.datab(!\sig_dgrb_state.s_wait_admin~q ),
	.datac(!\sig_dgrb_state~45_combout ),
	.datad(!\ctrl_dgrb_r.command.cmd_tr_due~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~51 .extended_lut = "off";
defparam \sig_dgrb_state~51 .lut_mask = 64'h0407040704070407;
defparam \sig_dgrb_state~51 .shared_arith = "off";

dffeas \sig_dgrb_state.s_track (
	.clk(clk),
	.d(\sig_dgrb_state~51_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgrb_state.s_track~q ),
	.prn(vcc));
defparam \sig_dgrb_state.s_track .is_wysiwyg = "true";
defparam \sig_dgrb_state.s_track .power_up = "low";

arriaii_lcell_comb \Add4~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sig_cdvw_state.current_bit[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~1_sumout ),
	.cout(\Add4~2 ),
	.shareout());
defparam \Add4~1 .extended_lut = "off";
defparam \Add4~1 .lut_mask = 64'h00000000000000FF;
defparam \Add4~1 .shared_arith = "off";

dffeas \ctrl_dgrb_r.command.cmd_read_mtp (
	.clk(clk),
	.d(\ctrl_dgrb.command.cmd_read_mtp ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_dgrb_r.command.cmd_read_mtp~q ),
	.prn(vcc));
defparam \ctrl_dgrb_r.command.cmd_read_mtp .is_wysiwyg = "true";
defparam \ctrl_dgrb_r.command.cmd_read_mtp .power_up = "low";

arriaii_lcell_comb \sig_dgrb_state~61 (
	.dataa(!\sig_dgrb_state.s_wait_admin~q ),
	.datab(!\sig_dgrb_state.s_read_mtp~q ),
	.datac(!\sig_dgrb_state~45_combout ),
	.datad(!\ctrl_dgrb_r.command.cmd_read_mtp~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~61_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~61 .extended_lut = "off";
defparam \sig_dgrb_state~61 .lut_mask = 64'h0207020702070207;
defparam \sig_dgrb_state~61 .shared_arith = "off";

dffeas \sig_dgrb_state.s_read_mtp (
	.clk(clk),
	.d(\sig_dgrb_state~61_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgrb_state.s_read_mtp~q ),
	.prn(vcc));
defparam \sig_dgrb_state.s_read_mtp .is_wysiwyg = "true";
defparam \sig_dgrb_state.s_read_mtp .power_up = "low";

dffeas \cdvw_block:sig_cdvw_calc_1t (
	.clk(clk),
	.d(\Selector33~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\cdvw_block:sig_cdvw_calc_1t~q ),
	.prn(vcc));
defparam \cdvw_block:sig_cdvw_calc_1t .is_wysiwyg = "true";
defparam \cdvw_block:sig_cdvw_calc_1t .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~2 (
	.dataa(!\cdvw_proc~1_combout ),
	.datab(!\cdvw_block:sig_cdvw_calc_1t~q ),
	.datac(!\Selector33~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~2 .extended_lut = "off";
defparam \v_cdvw_state~2 .lut_mask = 64'h5D5D5D5D5D5D5D5D;
defparam \v_cdvw_state~2 .shared_arith = "off";

dffeas \sig_dgrb_last_state.s_track (
	.clk(clk),
	.d(\sig_dgrb_state.s_track~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgrb_last_state.s_track~q ),
	.prn(vcc));
defparam \sig_dgrb_last_state.s_track .is_wysiwyg = "true";
defparam \sig_dgrb_last_state.s_track .power_up = "low";

arriaii_lcell_comb \cdvw_proc~2 (
	.dataa(!\cdvw_block:sig_cdvw_calc_1t~q ),
	.datab(!\Selector33~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cdvw_proc~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cdvw_proc~2 .extended_lut = "off";
defparam \cdvw_proc~2 .lut_mask = 64'h2222222222222222;
defparam \cdvw_proc~2 .shared_arith = "off";

dffeas \trk_block:mmc_seq_req_sync:v_mmc_seq_done_1r (
	.clk(clk),
	.d(mmc_seq_done),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:mmc_seq_req_sync:v_mmc_seq_done_1r~q ),
	.prn(vcc));
defparam \trk_block:mmc_seq_req_sync:v_mmc_seq_done_1r .is_wysiwyg = "true";
defparam \trk_block:mmc_seq_req_sync:v_mmc_seq_done_1r .power_up = "low";

dffeas \trk_block:mmc_seq_req_sync:v_mmc_seq_done_2r (
	.clk(clk),
	.d(\trk_block:mmc_seq_req_sync:v_mmc_seq_done_1r~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:mmc_seq_req_sync:v_mmc_seq_done_2r~q ),
	.prn(vcc));
defparam \trk_block:mmc_seq_req_sync:v_mmc_seq_done_2r .is_wysiwyg = "true";
defparam \trk_block:mmc_seq_req_sync:v_mmc_seq_done_2r .power_up = "low";

dffeas \trk_block:mmc_seq_req_sync:v_mmc_seq_done_3r (
	.clk(clk),
	.d(\trk_block:mmc_seq_req_sync:v_mmc_seq_done_2r~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:mmc_seq_req_sync:v_mmc_seq_done_3r~q ),
	.prn(vcc));
defparam \trk_block:mmc_seq_req_sync:v_mmc_seq_done_3r .is_wysiwyg = "true";
defparam \trk_block:mmc_seq_req_sync:v_mmc_seq_done_3r .power_up = "low";

dffeas \trk_block:sig_mmc_seq_done_1t (
	.clk(clk),
	.d(\trk_block:mmc_seq_req_sync:v_mmc_seq_done_3r~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_mmc_seq_done_1t~q ),
	.prn(vcc));
defparam \trk_block:sig_mmc_seq_done_1t .is_wysiwyg = "true";
defparam \trk_block:sig_mmc_seq_done_1t .power_up = "low";

arriaii_lcell_comb \shift_in_mmc_seq_value~0 (
	.dataa(!\trk_block:mmc_seq_req_sync:v_mmc_seq_done_3r~q ),
	.datab(!\trk_block:sig_mmc_seq_done_1t~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\shift_in_mmc_seq_value~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \shift_in_mmc_seq_value~0 .extended_lut = "off";
defparam \shift_in_mmc_seq_value~0 .lut_mask = 64'h2222222222222222;
defparam \shift_in_mmc_seq_value~0 .shared_arith = "off";

dffeas sig_trk_cdvw_shift_in(
	.clk(clk),
	.d(\shift_in_mmc_seq_value~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_trk_cdvw_shift_in~q ),
	.prn(vcc));
defparam sig_trk_cdvw_shift_in.is_wysiwyg = "true";
defparam sig_trk_cdvw_shift_in.power_up = "low";

arriaii_lcell_comb \Add7~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sig_dq_pin_ctr[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~1_sumout ),
	.cout(\Add7~2 ),
	.shareout());
defparam \Add7~1 .extended_lut = "off";
defparam \Add7~1 .lut_mask = 64'h00000000000000FF;
defparam \Add7~1 .shared_arith = "off";

arriaii_lcell_comb \single_bit_cal~_wirecell (
	.dataa(!\single_bit_cal~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\single_bit_cal~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \single_bit_cal~_wirecell .extended_lut = "off";
defparam \single_bit_cal~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \single_bit_cal~_wirecell .shared_arith = "off";

dffeas \phs_shft_busy_reg:phs_shft_busy_1r (
	.clk(clk),
	.d(phs_shft_busy),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\phs_shft_busy_reg:phs_shft_busy_1r~q ),
	.prn(vcc));
defparam \phs_shft_busy_reg:phs_shft_busy_1r .is_wysiwyg = "true";
defparam \phs_shft_busy_reg:phs_shft_busy_1r .power_up = "low";

dffeas \phs_shft_busy_reg:phs_shft_busy_2r (
	.clk(clk),
	.d(\phs_shft_busy_reg:phs_shft_busy_1r~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\phs_shft_busy_reg:phs_shft_busy_2r~q ),
	.prn(vcc));
defparam \phs_shft_busy_reg:phs_shft_busy_2r .is_wysiwyg = "true";
defparam \phs_shft_busy_reg:phs_shft_busy_2r .power_up = "low";

arriaii_lcell_comb \sig_phs_shft_end~0 (
	.dataa(!\sig_phs_shft_busy~q ),
	.datab(!\phs_shft_busy_reg:phs_shft_busy_2r~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_phs_shft_end~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_phs_shft_end~0 .extended_lut = "off";
defparam \sig_phs_shft_end~0 .lut_mask = 64'h4444444444444444;
defparam \sig_phs_shft_end~0 .shared_arith = "off";

dffeas sig_phs_shft_end(
	.clk(clk),
	.d(\sig_phs_shft_end~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_phs_shft_end~q ),
	.prn(vcc));
defparam sig_phs_shft_end.is_wysiwyg = "true";
defparam sig_phs_shft_end.power_up = "low";

arriaii_lcell_comb \Selector23~0 (
	.dataa(!\sig_dgrb_state.s_test_phases~q ),
	.datab(!\sig_rsc_ack~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector23~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector23~0 .extended_lut = "off";
defparam \Selector23~0 .lut_mask = 64'h4444444444444444;
defparam \Selector23~0 .shared_arith = "off";

dffeas \sig_rsc_req.s_rsc_test_phase (
	.clk(clk),
	.d(\Selector23~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_rsc_req.s_rsc_test_phase~q ),
	.prn(vcc));
defparam \sig_rsc_req.s_rsc_test_phase .is_wysiwyg = "true";
defparam \sig_rsc_req.s_rsc_test_phase .power_up = "low";

arriaii_lcell_comb \Selector51~0 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_next_phase~q ),
	.datab(!\sig_phs_shft_end~q ),
	.datac(!\rsc_block:sig_rsc_state.s_rsc_idle~q ),
	.datad(!\rsc_block:sig_rsc_last_state.s_rsc_idle~q ),
	.datae(!\sig_rsc_req.s_rsc_test_phase~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector51~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector51~0 .extended_lut = "off";
defparam \Selector51~0 .lut_mask = 64'h1111F1111111F111;
defparam \Selector51~0 .shared_arith = "off";

dffeas \rsc_block:sig_rsc_state.s_rsc_test_phase (
	.clk(clk),
	.d(\Selector51~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rsc_state.s_rsc_test_phase~q ),
	.prn(vcc));
defparam \rsc_block:sig_rsc_state.s_rsc_test_phase .is_wysiwyg = "true";
defparam \rsc_block:sig_rsc_state.s_rsc_test_phase .power_up = "low";

arriaii_lcell_comb \sig_dq_pin_ctr[0]~0 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_test_phase~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dq_pin_ctr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dq_pin_ctr[0]~0 .extended_lut = "off";
defparam \sig_dq_pin_ctr[0]~0 .lut_mask = 64'h8888888888888888;
defparam \sig_dq_pin_ctr[0]~0 .shared_arith = "off";

dffeas \rsc_block:sig_rsc_last_state.s_rsc_test_dq (
	.clk(clk),
	.d(\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rsc_last_state.s_rsc_test_dq~q ),
	.prn(vcc));
defparam \rsc_block:sig_rsc_last_state.s_rsc_test_dq .is_wysiwyg = "true";
defparam \rsc_block:sig_rsc_last_state.s_rsc_test_dq .power_up = "low";

dffeas \rsc_block:sig_rsc_last_state.s_rsc_seek_cdvw (
	.clk(clk),
	.d(\rsc_block:sig_rsc_state.s_rsc_seek_cdvw~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rsc_last_state.s_rsc_seek_cdvw~q ),
	.prn(vcc));
defparam \rsc_block:sig_rsc_last_state.s_rsc_seek_cdvw .is_wysiwyg = "true";
defparam \rsc_block:sig_rsc_last_state.s_rsc_seek_cdvw .power_up = "low";

dffeas \rsc_block:sig_rsc_last_state.s_rsc_cdvw_calc (
	.clk(clk),
	.d(\rsc_block:sig_rsc_state.s_rsc_cdvw_calc~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rsc_last_state.s_rsc_cdvw_calc~q ),
	.prn(vcc));
defparam \rsc_block:sig_rsc_last_state.s_rsc_cdvw_calc .is_wysiwyg = "true";
defparam \rsc_block:sig_rsc_last_state.s_rsc_cdvw_calc .power_up = "low";

arriaii_lcell_comb \Selector58~2 (
	.dataa(!\sig_cdvw_state.status.calculating~q ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_cdvw_wait~q ),
	.datac(!\rsc_block:sig_rsc_last_state.s_rsc_cdvw_calc~q ),
	.datad(!\rsc_block:sig_rsc_state.s_rsc_cdvw_calc~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector58~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector58~2 .extended_lut = "off";
defparam \Selector58~2 .lut_mask = 64'h111F111F111F111F;
defparam \Selector58~2 .shared_arith = "off";

dffeas \rsc_block:sig_rsc_state.s_rsc_cdvw_wait (
	.clk(clk),
	.d(\Selector58~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rsc_state.s_rsc_cdvw_wait~q ),
	.prn(vcc));
defparam \rsc_block:sig_rsc_state.s_rsc_cdvw_wait .is_wysiwyg = "true";
defparam \rsc_block:sig_rsc_state.s_rsc_cdvw_wait .power_up = "low";

arriaii_lcell_comb \Selector59~0 (
	.dataa(!\sig_dgrb_state.s_read_mtp~q ),
	.datab(!\Equal14~1_combout ),
	.datac(!\rsc_block:sig_rsc_last_state.s_rsc_seek_cdvw~q ),
	.datad(!\rsc_block:sig_rsc_state.s_rsc_seek_cdvw~q ),
	.datae(!\sig_cdvw_state.status.valid_result~q ),
	.dataf(!\rsc_block:sig_rsc_state.s_rsc_cdvw_wait~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector59~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector59~0 .extended_lut = "off";
defparam \Selector59~0 .lut_mask = 64'h00FC00FC00FCAAFE;
defparam \Selector59~0 .shared_arith = "off";

dffeas \rsc_block:sig_rsc_state.s_rsc_seek_cdvw (
	.clk(clk),
	.d(\Selector59~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rsc_state.s_rsc_seek_cdvw~q ),
	.prn(vcc));
defparam \rsc_block:sig_rsc_state.s_rsc_seek_cdvw .is_wysiwyg = "true";
defparam \rsc_block:sig_rsc_state.s_rsc_seek_cdvw .power_up = "low";

arriaii_lcell_comb \rsc_block:sig_count[6]~0 (
	.dataa(!\rsc_block:sig_rsc_last_state.s_rsc_seek_cdvw~q ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_seek_cdvw~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rsc_block:sig_count[6]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rsc_block:sig_count[6]~0 .extended_lut = "off";
defparam \rsc_block:sig_count[6]~0 .lut_mask = 64'h2222222222222222;
defparam \rsc_block:sig_count[6]~0 .shared_arith = "off";

arriaii_lcell_comb \Add2~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sig_cdvw_state.current_window_centre[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~1_sumout ),
	.cout(\Add2~2 ),
	.shareout());
defparam \Add2~1 .extended_lut = "off";
defparam \Add2~1 .lut_mask = 64'h00000000000000FF;
defparam \Add2~1 .shared_arith = "off";

arriaii_lcell_comb \cdvw_proc~1 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cdvw_proc~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cdvw_proc~1 .extended_lut = "off";
defparam \cdvw_proc~1 .lut_mask = 64'h7575757575757575;
defparam \cdvw_proc~1 .shared_arith = "off";

arriaii_lcell_comb \Add2~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sig_cdvw_state.current_window_centre[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~5_sumout ),
	.cout(\Add2~6 ),
	.shareout());
defparam \Add2~5 .extended_lut = "off";
defparam \Add2~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add2~5 .shared_arith = "off";

arriaii_lcell_comb \Add2~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sig_cdvw_state.current_window_centre[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~9_sumout ),
	.cout(\Add2~10 ),
	.shareout());
defparam \Add2~9 .extended_lut = "off";
defparam \Add2~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add2~9 .shared_arith = "off";

arriaii_lcell_comb \Add4~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sig_cdvw_state.current_bit[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~5_sumout ),
	.cout(\Add4~6 ),
	.shareout());
defparam \Add4~5 .extended_lut = "off";
defparam \Add4~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add4~5 .shared_arith = "off";

arriaii_lcell_comb \Add4~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sig_cdvw_state.current_bit[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~9_sumout ),
	.cout(\Add4~10 ),
	.shareout());
defparam \Add4~9 .extended_lut = "off";
defparam \Add4~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add4~9 .shared_arith = "off";

arriaii_lcell_comb \sig_cdvw_state.current_bit[5]~0 (
	.dataa(!\sig_cdvw_state.status.calculating~q ),
	.datab(!\cdvw_proc~1_combout ),
	.datac(!\cdvw_block:sig_cdvw_calc_1t~q ),
	.datad(!\Selector33~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_cdvw_state.current_bit[5]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_cdvw_state.current_bit[5]~0 .extended_lut = "off";
defparam \sig_cdvw_state.current_bit[5]~0 .lut_mask = 64'h77F777F777F777F7;
defparam \sig_cdvw_state.current_bit[5]~0 .shared_arith = "off";

dffeas \sig_cdvw_state.current_bit[2] (
	.clk(clk),
	.d(\Add4~9_sumout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_bit[5]~2_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.current_bit[5]~0_combout ),
	.q(\sig_cdvw_state.current_bit[2]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_bit[2] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_bit[2] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~21 (
	.dataa(!\v_cdvw_state~2_combout ),
	.datab(!\sig_cdvw_state.working_window[0]~q ),
	.datac(!\sig_cdvw_state.last_bit_value~q ),
	.datad(!\sig_cdvw_state.working_window[23]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~21 .extended_lut = "off";
defparam \v_cdvw_state~21 .lut_mask = 64'h220A220A220A220A;
defparam \v_cdvw_state~21 .shared_arith = "off";

dffeas \sig_cdvw_state.last_bit_value (
	.clk(clk),
	.d(\v_cdvw_state~21_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_cdvw_state.last_bit_value~q ),
	.prn(vcc));
defparam \sig_cdvw_state.last_bit_value .is_wysiwyg = "true";
defparam \sig_cdvw_state.last_bit_value .power_up = "low";

arriaii_lcell_comb \find_centre_of_largest_data_valid_window~2 (
	.dataa(!\sig_cdvw_state.working_window[0]~q ),
	.datab(!\sig_cdvw_state.last_bit_value~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\find_centre_of_largest_data_valid_window~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \find_centre_of_largest_data_valid_window~2 .extended_lut = "off";
defparam \find_centre_of_largest_data_valid_window~2 .lut_mask = 64'h2222222222222222;
defparam \find_centre_of_largest_data_valid_window~2 .shared_arith = "off";

arriaii_lcell_comb \v_cdvw_state~6 (
	.dataa(!\sig_cdvw_state.status.calculating~q ),
	.datab(!\sig_cdvw_state.found_a_good_edge~q ),
	.datac(!\v_cdvw_state~2_combout ),
	.datad(!\find_centre_of_largest_data_valid_window~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~6 .extended_lut = "off";
defparam \v_cdvw_state~6 .lut_mask = 64'h3070307030703070;
defparam \v_cdvw_state~6 .shared_arith = "off";

dffeas \sig_cdvw_state.found_a_good_edge (
	.clk(clk),
	.d(\v_cdvw_state~6_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_cdvw_state.found_a_good_edge~q ),
	.prn(vcc));
defparam \sig_cdvw_state.found_a_good_edge .is_wysiwyg = "true";
defparam \sig_cdvw_state.found_a_good_edge .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~22 (
	.dataa(!\sig_cdvw_state.status.calculating~q ),
	.datab(!\sig_cdvw_state.found_a_good_edge~q ),
	.datac(!\v_cdvw_state~2_combout ),
	.datad(!\sig_cdvw_state.working_window[0]~q ),
	.datae(!\sig_cdvw_state.last_bit_value~q ),
	.dataf(!\sig_cdvw_state.window_centre_update~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~22 .extended_lut = "off";
defparam \v_cdvw_state~22 .lut_mask = 64'h10005000E0F0A0F0;
defparam \v_cdvw_state~22 .shared_arith = "off";

dffeas \sig_cdvw_state.window_centre_update (
	.clk(clk),
	.d(\v_cdvw_state~22_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_cdvw_state.window_centre_update~q ),
	.prn(vcc));
defparam \sig_cdvw_state.window_centre_update .is_wysiwyg = "true";
defparam \sig_cdvw_state.window_centre_update .power_up = "low";

arriaii_lcell_comb \sig_cdvw_state.current_window_centre[4]~4 (
	.dataa(!\sig_cdvw_state.found_a_good_edge~q ),
	.datab(!\sig_cdvw_state.last_bit_value~q ),
	.datac(!\sig_cdvw_state.window_centre_update~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_cdvw_state.current_window_centre[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_cdvw_state.current_window_centre[4]~4 .extended_lut = "off";
defparam \sig_cdvw_state.current_window_centre[4]~4 .lut_mask = 64'h8C8C8C8C8C8C8C8C;
defparam \sig_cdvw_state.current_window_centre[4]~4 .shared_arith = "off";

arriaii_lcell_comb \sig_cdvw_state.current_window_centre[4]~1 (
	.dataa(!\sig_cdvw_state.status.calculating~q ),
	.datab(!\sig_cdvw_state.working_window[0]~q ),
	.datac(!\cdvw_proc~1_combout ),
	.datad(!\cdvw_block:sig_cdvw_calc_1t~q ),
	.datae(!\Selector33~0_combout ),
	.dataf(!\sig_cdvw_state.current_window_centre[4]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_cdvw_state.current_window_centre[4]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_cdvw_state.current_window_centre[4]~1 .extended_lut = "off";
defparam \sig_cdvw_state.current_window_centre[4]~1 .lut_mask = 64'h4F4FFF4F0F0FFF0F;
defparam \sig_cdvw_state.current_window_centre[4]~1 .shared_arith = "off";

dffeas \sig_cdvw_state.current_window_centre[2] (
	.clk(clk),
	.d(\Add2~9_sumout ),
	.asdata(\sig_cdvw_state.current_bit[2]~q ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_window_centre[4]~0_combout ),
	.sload(\find_centre_of_largest_data_valid_window~2_combout ),
	.ena(\sig_cdvw_state.current_window_centre[4]~1_combout ),
	.q(\sig_cdvw_state.current_window_centre[2]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_window_centre[2] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_window_centre[2] .power_up = "low";

arriaii_lcell_comb \Add2~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sig_cdvw_state.current_window_centre[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~13_sumout ),
	.cout(\Add2~14 ),
	.shareout());
defparam \Add2~13 .extended_lut = "off";
defparam \Add2~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add2~13 .shared_arith = "off";

arriaii_lcell_comb \Add4~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sig_cdvw_state.current_bit[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~13_sumout ),
	.cout(\Add4~14 ),
	.shareout());
defparam \Add4~13 .extended_lut = "off";
defparam \Add4~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add4~13 .shared_arith = "off";

dffeas \sig_cdvw_state.current_bit[3] (
	.clk(clk),
	.d(\Add4~13_sumout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_bit[5]~2_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.current_bit[5]~0_combout ),
	.q(\sig_cdvw_state.current_bit[3]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_bit[3] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_bit[3] .power_up = "low";

dffeas \sig_cdvw_state.current_window_centre[3] (
	.clk(clk),
	.d(\Add2~13_sumout ),
	.asdata(\sig_cdvw_state.current_bit[3]~q ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_window_centre[4]~0_combout ),
	.sload(\find_centre_of_largest_data_valid_window~2_combout ),
	.ena(\sig_cdvw_state.current_window_centre[4]~1_combout ),
	.q(\sig_cdvw_state.current_window_centre[3]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_window_centre[3] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_window_centre[3] .power_up = "low";

arriaii_lcell_comb \Add2~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sig_cdvw_state.current_window_centre[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~17_sumout ),
	.cout(\Add2~18 ),
	.shareout());
defparam \Add2~17 .extended_lut = "off";
defparam \Add2~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add2~17 .shared_arith = "off";

arriaii_lcell_comb \Add4~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sig_cdvw_state.current_bit[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~17_sumout ),
	.cout(\Add4~18 ),
	.shareout());
defparam \Add4~17 .extended_lut = "off";
defparam \Add4~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add4~17 .shared_arith = "off";

dffeas \sig_cdvw_state.current_bit[4] (
	.clk(clk),
	.d(\Add4~17_sumout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_bit[5]~2_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.current_bit[5]~0_combout ),
	.q(\sig_cdvw_state.current_bit[4]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_bit[4] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_bit[4] .power_up = "low";

dffeas \sig_cdvw_state.current_window_centre[4] (
	.clk(clk),
	.d(\Add2~17_sumout ),
	.asdata(\sig_cdvw_state.current_bit[4]~q ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_window_centre[4]~0_combout ),
	.sload(\find_centre_of_largest_data_valid_window~2_combout ),
	.ena(\sig_cdvw_state.current_window_centre[4]~1_combout ),
	.q(\sig_cdvw_state.current_window_centre[4]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_window_centre[4] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_window_centre[4] .power_up = "low";

arriaii_lcell_comb \Add2~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sig_cdvw_state.current_window_centre[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~21_sumout ),
	.cout(),
	.shareout());
defparam \Add2~21 .extended_lut = "off";
defparam \Add2~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add2~21 .shared_arith = "off";

arriaii_lcell_comb \Add4~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sig_cdvw_state.current_bit[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~21_sumout ),
	.cout(),
	.shareout());
defparam \Add4~21 .extended_lut = "off";
defparam \Add4~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add4~21 .shared_arith = "off";

dffeas \sig_cdvw_state.current_bit[5] (
	.clk(clk),
	.d(\Add4~21_sumout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_bit[5]~2_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.current_bit[5]~0_combout ),
	.q(\sig_cdvw_state.current_bit[5]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_bit[5] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_bit[5] .power_up = "low";

dffeas \sig_cdvw_state.current_window_centre[5] (
	.clk(clk),
	.d(\Add2~21_sumout ),
	.asdata(\sig_cdvw_state.current_bit[5]~q ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_window_centre[4]~0_combout ),
	.sload(\find_centre_of_largest_data_valid_window~2_combout ),
	.ena(\sig_cdvw_state.current_window_centre[4]~1_combout ),
	.q(\sig_cdvw_state.current_window_centre[5]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_window_centre[5] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_window_centre[5] .power_up = "low";

arriaii_lcell_comb \sig_cdvw_state.current_window_centre[4]~2 (
	.dataa(!\sig_dgrb_state.s_track~q ),
	.datab(!\sig_cdvw_state.current_window_centre[5]~q ),
	.datac(!\sig_cdvw_state.current_window_centre[1]~q ),
	.datad(!\sig_cdvw_state.current_window_centre[2]~q ),
	.datae(!\sig_cdvw_state.current_window_centre[3]~q ),
	.dataf(!\sig_cdvw_state.current_window_centre[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_cdvw_state.current_window_centre[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_cdvw_state.current_window_centre[4]~2 .extended_lut = "off";
defparam \sig_cdvw_state.current_window_centre[4]~2 .lut_mask = 64'h1111111111111117;
defparam \sig_cdvw_state.current_window_centre[4]~2 .shared_arith = "off";

arriaii_lcell_comb \sig_cdvw_state.current_window_centre[4]~3 (
	.dataa(!\sig_dgrb_state.s_track~q ),
	.datab(!\sig_cdvw_state.current_window_centre[5]~q ),
	.datac(!\sig_cdvw_state.current_window_centre[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_cdvw_state.current_window_centre[4]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_cdvw_state.current_window_centre[4]~3 .extended_lut = "off";
defparam \sig_cdvw_state.current_window_centre[4]~3 .lut_mask = 64'hE0E0E0E0E0E0E0E0;
defparam \sig_cdvw_state.current_window_centre[4]~3 .shared_arith = "off";

arriaii_lcell_comb \sig_cdvw_state.current_window_centre[4]~0 (
	.dataa(!\find_centre_of_largest_data_valid_window~2_combout ),
	.datab(!\cdvw_proc~1_combout ),
	.datac(!\cdvw_block:sig_cdvw_calc_1t~q ),
	.datad(!\Selector33~0_combout ),
	.datae(!\sig_cdvw_state.current_window_centre[4]~2_combout ),
	.dataf(!\sig_cdvw_state.current_window_centre[4]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_cdvw_state.current_window_centre[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_cdvw_state.current_window_centre[4]~0 .extended_lut = "off";
defparam \sig_cdvw_state.current_window_centre[4]~0 .lut_mask = 64'h33F3BBFB33F333F3;
defparam \sig_cdvw_state.current_window_centre[4]~0 .shared_arith = "off";

dffeas \sig_cdvw_state.current_window_centre[0] (
	.clk(clk),
	.d(\Add2~1_sumout ),
	.asdata(\sig_cdvw_state.current_bit[0]~q ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_window_centre[4]~0_combout ),
	.sload(\find_centre_of_largest_data_valid_window~2_combout ),
	.ena(\sig_cdvw_state.current_window_centre[4]~1_combout ),
	.q(\sig_cdvw_state.current_window_centre[0]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_window_centre[0] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_window_centre[0] .power_up = "low";

dffeas \sig_cdvw_state.current_window_centre[1] (
	.clk(clk),
	.d(\Add2~5_sumout ),
	.asdata(\sig_cdvw_state.current_bit[1]~q ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_window_centre[4]~0_combout ),
	.sload(\find_centre_of_largest_data_valid_window~2_combout ),
	.ena(\sig_cdvw_state.current_window_centre[4]~1_combout ),
	.q(\sig_cdvw_state.current_window_centre[1]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_window_centre[1] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_window_centre[1] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~5 (
	.dataa(!\sig_cdvw_state.status.calculating~q ),
	.datab(!\sig_cdvw_state.working_window[0]~q ),
	.datac(!\sig_cdvw_state.last_bit_value~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~5 .extended_lut = "off";
defparam \v_cdvw_state~5 .lut_mask = 64'h1010101010101010;
defparam \v_cdvw_state~5 .shared_arith = "off";

arriaii_lcell_comb \Add3~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sig_cdvw_state.current_window_size[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~1_sumout ),
	.cout(\Add3~2 ),
	.shareout());
defparam \Add3~1 .extended_lut = "off";
defparam \Add3~1 .lut_mask = 64'h00000000000000FF;
defparam \Add3~1 .shared_arith = "off";

arriaii_lcell_comb \sig_cdvw_state.current_window_size[0]~0 (
	.dataa(!\sig_cdvw_state.working_window[0]~q ),
	.datab(!\sig_cdvw_state.last_bit_value~q ),
	.datac(!\cdvw_proc~1_combout ),
	.datad(!\cdvw_block:sig_cdvw_calc_1t~q ),
	.datae(!\Selector33~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_cdvw_state.current_window_size[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_cdvw_state.current_window_size[0]~0 .extended_lut = "off";
defparam \sig_cdvw_state.current_window_size[0]~0 .lut_mask = 64'h4F4FFF4F4F4FFF4F;
defparam \sig_cdvw_state.current_window_size[0]~0 .shared_arith = "off";

arriaii_lcell_comb \sig_cdvw_state.current_window_size[0]~2 (
	.dataa(!\sig_cdvw_state.found_a_good_edge~q ),
	.datab(!\sig_cdvw_state.working_window[0]~q ),
	.datac(!\sig_cdvw_state.last_bit_value~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_cdvw_state.current_window_size[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_cdvw_state.current_window_size[0]~2 .extended_lut = "off";
defparam \sig_cdvw_state.current_window_size[0]~2 .lut_mask = 64'h8383838383838383;
defparam \sig_cdvw_state.current_window_size[0]~2 .shared_arith = "off";

arriaii_lcell_comb \sig_cdvw_state.current_window_size[0]~1 (
	.dataa(!\sig_cdvw_state.status.calculating~q ),
	.datab(!\cdvw_proc~1_combout ),
	.datac(!\cdvw_block:sig_cdvw_calc_1t~q ),
	.datad(!\Selector33~0_combout ),
	.datae(!\sig_cdvw_state.current_window_size[0]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_cdvw_state.current_window_size[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_cdvw_state.current_window_size[0]~1 .extended_lut = "off";
defparam \sig_cdvw_state.current_window_size[0]~1 .lut_mask = 64'h77F733F377F733F3;
defparam \sig_cdvw_state.current_window_size[0]~1 .shared_arith = "off";

dffeas \sig_cdvw_state.current_window_size[0] (
	.clk(clk),
	.d(\Add3~1_sumout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_window_size[0]~0_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.current_window_size[0]~1_combout ),
	.q(\sig_cdvw_state.current_window_size[0]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_window_size[0] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_window_size[0] .power_up = "low";

arriaii_lcell_comb \Add3~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sig_cdvw_state.current_window_size[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~5_sumout ),
	.cout(\Add3~6 ),
	.shareout());
defparam \Add3~5 .extended_lut = "off";
defparam \Add3~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add3~5 .shared_arith = "off";

dffeas \sig_cdvw_state.current_window_size[1] (
	.clk(clk),
	.d(\Add3~5_sumout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_window_size[0]~0_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.current_window_size[0]~1_combout ),
	.q(\sig_cdvw_state.current_window_size[1]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_window_size[1] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_window_size[1] .power_up = "low";

arriaii_lcell_comb \Add3~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sig_cdvw_state.current_window_size[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~9_sumout ),
	.cout(\Add3~10 ),
	.shareout());
defparam \Add3~9 .extended_lut = "off";
defparam \Add3~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add3~9 .shared_arith = "off";

dffeas \sig_cdvw_state.current_window_size[2] (
	.clk(clk),
	.d(\Add3~9_sumout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_window_size[0]~0_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.current_window_size[0]~1_combout ),
	.q(\sig_cdvw_state.current_window_size[2]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_window_size[2] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_window_size[2] .power_up = "low";

arriaii_lcell_comb \Add3~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sig_cdvw_state.current_window_size[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~13_sumout ),
	.cout(\Add3~14 ),
	.shareout());
defparam \Add3~13 .extended_lut = "off";
defparam \Add3~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add3~13 .shared_arith = "off";

dffeas \sig_cdvw_state.current_window_size[3] (
	.clk(clk),
	.d(\Add3~13_sumout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_window_size[0]~0_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.current_window_size[0]~1_combout ),
	.q(\sig_cdvw_state.current_window_size[3]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_window_size[3] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_window_size[3] .power_up = "low";

dffeas \sig_cdvw_state.largest_window_size[3] (
	.clk(clk),
	.d(\sig_cdvw_state.current_window_size[3]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\v_cdvw_state~2_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.largest_window_centre[1]~0_combout ),
	.q(\sig_cdvw_state.largest_window_size[3]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.largest_window_size[3] .is_wysiwyg = "true";
defparam \sig_cdvw_state.largest_window_size[3] .power_up = "low";

arriaii_lcell_comb \Add3~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sig_cdvw_state.current_window_size[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~17_sumout ),
	.cout(\Add3~18 ),
	.shareout());
defparam \Add3~17 .extended_lut = "off";
defparam \Add3~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add3~17 .shared_arith = "off";

dffeas \sig_cdvw_state.current_window_size[4] (
	.clk(clk),
	.d(\Add3~17_sumout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_window_size[0]~0_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.current_window_size[0]~1_combout ),
	.q(\sig_cdvw_state.current_window_size[4]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_window_size[4] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_window_size[4] .power_up = "low";

arriaii_lcell_comb \Add3~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sig_cdvw_state.current_window_size[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~21_sumout ),
	.cout(),
	.shareout());
defparam \Add3~21 .extended_lut = "off";
defparam \Add3~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add3~21 .shared_arith = "off";

dffeas \sig_cdvw_state.current_window_size[5] (
	.clk(clk),
	.d(\Add3~21_sumout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_window_size[0]~0_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.current_window_size[0]~1_combout ),
	.q(\sig_cdvw_state.current_window_size[5]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_window_size[5] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_window_size[5] .power_up = "low";

dffeas \sig_cdvw_state.largest_window_size[5] (
	.clk(clk),
	.d(\sig_cdvw_state.current_window_size[5]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\v_cdvw_state~2_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.largest_window_centre[1]~0_combout ),
	.q(\sig_cdvw_state.largest_window_size[5]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.largest_window_size[5] .is_wysiwyg = "true";
defparam \sig_cdvw_state.largest_window_size[5] .power_up = "low";

arriaii_lcell_comb \LessThan3~1 (
	.dataa(!\sig_cdvw_state.largest_window_size[4]~q ),
	.datab(!\sig_cdvw_state.current_window_size[4]~q ),
	.datac(!\sig_cdvw_state.largest_window_size[5]~q ),
	.datad(!\sig_cdvw_state.current_window_size[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan3~1 .extended_lut = "off";
defparam \LessThan3~1 .lut_mask = 64'h9009900990099009;
defparam \LessThan3~1 .shared_arith = "off";

arriaii_lcell_comb \LessThan3~2 (
	.dataa(!\sig_cdvw_state.largest_window_size[4]~q ),
	.datab(!\sig_cdvw_state.current_window_size[4]~q ),
	.datac(!\sig_cdvw_state.largest_window_size[5]~q ),
	.datad(!\sig_cdvw_state.current_window_size[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan3~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan3~2 .extended_lut = "off";
defparam \LessThan3~2 .lut_mask = 64'h20F220F220F220F2;
defparam \LessThan3~2 .shared_arith = "off";

arriaii_lcell_comb \LessThan3~3 (
	.dataa(!\LessThan3~0_combout ),
	.datab(!\sig_cdvw_state.largest_window_size[3]~q ),
	.datac(!\sig_cdvw_state.current_window_size[3]~q ),
	.datad(!\LessThan3~1_combout ),
	.datae(!\LessThan3~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan3~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan3~3 .extended_lut = "off";
defparam \LessThan3~3 .lut_mask = 64'hFFB20000FFB20000;
defparam \LessThan3~3 .shared_arith = "off";

arriaii_lcell_comb \sig_cdvw_state.largest_window_centre[1]~0 (
	.dataa(!\v_cdvw_state~2_combout ),
	.datab(!\v_cdvw_state~5_combout ),
	.datac(!\LessThan3~3_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_cdvw_state.largest_window_centre[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_cdvw_state.largest_window_centre[1]~0 .extended_lut = "off";
defparam \sig_cdvw_state.largest_window_centre[1]~0 .lut_mask = 64'h7575757575757575;
defparam \sig_cdvw_state.largest_window_centre[1]~0 .shared_arith = "off";

dffeas \sig_cdvw_state.largest_window_centre[1] (
	.clk(clk),
	.d(\sig_cdvw_state.current_window_centre[1]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\v_cdvw_state~2_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.largest_window_centre[1]~0_combout ),
	.q(\sig_cdvw_state.largest_window_centre[1]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.largest_window_centre[1] .is_wysiwyg = "true";
defparam \sig_cdvw_state.largest_window_centre[1] .power_up = "low";

dffeas \sig_cdvw_state.largest_window_centre[2] (
	.clk(clk),
	.d(\sig_cdvw_state.current_window_centre[2]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\v_cdvw_state~2_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.largest_window_centre[1]~0_combout ),
	.q(\sig_cdvw_state.largest_window_centre[2]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.largest_window_centre[2] .is_wysiwyg = "true";
defparam \sig_cdvw_state.largest_window_centre[2] .power_up = "low";

arriaii_lcell_comb \rsc_block:sig_count[2]~0 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_flush_datapath~q ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datac(!\rsc_block:sig_rsc_last_state.s_rsc_test_dq~q ),
	.datad(!\rsc_block:sig_rsc_last_state.s_rsc_flush_datapath~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rsc_block:sig_count[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rsc_block:sig_count[2]~0 .extended_lut = "off";
defparam \rsc_block:sig_count[2]~0 .lut_mask = 64'h7530753075307530;
defparam \rsc_block:sig_count[2]~0 .shared_arith = "off";

arriaii_lcell_comb \Add6~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\rsc_block:sig_count[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~1_sumout ),
	.cout(\Add6~2 ),
	.shareout());
defparam \Add6~1 .extended_lut = "off";
defparam \Add6~1 .lut_mask = 64'h00000000000000FF;
defparam \Add6~1 .shared_arith = "off";

dffeas \sig_cdvw_state.largest_window_centre[0] (
	.clk(clk),
	.d(\sig_cdvw_state.current_window_centre[0]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\v_cdvw_state~2_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.largest_window_centre[1]~0_combout ),
	.q(\sig_cdvw_state.largest_window_centre[0]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.largest_window_centre[0] .is_wysiwyg = "true";
defparam \sig_cdvw_state.largest_window_centre[0] .power_up = "low";

arriaii_lcell_comb \Selector48~0 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_idle~q ),
	.datab(!\rsc_block:sig_count[2]~0_combout ),
	.datac(!\rsc_block:sig_count[6]~0_combout ),
	.datad(!\Add6~1_sumout ),
	.datae(!\sig_cdvw_state.largest_window_centre[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector48~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector48~0 .extended_lut = "off";
defparam \Selector48~0 .lut_mask = 64'h0040044400400444;
defparam \Selector48~0 .shared_arith = "off";

dffeas \sig_cdvw_state.largest_window_centre[4] (
	.clk(clk),
	.d(\sig_cdvw_state.current_window_centre[4]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\v_cdvw_state~2_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.largest_window_centre[1]~0_combout ),
	.q(\sig_cdvw_state.largest_window_centre[4]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.largest_window_centre[4] .is_wysiwyg = "true";
defparam \sig_cdvw_state.largest_window_centre[4] .power_up = "low";

dffeas \sig_cdvw_state.largest_window_centre[3] (
	.clk(clk),
	.d(\sig_cdvw_state.current_window_centre[3]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\v_cdvw_state~2_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.largest_window_centre[1]~0_combout ),
	.q(\sig_cdvw_state.largest_window_centre[3]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.largest_window_centre[3] .is_wysiwyg = "true";
defparam \sig_cdvw_state.largest_window_centre[3] .power_up = "low";

arriaii_lcell_comb \Add6~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\rsc_block:sig_count[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~9_sumout ),
	.cout(\Add6~10 ),
	.shareout());
defparam \Add6~9 .extended_lut = "off";
defparam \Add6~9 .lut_mask = 64'h00000000000000FF;
defparam \Add6~9 .shared_arith = "off";

arriaii_lcell_comb \Add6~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\rsc_block:sig_count[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~13_sumout ),
	.cout(\Add6~14 ),
	.shareout());
defparam \Add6~13 .extended_lut = "off";
defparam \Add6~13 .lut_mask = 64'h00000000000000FF;
defparam \Add6~13 .shared_arith = "off";

arriaii_lcell_comb \Selector45~0 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_idle~q ),
	.datab(!\rsc_block:sig_count[2]~0_combout ),
	.datac(!\rsc_block:sig_count[6]~0_combout ),
	.datad(!\sig_cdvw_state.largest_window_centre[3]~q ),
	.datae(!\Add6~13_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector45~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector45~0 .extended_lut = "off";
defparam \Selector45~0 .lut_mask = 64'h303F707F303F707F;
defparam \Selector45~0 .shared_arith = "off";

dffeas \rsc_block:sig_count[3] (
	.clk(clk),
	.d(\Selector45~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rsc_block:sig_count[2]~2_combout ),
	.q(\rsc_block:sig_count[3]~q ),
	.prn(vcc));
defparam \rsc_block:sig_count[3] .is_wysiwyg = "true";
defparam \rsc_block:sig_count[3] .power_up = "low";

arriaii_lcell_comb \Add6~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\rsc_block:sig_count[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~17_sumout ),
	.cout(\Add6~18 ),
	.shareout());
defparam \Add6~17 .extended_lut = "off";
defparam \Add6~17 .lut_mask = 64'h00000000000000FF;
defparam \Add6~17 .shared_arith = "off";

arriaii_lcell_comb \Selector44~0 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_flush_datapath~q ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_idle~q ),
	.datac(!\rsc_block:sig_rsc_last_state.s_rsc_flush_datapath~q ),
	.datad(!\Add6~17_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector44~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector44~0 .extended_lut = "off";
defparam \Selector44~0 .lut_mask = 64'h5073507350735073;
defparam \Selector44~0 .shared_arith = "off";

arriaii_lcell_comb \Selector44~1 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datab(!\rsc_block:sig_rsc_last_state.s_rsc_test_dq~q ),
	.datac(!\rsc_block:sig_count[6]~0_combout ),
	.datad(!\sig_cdvw_state.largest_window_centre[4]~q ),
	.datae(!\Selector44~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector44~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector44~1 .extended_lut = "off";
defparam \Selector44~1 .lut_mask = 64'h000FB0BF000FB0BF;
defparam \Selector44~1 .shared_arith = "off";

dffeas \rsc_block:sig_count[4] (
	.clk(clk),
	.d(\Selector44~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rsc_block:sig_count[2]~2_combout ),
	.q(\rsc_block:sig_count[4]~q ),
	.prn(vcc));
defparam \rsc_block:sig_count[4] .is_wysiwyg = "true";
defparam \rsc_block:sig_count[4] .power_up = "low";

arriaii_lcell_comb \Add6~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\rsc_block:sig_count[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~21_sumout ),
	.cout(\Add6~22 ),
	.shareout());
defparam \Add6~21 .extended_lut = "off";
defparam \Add6~21 .lut_mask = 64'h00000000000000FF;
defparam \Add6~21 .shared_arith = "off";

dffeas \sig_cdvw_state.largest_window_centre[5] (
	.clk(clk),
	.d(\sig_cdvw_state.current_window_centre[5]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\v_cdvw_state~2_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.largest_window_centre[1]~0_combout ),
	.q(\sig_cdvw_state.largest_window_centre[5]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.largest_window_centre[5] .is_wysiwyg = "true";
defparam \sig_cdvw_state.largest_window_centre[5] .power_up = "low";

arriaii_lcell_comb \Selector43~0 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_idle~q ),
	.datab(!\rsc_block:sig_count[2]~0_combout ),
	.datac(!\rsc_block:sig_count[6]~0_combout ),
	.datad(!\Add6~21_sumout ),
	.datae(!\sig_cdvw_state.largest_window_centre[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector43~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector43~0 .extended_lut = "off";
defparam \Selector43~0 .lut_mask = 64'h0040044400400444;
defparam \Selector43~0 .shared_arith = "off";

dffeas \rsc_block:sig_count[5] (
	.clk(clk),
	.d(\Selector43~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rsc_block:sig_count[2]~2_combout ),
	.q(\rsc_block:sig_count[5]~q ),
	.prn(vcc));
defparam \rsc_block:sig_count[5] .is_wysiwyg = "true";
defparam \rsc_block:sig_count[5] .power_up = "low";

arriaii_lcell_comb \Add6~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\rsc_block:sig_count[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~25_sumout ),
	.cout(\Add6~26 ),
	.shareout());
defparam \Add6~25 .extended_lut = "off";
defparam \Add6~25 .lut_mask = 64'h00000000000000FF;
defparam \Add6~25 .shared_arith = "off";

arriaii_lcell_comb \Selector58~1 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datab(!\rsc_block:sig_rsc_last_state.s_rsc_test_dq~q ),
	.datac(!\rsc_block:sig_rsc_last_state.s_rsc_flush_datapath~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector58~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector58~1 .extended_lut = "off";
defparam \Selector58~1 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \Selector58~1 .shared_arith = "off";

arriaii_lcell_comb \Selector42~0 (
	.dataa(!\sig_rsc_ac_access_req~0_combout ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_idle~q ),
	.datac(!\rsc_block:sig_count[6]~0_combout ),
	.datad(!\Add6~25_sumout ),
	.datae(!\Selector58~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector42~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector42~0 .extended_lut = "off";
defparam \Selector42~0 .lut_mask = 64'h0020003000200030;
defparam \Selector42~0 .shared_arith = "off";

arriaii_lcell_comb \rsc_block:sig_count[2]~3 (
	.dataa(!\rsc_block:sig_count[0]~q ),
	.datab(!\rsc_block:sig_count[7]~q ),
	.datac(!\rsc_block:sig_count[6]~q ),
	.datad(!\rsc_block:sig_count[1]~q ),
	.datae(!\rsc_block:sig_count[2]~q ),
	.dataf(!\rsc_block:sig_count[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rsc_block:sig_count[2]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rsc_block:sig_count[2]~3 .extended_lut = "off";
defparam \rsc_block:sig_count[2]~3 .lut_mask = 64'h8000000000000000;
defparam \rsc_block:sig_count[2]~3 .shared_arith = "off";

arriaii_lcell_comb \rsc_block:sig_count[2]~4 (
	.dataa(!\rsc_block:sig_rsc_last_state.s_rsc_seek_cdvw~q ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_seek_cdvw~q ),
	.datac(!\rsc_block:sig_rsc_state.s_rsc_flush_datapath~q ),
	.datad(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datae(!\rsc_block:sig_rsc_state.s_rsc_idle~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rsc_block:sig_count[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rsc_block:sig_count[2]~4 .extended_lut = "off";
defparam \rsc_block:sig_count[2]~4 .lut_mask = 64'h1111D1111111D111;
defparam \rsc_block:sig_count[2]~4 .shared_arith = "off";

arriaii_lcell_comb \rsc_block:sig_count[2]~1 (
	.dataa(!\sig_phs_shft_end~q ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_seek_cdvw~q ),
	.datac(!\rsc_block:sig_count[4]~q ),
	.datad(!\rsc_block:sig_count[5]~q ),
	.datae(!\rsc_block:sig_count[2]~3_combout ),
	.dataf(!\rsc_block:sig_count[2]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rsc_block:sig_count[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rsc_block:sig_count[2]~1 .extended_lut = "off";
defparam \rsc_block:sig_count[2]~1 .lut_mask = 64'h00000000EEEEFEEE;
defparam \rsc_block:sig_count[2]~1 .shared_arith = "off";

arriaii_lcell_comb \rsc_block:sig_count[6]~2 (
	.dataa(!\sig_rsc_ac_access_req~0_combout ),
	.datab(!\rsc_block:sig_count[6]~1_combout ),
	.datac(!\rsc_block:sig_count[2]~1_combout ),
	.datad(!\Selector58~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rsc_block:sig_count[6]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rsc_block:sig_count[6]~2 .extended_lut = "off";
defparam \rsc_block:sig_count[6]~2 .lut_mask = 64'hF0B0F0B0F0B0F0B0;
defparam \rsc_block:sig_count[6]~2 .shared_arith = "off";

dffeas \rsc_block:sig_count[6] (
	.clk(clk),
	.d(\Selector42~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rsc_block:sig_count[6]~2_combout ),
	.q(\rsc_block:sig_count[6]~q ),
	.prn(vcc));
defparam \rsc_block:sig_count[6] .is_wysiwyg = "true";
defparam \rsc_block:sig_count[6] .power_up = "low";

arriaii_lcell_comb \Add6~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\rsc_block:sig_count[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~29_sumout ),
	.cout(),
	.shareout());
defparam \Add6~29 .extended_lut = "off";
defparam \Add6~29 .lut_mask = 64'h00000000000000FF;
defparam \Add6~29 .shared_arith = "off";

arriaii_lcell_comb \Selector41~0 (
	.dataa(!\sig_rsc_ac_access_req~0_combout ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_idle~q ),
	.datac(!\rsc_block:sig_count[6]~0_combout ),
	.datad(!\Add6~29_sumout ),
	.datae(!\Selector58~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector41~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector41~0 .extended_lut = "off";
defparam \Selector41~0 .lut_mask = 64'h0020003000200030;
defparam \Selector41~0 .shared_arith = "off";

dffeas \rsc_block:sig_count[7] (
	.clk(clk),
	.d(\Selector41~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rsc_block:sig_count[6]~2_combout ),
	.q(\rsc_block:sig_count[7]~q ),
	.prn(vcc));
defparam \rsc_block:sig_count[7] .is_wysiwyg = "true";
defparam \rsc_block:sig_count[7] .power_up = "low";

arriaii_lcell_comb \Equal14~0 (
	.dataa(!\rsc_block:sig_count[4]~q ),
	.datab(!\rsc_block:sig_count[5]~q ),
	.datac(!\rsc_block:sig_count[7]~q ),
	.datad(!\rsc_block:sig_count[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal14~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal14~0 .extended_lut = "off";
defparam \Equal14~0 .lut_mask = 64'h8000800080008000;
defparam \Equal14~0 .shared_arith = "off";

dffeas \rsc_block:sig_curr_byte_ln_dis (
	.clk(clk),
	.d(sig_addr_cmd0cke0),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_curr_byte_ln_dis~q ),
	.prn(vcc));
defparam \rsc_block:sig_curr_byte_ln_dis .is_wysiwyg = "true";
defparam \rsc_block:sig_curr_byte_ln_dis .power_up = "low";

arriaii_lcell_comb \Add7~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sig_dq_pin_ctr[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~5_sumout ),
	.cout(\Add7~6 ),
	.shareout());
defparam \Add7~5 .extended_lut = "off";
defparam \Add7~5 .lut_mask = 64'h00000000000000FF;
defparam \Add7~5 .shared_arith = "off";

arriaii_lcell_comb \Add7~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sig_dq_pin_ctr[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~9_sumout ),
	.cout(\Add7~10 ),
	.shareout());
defparam \Add7~9 .extended_lut = "off";
defparam \Add7~9 .lut_mask = 64'h00000000000000FF;
defparam \Add7~9 .shared_arith = "off";

arriaii_lcell_comb \sig_dq_pin_ctr[0]~1 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datab(!\rsc_block:sig_chkd_all_dq_pins~q ),
	.datac(!\Selector53~0_combout ),
	.datad(!\rsc_block:sig_rsc_state.s_rsc_idle~q ),
	.datae(!\rsc_block:sig_rsc_state.s_rsc_test_phase~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dq_pin_ctr[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dq_pin_ctr[0]~1 .extended_lut = "off";
defparam \sig_dq_pin_ctr[0]~1 .lut_mask = 64'hAE04AEAEAE04AEAE;
defparam \sig_dq_pin_ctr[0]~1 .shared_arith = "off";

dffeas \sig_dq_pin_ctr[2] (
	.clk(clk),
	.d(\Add7~9_sumout ),
	.asdata(\single_bit_cal~_wirecell_combout ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_dq_pin_ctr[0]~0_combout ),
	.sload(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.ena(\sig_dq_pin_ctr[0]~1_combout ),
	.q(\sig_dq_pin_ctr[2]~q ),
	.prn(vcc));
defparam \sig_dq_pin_ctr[2] .is_wysiwyg = "true";
defparam \sig_dq_pin_ctr[2] .power_up = "low";

arriaii_lcell_comb \tp_match_block:sig_rdata_current_pin[15]~0 (
	.dataa(!\sig_dq_pin_ctr[1]~q ),
	.datab(!\sig_dq_pin_ctr[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\tp_match_block:sig_rdata_current_pin[15]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \tp_match_block:sig_rdata_current_pin[15]~0 .extended_lut = "off";
defparam \tp_match_block:sig_rdata_current_pin[15]~0 .lut_mask = 64'h4444444444444444;
defparam \tp_match_block:sig_rdata_current_pin[15]~0 .shared_arith = "off";

arriaii_lcell_comb \Add7~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sig_dq_pin_ctr[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~13_sumout ),
	.cout(\Add7~14 ),
	.shareout());
defparam \Add7~13 .extended_lut = "off";
defparam \Add7~13 .lut_mask = 64'h00000000000000FF;
defparam \Add7~13 .shared_arith = "off";

dffeas \sig_dq_pin_ctr[3] (
	.clk(clk),
	.d(\Add7~13_sumout ),
	.asdata(\single_bit_cal~_wirecell_combout ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_dq_pin_ctr[0]~0_combout ),
	.sload(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.ena(\sig_dq_pin_ctr[0]~1_combout ),
	.q(\sig_dq_pin_ctr[3]~q ),
	.prn(vcc));
defparam \sig_dq_pin_ctr[3] .is_wysiwyg = "true";
defparam \sig_dq_pin_ctr[3] .power_up = "low";

arriaii_lcell_comb \Add7~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\sig_dq_pin_ctr[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add7~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add7~17_sumout ),
	.cout(),
	.shareout());
defparam \Add7~17 .extended_lut = "off";
defparam \Add7~17 .lut_mask = 64'h00000000000000FF;
defparam \Add7~17 .shared_arith = "off";

dffeas \sig_dq_pin_ctr[4] (
	.clk(clk),
	.d(\Add7~17_sumout ),
	.asdata(\single_bit_cal~_wirecell_combout ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_dq_pin_ctr[0]~0_combout ),
	.sload(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.ena(\sig_dq_pin_ctr[0]~1_combout ),
	.q(\sig_dq_pin_ctr[4]~q ),
	.prn(vcc));
defparam \sig_dq_pin_ctr[4] .is_wysiwyg = "true";
defparam \sig_dq_pin_ctr[4] .power_up = "low";

arriaii_lcell_comb \Mux7~0 (
	.dataa(!q_b_66),
	.datab(!q_b_98),
	.datac(!q_b_82),
	.datad(!q_b_114),
	.datae(!\sig_dq_pin_ctr[4]~q ),
	.dataf(!\sig_dq_pin_ctr[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux7~0 .extended_lut = "off";
defparam \Mux7~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux7~0 .shared_arith = "off";

arriaii_lcell_comb \Mux7~2 (
	.dataa(!q_b_97),
	.datab(!q_b_101),
	.datac(!q_b_99),
	.datad(!q_b_103),
	.datae(!\sig_dq_pin_ctr[2]~q ),
	.dataf(!\sig_dq_pin_ctr[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux7~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux7~2 .extended_lut = "off";
defparam \Mux7~2 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux7~2 .shared_arith = "off";

arriaii_lcell_comb \Mux7~3 (
	.dataa(!q_b_81),
	.datab(!q_b_85),
	.datac(!q_b_83),
	.datad(!q_b_87),
	.datae(!\sig_dq_pin_ctr[2]~q ),
	.dataf(!\sig_dq_pin_ctr[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux7~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux7~3 .extended_lut = "off";
defparam \Mux7~3 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux7~3 .shared_arith = "off";

arriaii_lcell_comb \Mux7~4 (
	.dataa(!q_b_113),
	.datab(!q_b_117),
	.datac(!q_b_115),
	.datad(!q_b_119),
	.datae(!\sig_dq_pin_ctr[2]~q ),
	.dataf(!\sig_dq_pin_ctr[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux7~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux7~4 .extended_lut = "off";
defparam \Mux7~4 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux7~4 .shared_arith = "off";

arriaii_lcell_comb \Mux7~5 (
	.dataa(!\Mux7~1_combout ),
	.datab(!\Mux7~2_combout ),
	.datac(!\Mux7~3_combout ),
	.datad(!\Mux7~4_combout ),
	.datae(!\sig_dq_pin_ctr[4]~q ),
	.dataf(!\sig_dq_pin_ctr[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux7~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux7~5 .extended_lut = "off";
defparam \Mux7~5 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux7~5 .shared_arith = "off";

arriaii_lcell_comb \Mux7~6 (
	.dataa(!q_b_70),
	.datab(!q_b_102),
	.datac(!q_b_86),
	.datad(!q_b_118),
	.datae(!\sig_dq_pin_ctr[4]~q ),
	.dataf(!\sig_dq_pin_ctr[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux7~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux7~6 .extended_lut = "off";
defparam \Mux7~6 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux7~6 .shared_arith = "off";

arriaii_lcell_comb \Mux7~7 (
	.dataa(!q_b_68),
	.datab(!q_b_100),
	.datac(!q_b_84),
	.datad(!q_b_116),
	.datae(!\sig_dq_pin_ctr[4]~q ),
	.dataf(!\sig_dq_pin_ctr[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux7~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux7~7 .extended_lut = "off";
defparam \Mux7~7 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux7~7 .shared_arith = "off";

arriaii_lcell_comb \Mux7~8 (
	.dataa(!q_b_64),
	.datab(!q_b_96),
	.datac(!q_b_80),
	.datad(!q_b_112),
	.datae(!\sig_dq_pin_ctr[4]~q ),
	.dataf(!\sig_dq_pin_ctr[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux7~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux7~8 .extended_lut = "off";
defparam \Mux7~8 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux7~8 .shared_arith = "off";

arriaii_lcell_comb \Mux7~9 (
	.dataa(!\sig_dq_pin_ctr[1]~q ),
	.datab(!\sig_dq_pin_ctr[2]~q ),
	.datac(!\Mux7~6_combout ),
	.datad(!\Mux7~7_combout ),
	.datae(!\Mux7~8_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux7~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux7~9 .extended_lut = "off";
defparam \Mux7~9 .lut_mask = 64'h05278DAF05278DAF;
defparam \Mux7~9 .shared_arith = "off";

arriaii_lcell_comb \Mux7~10 (
	.dataa(!\sig_dq_pin_ctr[0]~q ),
	.datab(!\tp_match_block:sig_rdata_current_pin[15]~0_combout ),
	.datac(!\Mux7~0_combout ),
	.datad(!\Mux7~5_combout ),
	.datae(!\Mux7~9_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux7~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux7~10 .extended_lut = "off";
defparam \Mux7~10 .lut_mask = 64'h02578ADF02578ADF;
defparam \Mux7~10 .shared_arith = "off";

dffeas \tp_match_block:sig_rdata_current_pin[14] (
	.clk(clk),
	.d(\Mux7~10_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_current_pin[14]~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_current_pin[14] .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_current_pin[14] .power_up = "low";

dffeas \tp_match_block:sig_rdata_current_pin[10] (
	.clk(clk),
	.d(\tp_match_block:sig_rdata_current_pin[14]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_current_pin[10]~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_current_pin[10] .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_current_pin[10] .power_up = "low";

dffeas \tp_match_block:sig_rdata_current_pin[6] (
	.clk(clk),
	.d(\tp_match_block:sig_rdata_current_pin[10]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_current_pin[6]~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_current_pin[6] .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_current_pin[6] .power_up = "low";

arriaii_lcell_comb \Mux8~0 (
	.dataa(!q_b_74),
	.datab(!q_b_106),
	.datac(!q_b_90),
	.datad(!q_b_122),
	.datae(!\sig_dq_pin_ctr[4]~q ),
	.dataf(!\sig_dq_pin_ctr[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux8~0 .extended_lut = "off";
defparam \Mux8~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux8~0 .shared_arith = "off";

arriaii_lcell_comb \Mux8~2 (
	.dataa(!q_b_105),
	.datab(!q_b_109),
	.datac(!q_b_107),
	.datad(!q_b_111),
	.datae(!\sig_dq_pin_ctr[2]~q ),
	.dataf(!\sig_dq_pin_ctr[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux8~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux8~2 .extended_lut = "off";
defparam \Mux8~2 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux8~2 .shared_arith = "off";

arriaii_lcell_comb \Mux8~3 (
	.dataa(!q_b_89),
	.datab(!q_b_93),
	.datac(!q_b_91),
	.datad(!q_b_95),
	.datae(!\sig_dq_pin_ctr[2]~q ),
	.dataf(!\sig_dq_pin_ctr[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux8~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux8~3 .extended_lut = "off";
defparam \Mux8~3 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux8~3 .shared_arith = "off";

arriaii_lcell_comb \Mux8~4 (
	.dataa(!q_b_121),
	.datab(!q_b_125),
	.datac(!q_b_123),
	.datad(!q_b_127),
	.datae(!\sig_dq_pin_ctr[2]~q ),
	.dataf(!\sig_dq_pin_ctr[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux8~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux8~4 .extended_lut = "off";
defparam \Mux8~4 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux8~4 .shared_arith = "off";

arriaii_lcell_comb \Mux8~5 (
	.dataa(!\Mux8~1_combout ),
	.datab(!\Mux8~2_combout ),
	.datac(!\Mux8~3_combout ),
	.datad(!\Mux8~4_combout ),
	.datae(!\sig_dq_pin_ctr[4]~q ),
	.dataf(!\sig_dq_pin_ctr[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux8~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux8~5 .extended_lut = "off";
defparam \Mux8~5 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux8~5 .shared_arith = "off";

arriaii_lcell_comb \Mux8~6 (
	.dataa(!q_b_78),
	.datab(!q_b_110),
	.datac(!q_b_94),
	.datad(!q_b_126),
	.datae(!\sig_dq_pin_ctr[4]~q ),
	.dataf(!\sig_dq_pin_ctr[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux8~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux8~6 .extended_lut = "off";
defparam \Mux8~6 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux8~6 .shared_arith = "off";

arriaii_lcell_comb \Mux8~7 (
	.dataa(!q_b_76),
	.datab(!q_b_108),
	.datac(!q_b_92),
	.datad(!q_b_124),
	.datae(!\sig_dq_pin_ctr[4]~q ),
	.dataf(!\sig_dq_pin_ctr[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux8~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux8~7 .extended_lut = "off";
defparam \Mux8~7 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux8~7 .shared_arith = "off";

arriaii_lcell_comb \Mux8~8 (
	.dataa(!q_b_72),
	.datab(!q_b_104),
	.datac(!q_b_88),
	.datad(!q_b_120),
	.datae(!\sig_dq_pin_ctr[4]~q ),
	.dataf(!\sig_dq_pin_ctr[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux8~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux8~8 .extended_lut = "off";
defparam \Mux8~8 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux8~8 .shared_arith = "off";

arriaii_lcell_comb \Mux8~9 (
	.dataa(!\sig_dq_pin_ctr[1]~q ),
	.datab(!\sig_dq_pin_ctr[2]~q ),
	.datac(!\Mux8~6_combout ),
	.datad(!\Mux8~7_combout ),
	.datae(!\Mux8~8_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux8~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux8~9 .extended_lut = "off";
defparam \Mux8~9 .lut_mask = 64'h05278DAF05278DAF;
defparam \Mux8~9 .shared_arith = "off";

arriaii_lcell_comb \Mux8~10 (
	.dataa(!\sig_dq_pin_ctr[0]~q ),
	.datab(!\tp_match_block:sig_rdata_current_pin[15]~0_combout ),
	.datac(!\Mux8~0_combout ),
	.datad(!\Mux8~5_combout ),
	.datae(!\Mux8~9_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux8~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux8~10 .extended_lut = "off";
defparam \Mux8~10 .lut_mask = 64'h02578ADF02578ADF;
defparam \Mux8~10 .shared_arith = "off";

dffeas \tp_match_block:sig_rdata_current_pin[15] (
	.clk(clk),
	.d(\Mux8~10_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_current_pin[15]~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_current_pin[15] .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_current_pin[15] .power_up = "low";

dffeas \tp_match_block:sig_rdata_current_pin[11] (
	.clk(clk),
	.d(\tp_match_block:sig_rdata_current_pin[15]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_current_pin[11]~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_current_pin[11] .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_current_pin[11] .power_up = "low";

arriaii_lcell_comb \Equal15~1 (
	.dataa(!\tp_match_block:sig_rdata_current_pin[7]~q ),
	.datab(!\tp_match_block:sig_rdata_current_pin[10]~q ),
	.datac(!\tp_match_block:sig_rdata_current_pin[11]~q ),
	.datad(!\tp_match_block:sig_rdata_current_pin[15]~q ),
	.datae(!\tp_match_block:sig_rdata_current_pin[14]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal15~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal15~1 .extended_lut = "off";
defparam \Equal15~1 .lut_mask = 64'h4000000040000000;
defparam \Equal15~1 .shared_arith = "off";

arriaii_lcell_comb \Mux5~0 (
	.dataa(!q_b_2),
	.datab(!q_b_34),
	.datac(!q_b_18),
	.datad(!q_b_50),
	.datae(!\sig_dq_pin_ctr[4]~q ),
	.dataf(!\sig_dq_pin_ctr[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux5~0 .extended_lut = "off";
defparam \Mux5~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux5~0 .shared_arith = "off";

arriaii_lcell_comb \Mux5~2 (
	.dataa(!q_b_33),
	.datab(!q_b_37),
	.datac(!q_b_35),
	.datad(!q_b_39),
	.datae(!\sig_dq_pin_ctr[2]~q ),
	.dataf(!\sig_dq_pin_ctr[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux5~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux5~2 .extended_lut = "off";
defparam \Mux5~2 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux5~2 .shared_arith = "off";

arriaii_lcell_comb \Mux5~3 (
	.dataa(!q_b_17),
	.datab(!q_b_21),
	.datac(!q_b_19),
	.datad(!q_b_23),
	.datae(!\sig_dq_pin_ctr[2]~q ),
	.dataf(!\sig_dq_pin_ctr[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux5~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux5~3 .extended_lut = "off";
defparam \Mux5~3 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux5~3 .shared_arith = "off";

arriaii_lcell_comb \Mux5~4 (
	.dataa(!q_b_49),
	.datab(!q_b_53),
	.datac(!q_b_51),
	.datad(!q_b_55),
	.datae(!\sig_dq_pin_ctr[2]~q ),
	.dataf(!\sig_dq_pin_ctr[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux5~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux5~4 .extended_lut = "off";
defparam \Mux5~4 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux5~4 .shared_arith = "off";

arriaii_lcell_comb \Mux5~5 (
	.dataa(!\Mux5~1_combout ),
	.datab(!\Mux5~2_combout ),
	.datac(!\Mux5~3_combout ),
	.datad(!\Mux5~4_combout ),
	.datae(!\sig_dq_pin_ctr[4]~q ),
	.dataf(!\sig_dq_pin_ctr[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux5~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux5~5 .extended_lut = "off";
defparam \Mux5~5 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux5~5 .shared_arith = "off";

arriaii_lcell_comb \Mux5~6 (
	.dataa(!q_b_6),
	.datab(!q_b_38),
	.datac(!q_b_22),
	.datad(!q_b_54),
	.datae(!\sig_dq_pin_ctr[4]~q ),
	.dataf(!\sig_dq_pin_ctr[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux5~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux5~6 .extended_lut = "off";
defparam \Mux5~6 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux5~6 .shared_arith = "off";

arriaii_lcell_comb \Mux5~7 (
	.dataa(!q_b_4),
	.datab(!q_b_36),
	.datac(!q_b_20),
	.datad(!q_b_52),
	.datae(!\sig_dq_pin_ctr[4]~q ),
	.dataf(!\sig_dq_pin_ctr[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux5~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux5~7 .extended_lut = "off";
defparam \Mux5~7 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux5~7 .shared_arith = "off";

arriaii_lcell_comb \Mux5~8 (
	.dataa(!q_b_0),
	.datab(!q_b_32),
	.datac(!q_b_16),
	.datad(!q_b_48),
	.datae(!\sig_dq_pin_ctr[4]~q ),
	.dataf(!\sig_dq_pin_ctr[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux5~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux5~8 .extended_lut = "off";
defparam \Mux5~8 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux5~8 .shared_arith = "off";

arriaii_lcell_comb \Mux5~9 (
	.dataa(!\sig_dq_pin_ctr[1]~q ),
	.datab(!\sig_dq_pin_ctr[2]~q ),
	.datac(!\Mux5~6_combout ),
	.datad(!\Mux5~7_combout ),
	.datae(!\Mux5~8_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux5~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux5~9 .extended_lut = "off";
defparam \Mux5~9 .lut_mask = 64'h05278DAF05278DAF;
defparam \Mux5~9 .shared_arith = "off";

arriaii_lcell_comb \Mux5~10 (
	.dataa(!\sig_dq_pin_ctr[0]~q ),
	.datab(!\tp_match_block:sig_rdata_current_pin[15]~0_combout ),
	.datac(!\Mux5~0_combout ),
	.datad(!\Mux5~5_combout ),
	.datae(!\Mux5~9_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux5~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux5~10 .extended_lut = "off";
defparam \Mux5~10 .lut_mask = 64'h02578ADF02578ADF;
defparam \Mux5~10 .shared_arith = "off";

dffeas \tp_match_block:sig_rdata_current_pin[12] (
	.clk(clk),
	.d(\Mux5~10_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_current_pin[12]~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_current_pin[12] .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_current_pin[12] .power_up = "low";

dffeas \tp_match_block:sig_rdata_current_pin[8] (
	.clk(clk),
	.d(\tp_match_block:sig_rdata_current_pin[12]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_current_pin[8]~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_current_pin[8] .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_current_pin[8] .power_up = "low";

dffeas \tp_match_block:sig_rdata_current_pin[4] (
	.clk(clk),
	.d(\tp_match_block:sig_rdata_current_pin[8]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_current_pin[4]~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_current_pin[4] .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_current_pin[4] .power_up = "low";

dffeas \tp_match_block:sig_rdata_current_pin[0] (
	.clk(clk),
	.d(\tp_match_block:sig_rdata_current_pin[4]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_current_pin[0]~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_current_pin[0] .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_current_pin[0] .power_up = "low";

dffeas \tp_match_block:sig_rdata_current_pin[2] (
	.clk(clk),
	.d(\tp_match_block:sig_rdata_current_pin[6]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_current_pin[2]~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_current_pin[2] .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_current_pin[2] .power_up = "low";

dffeas \tp_match_block:sig_rdata_current_pin[7] (
	.clk(clk),
	.d(\tp_match_block:sig_rdata_current_pin[11]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_current_pin[7]~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_current_pin[7] .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_current_pin[7] .power_up = "low";

dffeas \tp_match_block:sig_rdata_current_pin[3] (
	.clk(clk),
	.d(\tp_match_block:sig_rdata_current_pin[7]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_current_pin[3]~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_current_pin[3] .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_current_pin[3] .power_up = "low";

arriaii_lcell_comb \Mux6~0 (
	.dataa(!q_b_10),
	.datab(!q_b_42),
	.datac(!q_b_26),
	.datad(!q_b_58),
	.datae(!\sig_dq_pin_ctr[4]~q ),
	.dataf(!\sig_dq_pin_ctr[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux6~0 .extended_lut = "off";
defparam \Mux6~0 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux6~0 .shared_arith = "off";

arriaii_lcell_comb \Mux6~2 (
	.dataa(!q_b_41),
	.datab(!q_b_45),
	.datac(!q_b_43),
	.datad(!q_b_47),
	.datae(!\sig_dq_pin_ctr[2]~q ),
	.dataf(!\sig_dq_pin_ctr[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux6~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux6~2 .extended_lut = "off";
defparam \Mux6~2 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux6~2 .shared_arith = "off";

arriaii_lcell_comb \Mux6~3 (
	.dataa(!q_b_25),
	.datab(!q_b_29),
	.datac(!q_b_27),
	.datad(!q_b_31),
	.datae(!\sig_dq_pin_ctr[2]~q ),
	.dataf(!\sig_dq_pin_ctr[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux6~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux6~3 .extended_lut = "off";
defparam \Mux6~3 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux6~3 .shared_arith = "off";

arriaii_lcell_comb \Mux6~4 (
	.dataa(!q_b_57),
	.datab(!q_b_61),
	.datac(!q_b_59),
	.datad(!q_b_63),
	.datae(!\sig_dq_pin_ctr[2]~q ),
	.dataf(!\sig_dq_pin_ctr[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux6~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux6~4 .extended_lut = "off";
defparam \Mux6~4 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux6~4 .shared_arith = "off";

arriaii_lcell_comb \Mux6~5 (
	.dataa(!\Mux6~1_combout ),
	.datab(!\Mux6~2_combout ),
	.datac(!\Mux6~3_combout ),
	.datad(!\Mux6~4_combout ),
	.datae(!\sig_dq_pin_ctr[4]~q ),
	.dataf(!\sig_dq_pin_ctr[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux6~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux6~5 .extended_lut = "off";
defparam \Mux6~5 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux6~5 .shared_arith = "off";

arriaii_lcell_comb \Mux6~6 (
	.dataa(!q_b_14),
	.datab(!q_b_46),
	.datac(!q_b_30),
	.datad(!q_b_62),
	.datae(!\sig_dq_pin_ctr[4]~q ),
	.dataf(!\sig_dq_pin_ctr[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux6~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux6~6 .extended_lut = "off";
defparam \Mux6~6 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux6~6 .shared_arith = "off";

arriaii_lcell_comb \Mux6~7 (
	.dataa(!q_b_12),
	.datab(!q_b_44),
	.datac(!q_b_28),
	.datad(!q_b_60),
	.datae(!\sig_dq_pin_ctr[4]~q ),
	.dataf(!\sig_dq_pin_ctr[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux6~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux6~7 .extended_lut = "off";
defparam \Mux6~7 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux6~7 .shared_arith = "off";

arriaii_lcell_comb \Mux6~8 (
	.dataa(!q_b_8),
	.datab(!q_b_40),
	.datac(!q_b_24),
	.datad(!q_b_56),
	.datae(!\sig_dq_pin_ctr[4]~q ),
	.dataf(!\sig_dq_pin_ctr[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux6~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux6~8 .extended_lut = "off";
defparam \Mux6~8 .lut_mask = 64'h555533330F0F00FF;
defparam \Mux6~8 .shared_arith = "off";

arriaii_lcell_comb \Mux6~9 (
	.dataa(!\sig_dq_pin_ctr[1]~q ),
	.datab(!\sig_dq_pin_ctr[2]~q ),
	.datac(!\Mux6~6_combout ),
	.datad(!\Mux6~7_combout ),
	.datae(!\Mux6~8_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux6~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux6~9 .extended_lut = "off";
defparam \Mux6~9 .lut_mask = 64'h05278DAF05278DAF;
defparam \Mux6~9 .shared_arith = "off";

arriaii_lcell_comb \Mux6~10 (
	.dataa(!\sig_dq_pin_ctr[0]~q ),
	.datab(!\Mux6~0_combout ),
	.datac(!\tp_match_block:sig_rdata_current_pin[15]~0_combout ),
	.datad(!\Mux6~5_combout ),
	.datae(!\Mux6~9_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux6~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux6~10 .extended_lut = "off";
defparam \Mux6~10 .lut_mask = 64'h0257A2F70257A2F7;
defparam \Mux6~10 .shared_arith = "off";

dffeas \tp_match_block:sig_rdata_current_pin[13] (
	.clk(clk),
	.d(\Mux6~10_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_current_pin[13]~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_current_pin[13] .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_current_pin[13] .power_up = "low";

dffeas \tp_match_block:sig_rdata_current_pin[9] (
	.clk(clk),
	.d(\tp_match_block:sig_rdata_current_pin[13]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_current_pin[9]~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_current_pin[9] .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_current_pin[9] .power_up = "low";

dffeas \tp_match_block:sig_rdata_current_pin[5] (
	.clk(clk),
	.d(\tp_match_block:sig_rdata_current_pin[9]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_current_pin[5]~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_current_pin[5] .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_current_pin[5] .power_up = "low";

arriaii_lcell_comb \Equal15~2 (
	.dataa(!\tp_match_block:sig_rdata_current_pin[1]~q ),
	.datab(!\tp_match_block:sig_rdata_current_pin[2]~q ),
	.datac(!\tp_match_block:sig_rdata_current_pin[3]~q ),
	.datad(!\tp_match_block:sig_rdata_current_pin[5]~q ),
	.datae(!\tp_match_block:sig_rdata_current_pin[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal15~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal15~2 .extended_lut = "off";
defparam \Equal15~2 .lut_mask = 64'h0000002000000020;
defparam \Equal15~2 .shared_arith = "off";

arriaii_lcell_comb \Equal15~3 (
	.dataa(!\Equal15~0_combout ),
	.datab(!\tp_match_block:sig_rdata_current_pin[6]~q ),
	.datac(!\Equal15~1_combout ),
	.datad(!\tp_match_block:sig_rdata_current_pin[0]~q ),
	.datae(!\Equal15~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal15~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal15~3 .extended_lut = "off";
defparam \Equal15~3 .lut_mask = 64'h0000000100000001;
defparam \Equal15~3 .shared_arith = "off";

dffeas sig_mtp_match(
	.clk(clk),
	.d(\Equal15~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_mtp_match~q ),
	.prn(vcc));
defparam sig_mtp_match.is_wysiwyg = "true";
defparam sig_mtp_match.power_up = "low";

arriaii_lcell_comb \rsc_block:sig_count[6]~3 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datab(!\rsc_block:sig_test_dq_expired~q ),
	.datac(!\rsc_block:sig_curr_byte_ln_dis~q ),
	.datad(!\sig_mtp_match~q ),
	.datae(!\rsc_block:sig_count[2]~q ),
	.dataf(!\rsc_block:sig_count[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rsc_block:sig_count[6]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rsc_block:sig_count[6]~3 .extended_lut = "off";
defparam \rsc_block:sig_count[6]~3 .lut_mask = 64'h0400AEAAAEAAAEAA;
defparam \rsc_block:sig_count[6]~3 .shared_arith = "off";

arriaii_lcell_comb \rsc_block:sig_count[6]~1 (
	.dataa(!\sig_dimm_driving_dq~q ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datac(!\rsc_block:sig_count[0]~q ),
	.datad(!\rsc_block:sig_count[1]~q ),
	.datae(!\Equal14~0_combout ),
	.dataf(!\rsc_block:sig_count[6]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rsc_block:sig_count[6]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rsc_block:sig_count[6]~1 .extended_lut = "off";
defparam \rsc_block:sig_count[6]~1 .lut_mask = 64'h88880888AAAAAAAA;
defparam \rsc_block:sig_count[6]~1 .shared_arith = "off";

arriaii_lcell_comb \rsc_block:sig_count[2]~2 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_flush_datapath~q ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datac(!\rsc_block:sig_rsc_last_state.s_rsc_test_dq~q ),
	.datad(!\rsc_block:sig_rsc_last_state.s_rsc_flush_datapath~q ),
	.datae(!\rsc_block:sig_count[6]~1_combout ),
	.dataf(!\rsc_block:sig_count[2]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rsc_block:sig_count[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rsc_block:sig_count[2]~2 .extended_lut = "off";
defparam \rsc_block:sig_count[2]~2 .lut_mask = 64'hFCA8FFFF00000000;
defparam \rsc_block:sig_count[2]~2 .shared_arith = "off";

dffeas \rsc_block:sig_count[0] (
	.clk(clk),
	.d(\Selector48~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rsc_block:sig_count[2]~2_combout ),
	.q(\rsc_block:sig_count[0]~q ),
	.prn(vcc));
defparam \rsc_block:sig_count[0] .is_wysiwyg = "true";
defparam \rsc_block:sig_count[0] .power_up = "low";

arriaii_lcell_comb \Add6~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\rsc_block:sig_count[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~5_sumout ),
	.cout(\Add6~6 ),
	.shareout());
defparam \Add6~5 .extended_lut = "off";
defparam \Add6~5 .lut_mask = 64'h00000000000000FF;
defparam \Add6~5 .shared_arith = "off";

arriaii_lcell_comb \Selector46~0 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_flush_datapath~q ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_idle~q ),
	.datac(!\rsc_block:sig_rsc_last_state.s_rsc_flush_datapath~q ),
	.datad(!\Add6~9_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector46~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector46~0 .extended_lut = "off";
defparam \Selector46~0 .lut_mask = 64'h5073507350735073;
defparam \Selector46~0 .shared_arith = "off";

arriaii_lcell_comb \Selector46~1 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datab(!\rsc_block:sig_rsc_last_state.s_rsc_test_dq~q ),
	.datac(!\rsc_block:sig_count[6]~0_combout ),
	.datad(!\sig_cdvw_state.largest_window_centre[2]~q ),
	.datae(!\Selector46~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector46~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector46~1 .extended_lut = "off";
defparam \Selector46~1 .lut_mask = 64'h000FB0BF000FB0BF;
defparam \Selector46~1 .shared_arith = "off";

dffeas \rsc_block:sig_count[2] (
	.clk(clk),
	.d(\Selector46~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rsc_block:sig_count[2]~2_combout ),
	.q(\rsc_block:sig_count[2]~q ),
	.prn(vcc));
defparam \rsc_block:sig_count[2] .is_wysiwyg = "true";
defparam \rsc_block:sig_count[2] .power_up = "low";

arriaii_lcell_comb \sig_test_dq_expired~0 (
	.dataa(!\sig_dimm_driving_dq~q ),
	.datab(!\rsc_block:sig_count[0]~q ),
	.datac(!\rsc_block:sig_test_dq_expired~q ),
	.datad(!\rsc_block:sig_curr_byte_ln_dis~q ),
	.datae(!\sig_mtp_match~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_test_dq_expired~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_test_dq_expired~0 .extended_lut = "off";
defparam \sig_test_dq_expired~0 .lut_mask = 64'h0020000000200000;
defparam \sig_test_dq_expired~0 .shared_arith = "off";

arriaii_lcell_comb \sig_test_dq_expired~1 (
	.dataa(!\rsc_block:sig_count[1]~q ),
	.datab(!\rsc_block:sig_count[2]~q ),
	.datac(!\rsc_block:sig_count[3]~q ),
	.datad(!\Equal14~0_combout ),
	.datae(!\sig_test_dq_expired~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_test_dq_expired~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_test_dq_expired~1 .extended_lut = "off";
defparam \sig_test_dq_expired~1 .lut_mask = 64'h0000008000000080;
defparam \sig_test_dq_expired~1 .shared_arith = "off";

dffeas \rsc_block:sig_test_dq_expired (
	.clk(clk),
	.d(\sig_test_dq_expired~1_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.sload(!\rsc_block:sig_rsc_last_state.s_rsc_test_dq~q ),
	.ena(vcc),
	.q(\rsc_block:sig_test_dq_expired~q ),
	.prn(vcc));
defparam \rsc_block:sig_test_dq_expired .is_wysiwyg = "true";
defparam \rsc_block:sig_test_dq_expired .power_up = "low";

arriaii_lcell_comb \Selector53~0 (
	.dataa(!\sig_dimm_driving_dq~q ),
	.datab(!\rsc_block:sig_rsc_last_state.s_rsc_test_dq~q ),
	.datac(!\rsc_block:sig_test_dq_expired~q ),
	.datad(!\rsc_block:sig_curr_byte_ln_dis~q ),
	.datae(!\sig_mtp_match~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector53~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector53~0 .extended_lut = "off";
defparam \Selector53~0 .lut_mask = 64'h2202222222022222;
defparam \Selector53~0 .shared_arith = "off";

arriaii_lcell_comb \Selector52~0 (
	.dataa(!\sig_dimm_driving_dq~q ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_wait_for_idle_dimm~q ),
	.datac(!\rsc_block:sig_rsc_state.s_rsc_test_phase~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector52~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector52~0 .extended_lut = "off";
defparam \Selector52~0 .lut_mask = 64'h2F2F2F2F2F2F2F2F;
defparam \Selector52~0 .shared_arith = "off";

dffeas \rsc_block:sig_rsc_state.s_rsc_wait_for_idle_dimm (
	.clk(clk),
	.d(\Selector52~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rsc_state.s_rsc_wait_for_idle_dimm~q ),
	.prn(vcc));
defparam \rsc_block:sig_rsc_state.s_rsc_wait_for_idle_dimm .is_wysiwyg = "true";
defparam \rsc_block:sig_rsc_state.s_rsc_wait_for_idle_dimm .power_up = "low";

arriaii_lcell_comb \Selector53~1 (
	.dataa(!\sig_dimm_driving_dq~q ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datac(!\rsc_block:sig_chkd_all_dq_pins~q ),
	.datad(!\Selector53~0_combout ),
	.datae(!\rsc_block:sig_rsc_state.s_rsc_wait_for_idle_dimm~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector53~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector53~1 .extended_lut = "off";
defparam \Selector53~1 .lut_mask = 64'h0030557500305575;
defparam \Selector53~1 .shared_arith = "off";

arriaii_lcell_comb \Selector53~2 (
	.dataa(!\sig_dimm_driving_dq~q ),
	.datab(!\Equal14~1_combout ),
	.datac(!\rsc_block:sig_rsc_state.s_rsc_flush_datapath~q ),
	.datad(!\rsc_block:sig_rsc_last_state.s_rsc_flush_datapath~q ),
	.datae(!\Selector53~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector53~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector53~2 .extended_lut = "off";
defparam \Selector53~2 .lut_mask = 64'h0F0DFFFF0F0DFFFF;
defparam \Selector53~2 .shared_arith = "off";

dffeas \rsc_block:sig_rsc_state.s_rsc_flush_datapath (
	.clk(clk),
	.d(\Selector53~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rsc_state.s_rsc_flush_datapath~q ),
	.prn(vcc));
defparam \rsc_block:sig_rsc_state.s_rsc_flush_datapath .is_wysiwyg = "true";
defparam \rsc_block:sig_rsc_state.s_rsc_flush_datapath .power_up = "low";

dffeas \rsc_block:sig_rsc_last_state.s_rsc_flush_datapath (
	.clk(clk),
	.d(\rsc_block:sig_rsc_state.s_rsc_flush_datapath~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rsc_last_state.s_rsc_flush_datapath~q ),
	.prn(vcc));
defparam \rsc_block:sig_rsc_last_state.s_rsc_flush_datapath .is_wysiwyg = "true";
defparam \rsc_block:sig_rsc_last_state.s_rsc_flush_datapath .power_up = "low";

arriaii_lcell_comb \Selector47~0 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_flush_datapath~q ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_idle~q ),
	.datac(!\rsc_block:sig_rsc_last_state.s_rsc_flush_datapath~q ),
	.datad(!\Add6~5_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector47~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector47~0 .extended_lut = "off";
defparam \Selector47~0 .lut_mask = 64'h5073507350735073;
defparam \Selector47~0 .shared_arith = "off";

arriaii_lcell_comb \Selector47~1 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datab(!\rsc_block:sig_rsc_last_state.s_rsc_test_dq~q ),
	.datac(!\rsc_block:sig_count[6]~0_combout ),
	.datad(!\sig_cdvw_state.largest_window_centre[1]~q ),
	.datae(!\Selector47~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector47~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector47~1 .extended_lut = "off";
defparam \Selector47~1 .lut_mask = 64'h000FB0BF000FB0BF;
defparam \Selector47~1 .shared_arith = "off";

dffeas \rsc_block:sig_count[1] (
	.clk(clk),
	.d(\Selector47~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rsc_block:sig_count[2]~2_combout ),
	.q(\rsc_block:sig_count[1]~q ),
	.prn(vcc));
defparam \rsc_block:sig_count[1] .is_wysiwyg = "true";
defparam \rsc_block:sig_count[1] .power_up = "low";

arriaii_lcell_comb \Equal14~1 (
	.dataa(!\rsc_block:sig_count[0]~q ),
	.datab(!\rsc_block:sig_count[1]~q ),
	.datac(!\rsc_block:sig_count[2]~q ),
	.datad(!\rsc_block:sig_count[3]~q ),
	.datae(!\Equal14~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal14~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal14~1 .extended_lut = "off";
defparam \Equal14~1 .lut_mask = 64'h0000800000008000;
defparam \Equal14~1 .shared_arith = "off";

arriaii_lcell_comb \Selector54~0 (
	.dataa(!\sig_dimm_driving_dq~q ),
	.datab(!\Equal14~1_combout ),
	.datac(!\rsc_block:sig_rsc_state.s_rsc_flush_datapath~q ),
	.datad(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datae(!\Selector53~0_combout ),
	.dataf(!\rsc_block:sig_rsc_last_state.s_rsc_flush_datapath~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector54~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector54~0 .extended_lut = "off";
defparam \Selector54~0 .lut_mask = 64'h00FF000002FF0202;
defparam \Selector54~0 .shared_arith = "off";

dffeas \rsc_block:sig_rsc_state.s_rsc_test_dq (
	.clk(clk),
	.d(\Selector54~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.prn(vcc));
defparam \rsc_block:sig_rsc_state.s_rsc_test_dq .is_wysiwyg = "true";
defparam \rsc_block:sig_rsc_state.s_rsc_test_dq .power_up = "low";

dffeas \sig_dq_pin_ctr[0] (
	.clk(clk),
	.d(\Add7~1_sumout ),
	.asdata(\single_bit_cal~_wirecell_combout ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_dq_pin_ctr[0]~0_combout ),
	.sload(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.ena(\sig_dq_pin_ctr[0]~1_combout ),
	.q(\sig_dq_pin_ctr[0]~q ),
	.prn(vcc));
defparam \sig_dq_pin_ctr[0] .is_wysiwyg = "true";
defparam \sig_dq_pin_ctr[0] .power_up = "low";

dffeas \sig_dq_pin_ctr[1] (
	.clk(clk),
	.d(\Add7~5_sumout ),
	.asdata(\single_bit_cal~_wirecell_combout ),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_dq_pin_ctr[0]~0_combout ),
	.sload(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.ena(\sig_dq_pin_ctr[0]~1_combout ),
	.q(\sig_dq_pin_ctr[1]~q ),
	.prn(vcc));
defparam \sig_dq_pin_ctr[1] .is_wysiwyg = "true";
defparam \sig_dq_pin_ctr[1] .power_up = "low";

arriaii_lcell_comb \Equal11~0 (
	.dataa(!\sig_dq_pin_ctr[0]~q ),
	.datab(!\sig_dq_pin_ctr[1]~q ),
	.datac(!\sig_dq_pin_ctr[2]~q ),
	.datad(!\sig_dq_pin_ctr[4]~q ),
	.datae(!\sig_dq_pin_ctr[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal11~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal11~0 .extended_lut = "off";
defparam \Equal11~0 .lut_mask = 64'h8000000080000000;
defparam \Equal11~0 .shared_arith = "off";

dffeas \rsc_block:sig_chkd_all_dq_pins (
	.clk(clk),
	.d(\Equal11~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_chkd_all_dq_pins~q ),
	.prn(vcc));
defparam \rsc_block:sig_chkd_all_dq_pins .is_wysiwyg = "true";
defparam \rsc_block:sig_chkd_all_dq_pins .power_up = "low";

arriaii_lcell_comb \sig_rsc_cdvw_shift_in~0 (
	.dataa(!\sig_dimm_driving_dq~q ),
	.datab(!\rsc_block:sig_chkd_all_dq_pins~q ),
	.datac(!\rsc_block:sig_test_dq_expired~q ),
	.datad(!\rsc_block:sig_curr_byte_ln_dis~q ),
	.datae(!\sig_mtp_match~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_rsc_cdvw_shift_in~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_rsc_cdvw_shift_in~0 .extended_lut = "off";
defparam \sig_rsc_cdvw_shift_in~0 .lut_mask = 64'h2202222222022222;
defparam \sig_rsc_cdvw_shift_in~0 .shared_arith = "off";

dffeas sig_rsc_cdvw_shift_in(
	.clk(clk),
	.d(\sig_rsc_cdvw_shift_in~0_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.sload(!\rsc_block:sig_rsc_last_state.s_rsc_test_dq~q ),
	.ena(vcc),
	.q(\sig_rsc_cdvw_shift_in~q ),
	.prn(vcc));
defparam sig_rsc_cdvw_shift_in.is_wysiwyg = "true";
defparam sig_rsc_cdvw_shift_in.power_up = "low";

arriaii_lcell_comb \v_cdvw_state~20 (
	.dataa(!\sig_dgrb_state.s_seek_cdvw~q ),
	.datab(!\sig_dgrb_state.s_test_phases~q ),
	.datac(!\sig_dgrb_state.s_read_mtp~q ),
	.datad(!\sig_rsc_cdvw_shift_in~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~20 .extended_lut = "off";
defparam \v_cdvw_state~20 .lut_mask = 64'h007F007F007F007F;
defparam \v_cdvw_state~20 .shared_arith = "off";

arriaii_lcell_comb \sig_cdvw_state.working_window[23]~0 (
	.dataa(!\sig_dgrb_state.s_track~q ),
	.datab(!\sig_cdvw_state.status.calculating~q ),
	.datac(!\sig_trk_cdvw_shift_in~q ),
	.datad(!\v_cdvw_state~20_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_cdvw_state.working_window[23]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_cdvw_state.working_window[23]~0 .extended_lut = "off";
defparam \sig_cdvw_state.working_window[23]~0 .lut_mask = 64'hC800C800C800C800;
defparam \sig_cdvw_state.working_window[23]~0 .shared_arith = "off";

arriaii_lcell_comb \Selector35~0 (
	.dataa(!\sig_dgrb_state.s_track~q ),
	.datab(!\sig_trk_cdvw_shift_in~q ),
	.datac(!\v_cdvw_state~20_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector35~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector35~0 .extended_lut = "off";
defparam \Selector35~0 .lut_mask = 64'hE0E0E0E0E0E0E0E0;
defparam \Selector35~0 .shared_arith = "off";

arriaii_lcell_comb \Selector68~0 (
	.dataa(!\sig_dimm_driving_dq~q ),
	.datab(!\rsc_block:sig_test_dq_expired~q ),
	.datac(!\rsc_block:sig_curr_byte_ln_dis~q ),
	.datad(!\sig_mtp_match~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector68~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector68~0 .extended_lut = "off";
defparam \Selector68~0 .lut_mask = 64'h0200020002000200;
defparam \Selector68~0 .shared_arith = "off";

arriaii_lcell_comb \Selector68~1 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datab(!\rsc_block:sig_rsc_last_state.s_rsc_test_dq~q ),
	.datac(!\rsc_block:sig_rsc_state.s_rsc_test_phase~q ),
	.datad(!\rsc_block:rsc_proc:v_phase_works~q ),
	.datae(!\Selector68~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector68~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector68~1 .extended_lut = "off";
defparam \Selector68~1 .lut_mask = 64'h0AFF0AEE0AFF0AEE;
defparam \Selector68~1 .shared_arith = "off";

dffeas \rsc_block:rsc_proc:v_phase_works (
	.clk(clk),
	.d(\Selector68~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:rsc_proc:v_phase_works~q ),
	.prn(vcc));
defparam \rsc_block:rsc_proc:v_phase_works .is_wysiwyg = "true";
defparam \rsc_block:rsc_proc:v_phase_works .power_up = "low";

arriaii_lcell_comb \sig_rsc_cdvw_phase~0 (
	.dataa(!\sig_dimm_driving_dq~q ),
	.datab(!\rsc_block:sig_chkd_all_dq_pins~q ),
	.datac(!\rsc_block:sig_curr_byte_ln_dis~q ),
	.datad(!\sig_mtp_match~q ),
	.datae(!\rsc_block:rsc_proc:v_phase_works~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_rsc_cdvw_phase~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_rsc_cdvw_phase~0 .extended_lut = "off";
defparam \sig_rsc_cdvw_phase~0 .lut_mask = 64'h0000202200002022;
defparam \sig_rsc_cdvw_phase~0 .shared_arith = "off";

dffeas sig_rsc_cdvw_phase(
	.clk(clk),
	.d(\sig_rsc_cdvw_phase~0_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.sload(!\rsc_block:sig_rsc_last_state.s_rsc_test_dq~q ),
	.ena(vcc),
	.q(\sig_rsc_cdvw_phase~q ),
	.prn(vcc));
defparam sig_rsc_cdvw_phase.is_wysiwyg = "true";
defparam sig_rsc_cdvw_phase.power_up = "low";

arriaii_lcell_comb \working_window~0 (
	.dataa(!\sig_dgrb_state.s_seek_cdvw~q ),
	.datab(!\sig_dgrb_state.s_test_phases~q ),
	.datac(!\sig_dgrb_state.s_read_mtp~q ),
	.datad(!\sig_rsc_cdvw_phase~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\working_window~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \working_window~0 .extended_lut = "off";
defparam \working_window~0 .lut_mask = 64'h007F007F007F007F;
defparam \working_window~0 .shared_arith = "off";

dffeas \trk_block:mmc_seq_value_r (
	.clk(clk),
	.d(mmc_seq_value),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rst_n),
	.q(\trk_block:mmc_seq_value_r~q ),
	.prn(vcc));
defparam \trk_block:mmc_seq_value_r .is_wysiwyg = "true";
defparam \trk_block:mmc_seq_value_r .power_up = "low";

arriaii_lcell_comb \sig_trk_cdvw_phase~0 (
	.dataa(!\trk_block:mmc_seq_req_sync:v_mmc_seq_done_3r~q ),
	.datab(!\trk_block:sig_mmc_seq_done_1t~q ),
	.datac(!\trk_block:mmc_seq_value_r~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_trk_cdvw_phase~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_trk_cdvw_phase~0 .extended_lut = "off";
defparam \sig_trk_cdvw_phase~0 .lut_mask = 64'h0202020202020202;
defparam \sig_trk_cdvw_phase~0 .shared_arith = "off";

dffeas sig_trk_cdvw_phase(
	.clk(clk),
	.d(\sig_trk_cdvw_phase~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_trk_cdvw_phase~q ),
	.prn(vcc));
defparam sig_trk_cdvw_phase.is_wysiwyg = "true";
defparam sig_trk_cdvw_phase.power_up = "low";

arriaii_lcell_comb \v_cdvw_state~56 (
	.dataa(!\sig_dgrb_state.s_track~q ),
	.datab(!\sig_cdvw_state.status.calculating~q ),
	.datac(!\sig_cdvw_state.working_window[0]~q ),
	.datad(!\working_window~0_combout ),
	.datae(!\sig_trk_cdvw_phase~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~56_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~56 .extended_lut = "off";
defparam \v_cdvw_state~56 .lut_mask = 64'h00C040C000C040C0;
defparam \v_cdvw_state~56 .shared_arith = "off";

dffeas \ctrl_dgrb_r.command.cmd_rrp_seek (
	.clk(clk),
	.d(\ctrl_dgrb.command.cmd_rrp_seek ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_dgrb_r.command.cmd_rrp_seek~q ),
	.prn(vcc));
defparam \ctrl_dgrb_r.command.cmd_rrp_seek .is_wysiwyg = "true";
defparam \ctrl_dgrb_r.command.cmd_rrp_seek .power_up = "low";

arriaii_lcell_comb \sig_dgrb_state~48 (
	.dataa(!\sig_dgrb_state.s_seek_cdvw~q ),
	.datab(!\sig_dgrb_state.s_wait_admin~q ),
	.datac(!\sig_dgrb_state~45_combout ),
	.datad(!\ctrl_dgrb_r.command.cmd_rrp_seek~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~48 .extended_lut = "off";
defparam \sig_dgrb_state~48 .lut_mask = 64'h0407040704070407;
defparam \sig_dgrb_state~48 .shared_arith = "off";

dffeas \sig_dgrb_state.s_seek_cdvw (
	.clk(clk),
	.d(\sig_dgrb_state~48_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgrb_state.s_seek_cdvw~q ),
	.prn(vcc));
defparam \sig_dgrb_state.s_seek_cdvw .is_wysiwyg = "true";
defparam \sig_dgrb_state.s_seek_cdvw .power_up = "low";

arriaii_lcell_comb \sig_cdvw_state.working_window[32]~2 (
	.dataa(!\sig_dgrb_state.s_track~q ),
	.datab(!\sig_cdvw_state.status.calculating~q ),
	.datac(!\sig_dgrb_state.s_seek_cdvw~q ),
	.datad(!\sig_dgrb_state.s_test_phases~q ),
	.datae(!\sig_dgrb_state.s_read_mtp~q ),
	.dataf(!\sig_rsc_cdvw_shift_in~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_cdvw_state.working_window[32]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_cdvw_state.working_window[32]~2 .extended_lut = "off";
defparam \sig_cdvw_state.working_window[32]~2 .lut_mask = 64'hCCCCCCCCC4444444;
defparam \sig_cdvw_state.working_window[32]~2 .shared_arith = "off";

arriaii_lcell_comb \v_cdvw_state~90 (
	.dataa(!\sig_dgrb_state.s_track~q ),
	.datab(!\sig_cdvw_state.status.calculating~q ),
	.datac(!\sig_cdvw_state.working_window[0]~q ),
	.datad(!\v_cdvw_state~20_combout ),
	.datae(!\v_cdvw_state~56_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~90_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~90 .extended_lut = "off";
defparam \v_cdvw_state~90 .lut_mask = 64'h313131BB313131BB;
defparam \v_cdvw_state~90 .shared_arith = "off";

arriaii_lcell_comb \v_cdvw_state~91 (
	.dataa(!\cdvw_proc~1_combout ),
	.datab(!\cdvw_proc~2_combout ),
	.datac(!\sig_cdvw_state.working_window[32]~2_combout ),
	.datad(!\sig_cdvw_state.working_window[63]~q ),
	.datae(!\v_cdvw_state~90_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~91_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~91 .extended_lut = "off";
defparam \v_cdvw_state~91 .lut_mask = 64'h80AA002280AA0022;
defparam \v_cdvw_state~91 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[63] (
	.clk(clk),
	.d(\v_cdvw_state~91_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_cdvw_state.working_window[63]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[63] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[63] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~89 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[63]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~89_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~89 .extended_lut = "off";
defparam \v_cdvw_state~89 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~89 .shared_arith = "off";

arriaii_lcell_comb \sig_cdvw_state.working_window[32]~3 (
	.dataa(!\cdvw_proc~1_combout ),
	.datab(!\sig_cdvw_state.working_window[32]~2_combout ),
	.datac(!\cdvw_block:sig_cdvw_calc_1t~q ),
	.datad(!\Selector33~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_cdvw_state.working_window[32]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_cdvw_state.working_window[32]~3 .extended_lut = "off";
defparam \sig_cdvw_state.working_window[32]~3 .lut_mask = 64'hDD5DDD5DDD5DDD5D;
defparam \sig_cdvw_state.working_window[32]~3 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[62] (
	.clk(clk),
	.d(\v_cdvw_state~89_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[32]~3_combout ),
	.q(\sig_cdvw_state.working_window[62]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[62] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[62] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~88 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[62]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~88_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~88 .extended_lut = "off";
defparam \v_cdvw_state~88 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~88 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[61] (
	.clk(clk),
	.d(\v_cdvw_state~88_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[32]~3_combout ),
	.q(\sig_cdvw_state.working_window[61]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[61] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[61] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~87 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[61]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~87_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~87 .extended_lut = "off";
defparam \v_cdvw_state~87 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~87 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[60] (
	.clk(clk),
	.d(\v_cdvw_state~87_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[32]~3_combout ),
	.q(\sig_cdvw_state.working_window[60]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[60] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[60] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~86 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[60]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~86_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~86 .extended_lut = "off";
defparam \v_cdvw_state~86 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~86 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[59] (
	.clk(clk),
	.d(\v_cdvw_state~86_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[32]~3_combout ),
	.q(\sig_cdvw_state.working_window[59]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[59] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[59] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~85 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[59]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~85_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~85 .extended_lut = "off";
defparam \v_cdvw_state~85 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~85 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[58] (
	.clk(clk),
	.d(\v_cdvw_state~85_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[32]~3_combout ),
	.q(\sig_cdvw_state.working_window[58]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[58] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[58] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~84 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[58]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~84_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~84 .extended_lut = "off";
defparam \v_cdvw_state~84 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~84 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[57] (
	.clk(clk),
	.d(\v_cdvw_state~84_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[32]~3_combout ),
	.q(\sig_cdvw_state.working_window[57]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[57] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[57] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~83 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[57]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~83_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~83 .extended_lut = "off";
defparam \v_cdvw_state~83 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~83 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[56] (
	.clk(clk),
	.d(\v_cdvw_state~83_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[32]~3_combout ),
	.q(\sig_cdvw_state.working_window[56]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[56] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[56] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~82 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[56]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~82_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~82 .extended_lut = "off";
defparam \v_cdvw_state~82 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~82 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[55] (
	.clk(clk),
	.d(\v_cdvw_state~82_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[32]~3_combout ),
	.q(\sig_cdvw_state.working_window[55]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[55] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[55] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~81 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[55]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~81_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~81 .extended_lut = "off";
defparam \v_cdvw_state~81 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~81 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[54] (
	.clk(clk),
	.d(\v_cdvw_state~81_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[32]~3_combout ),
	.q(\sig_cdvw_state.working_window[54]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[54] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[54] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~80 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[54]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~80_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~80 .extended_lut = "off";
defparam \v_cdvw_state~80 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~80 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[53] (
	.clk(clk),
	.d(\v_cdvw_state~80_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[32]~3_combout ),
	.q(\sig_cdvw_state.working_window[53]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[53] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[53] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~79 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[53]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~79_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~79 .extended_lut = "off";
defparam \v_cdvw_state~79 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~79 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[52] (
	.clk(clk),
	.d(\v_cdvw_state~79_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[32]~3_combout ),
	.q(\sig_cdvw_state.working_window[52]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[52] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[52] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~78 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[52]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~78_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~78 .extended_lut = "off";
defparam \v_cdvw_state~78 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~78 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[51] (
	.clk(clk),
	.d(\v_cdvw_state~78_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[32]~3_combout ),
	.q(\sig_cdvw_state.working_window[51]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[51] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[51] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~77 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[51]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~77_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~77 .extended_lut = "off";
defparam \v_cdvw_state~77 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~77 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[50] (
	.clk(clk),
	.d(\v_cdvw_state~77_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[32]~3_combout ),
	.q(\sig_cdvw_state.working_window[50]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[50] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[50] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~76 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[50]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~76_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~76 .extended_lut = "off";
defparam \v_cdvw_state~76 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~76 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[49] (
	.clk(clk),
	.d(\v_cdvw_state~76_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[32]~3_combout ),
	.q(\sig_cdvw_state.working_window[49]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[49] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[49] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~75 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[49]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~75_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~75 .extended_lut = "off";
defparam \v_cdvw_state~75 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~75 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[48] (
	.clk(clk),
	.d(\v_cdvw_state~75_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[32]~3_combout ),
	.q(\sig_cdvw_state.working_window[48]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[48] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[48] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~74 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[48]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~74_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~74 .extended_lut = "off";
defparam \v_cdvw_state~74 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~74 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[47] (
	.clk(clk),
	.d(\v_cdvw_state~74_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[32]~3_combout ),
	.q(\sig_cdvw_state.working_window[47]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[47] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[47] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~73 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[47]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~73_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~73 .extended_lut = "off";
defparam \v_cdvw_state~73 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~73 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[46] (
	.clk(clk),
	.d(\v_cdvw_state~73_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[32]~3_combout ),
	.q(\sig_cdvw_state.working_window[46]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[46] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[46] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~72 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[46]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~72_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~72 .extended_lut = "off";
defparam \v_cdvw_state~72 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~72 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[45] (
	.clk(clk),
	.d(\v_cdvw_state~72_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[32]~3_combout ),
	.q(\sig_cdvw_state.working_window[45]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[45] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[45] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~71 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[45]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~71_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~71 .extended_lut = "off";
defparam \v_cdvw_state~71 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~71 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[44] (
	.clk(clk),
	.d(\v_cdvw_state~71_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[32]~3_combout ),
	.q(\sig_cdvw_state.working_window[44]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[44] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[44] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~70 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[44]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~70_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~70 .extended_lut = "off";
defparam \v_cdvw_state~70 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~70 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[43] (
	.clk(clk),
	.d(\v_cdvw_state~70_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[32]~3_combout ),
	.q(\sig_cdvw_state.working_window[43]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[43] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[43] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~69 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[43]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~69_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~69 .extended_lut = "off";
defparam \v_cdvw_state~69 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~69 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[42] (
	.clk(clk),
	.d(\v_cdvw_state~69_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[32]~3_combout ),
	.q(\sig_cdvw_state.working_window[42]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[42] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[42] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~68 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[42]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~68_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~68 .extended_lut = "off";
defparam \v_cdvw_state~68 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~68 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[41] (
	.clk(clk),
	.d(\v_cdvw_state~68_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[32]~3_combout ),
	.q(\sig_cdvw_state.working_window[41]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[41] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[41] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~67 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[41]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~67_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~67 .extended_lut = "off";
defparam \v_cdvw_state~67 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~67 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[40] (
	.clk(clk),
	.d(\v_cdvw_state~67_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[32]~3_combout ),
	.q(\sig_cdvw_state.working_window[40]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[40] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[40] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~66 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[40]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~66_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~66 .extended_lut = "off";
defparam \v_cdvw_state~66 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~66 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[39] (
	.clk(clk),
	.d(\v_cdvw_state~66_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[32]~3_combout ),
	.q(\sig_cdvw_state.working_window[39]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[39] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[39] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~65 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[39]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~65_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~65 .extended_lut = "off";
defparam \v_cdvw_state~65 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~65 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[38] (
	.clk(clk),
	.d(\v_cdvw_state~65_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[32]~3_combout ),
	.q(\sig_cdvw_state.working_window[38]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[38] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[38] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~64 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[38]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~64_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~64 .extended_lut = "off";
defparam \v_cdvw_state~64 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~64 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[37] (
	.clk(clk),
	.d(\v_cdvw_state~64_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[32]~3_combout ),
	.q(\sig_cdvw_state.working_window[37]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[37] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[37] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~63 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[37]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~63_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~63 .extended_lut = "off";
defparam \v_cdvw_state~63 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~63 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[36] (
	.clk(clk),
	.d(\v_cdvw_state~63_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[32]~3_combout ),
	.q(\sig_cdvw_state.working_window[36]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[36] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[36] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~62 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[36]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~62_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~62 .extended_lut = "off";
defparam \v_cdvw_state~62 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~62 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[35] (
	.clk(clk),
	.d(\v_cdvw_state~62_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[32]~3_combout ),
	.q(\sig_cdvw_state.working_window[35]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[35] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[35] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~61 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[35]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~61_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~61 .extended_lut = "off";
defparam \v_cdvw_state~61 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~61 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[34] (
	.clk(clk),
	.d(\v_cdvw_state~61_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[32]~3_combout ),
	.q(\sig_cdvw_state.working_window[34]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[34] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[34] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~60 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[34]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~60_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~60 .extended_lut = "off";
defparam \v_cdvw_state~60 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~60 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[33] (
	.clk(clk),
	.d(\v_cdvw_state~60_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[32]~3_combout ),
	.q(\sig_cdvw_state.working_window[33]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[33] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[33] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~59 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[33]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~59_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~59 .extended_lut = "off";
defparam \v_cdvw_state~59 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~59 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[32] (
	.clk(clk),
	.d(\v_cdvw_state~59_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[32]~3_combout ),
	.q(\sig_cdvw_state.working_window[32]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[32] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[32] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~57 (
	.dataa(!\sig_dgrb_state.s_track~q ),
	.datab(!\sig_cdvw_state.status.calculating~q ),
	.datac(!\sig_cdvw_state.working_window[0]~q ),
	.datad(!\Selector35~0_combout ),
	.datae(!\v_cdvw_state~56_combout ),
	.dataf(!\sig_cdvw_state.working_window[32]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~57_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~57 .extended_lut = "off";
defparam \v_cdvw_state~57 .lut_mask = 64'hBA32FF3210105510;
defparam \v_cdvw_state~57 .shared_arith = "off";

arriaii_lcell_comb \v_cdvw_state~58 (
	.dataa(!\cdvw_proc~1_combout ),
	.datab(!\cdvw_proc~2_combout ),
	.datac(!\sig_cdvw_state.working_window[23]~0_combout ),
	.datad(!\sig_cdvw_state.working_window[31]~q ),
	.datae(!\v_cdvw_state~57_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~58_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~58 .extended_lut = "off";
defparam \v_cdvw_state~58 .lut_mask = 64'h80AA002280AA0022;
defparam \v_cdvw_state~58 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[31] (
	.clk(clk),
	.d(\v_cdvw_state~58_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_cdvw_state.working_window[31]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[31] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[31] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~55 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[31]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~55_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~55 .extended_lut = "off";
defparam \v_cdvw_state~55 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~55 .shared_arith = "off";

arriaii_lcell_comb \sig_cdvw_state.working_window[23]~4 (
	.dataa(!\sig_dgrb_state.s_track~q ),
	.datab(!\sig_trk_cdvw_shift_in~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_cdvw_state.working_window[23]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_cdvw_state.working_window[23]~4 .extended_lut = "off";
defparam \sig_cdvw_state.working_window[23]~4 .lut_mask = 64'h1111111111111111;
defparam \sig_cdvw_state.working_window[23]~4 .shared_arith = "off";

arriaii_lcell_comb \sig_cdvw_state.working_window[23]~1 (
	.dataa(!\cdvw_proc~1_combout ),
	.datab(!\cdvw_block:sig_cdvw_calc_1t~q ),
	.datac(!\Selector33~0_combout ),
	.datad(!\sig_cdvw_state.status.calculating~q ),
	.datae(!\v_cdvw_state~20_combout ),
	.dataf(!\sig_cdvw_state.working_window[23]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_cdvw_state.working_window[23]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_cdvw_state.working_window[23]~1 .extended_lut = "off";
defparam \sig_cdvw_state.working_window[23]~1 .lut_mask = 64'h55F7F7F7F7F7F7F7;
defparam \sig_cdvw_state.working_window[23]~1 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[30] (
	.clk(clk),
	.d(\v_cdvw_state~55_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[23]~1_combout ),
	.q(\sig_cdvw_state.working_window[30]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[30] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[30] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~54 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[30]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~54_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~54 .extended_lut = "off";
defparam \v_cdvw_state~54 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~54 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[29] (
	.clk(clk),
	.d(\v_cdvw_state~54_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[23]~1_combout ),
	.q(\sig_cdvw_state.working_window[29]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[29] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[29] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~53 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[29]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~53_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~53 .extended_lut = "off";
defparam \v_cdvw_state~53 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~53 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[28] (
	.clk(clk),
	.d(\v_cdvw_state~53_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[23]~1_combout ),
	.q(\sig_cdvw_state.working_window[28]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[28] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[28] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~52 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[28]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~52 .extended_lut = "off";
defparam \v_cdvw_state~52 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~52 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[27] (
	.clk(clk),
	.d(\v_cdvw_state~52_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[23]~1_combout ),
	.q(\sig_cdvw_state.working_window[27]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[27] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[27] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~51 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[27]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~51 .extended_lut = "off";
defparam \v_cdvw_state~51 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~51 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[26] (
	.clk(clk),
	.d(\v_cdvw_state~51_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[23]~1_combout ),
	.q(\sig_cdvw_state.working_window[26]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[26] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[26] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~50 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[26]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~50_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~50 .extended_lut = "off";
defparam \v_cdvw_state~50 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~50 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[25] (
	.clk(clk),
	.d(\v_cdvw_state~50_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[23]~1_combout ),
	.q(\sig_cdvw_state.working_window[25]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[25] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[25] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~49 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[25]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~49 .extended_lut = "off";
defparam \v_cdvw_state~49 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~49 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[24] (
	.clk(clk),
	.d(\v_cdvw_state~49_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[23]~1_combout ),
	.q(\sig_cdvw_state.working_window[24]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[24] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[24] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~48 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[24]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~48 .extended_lut = "off";
defparam \v_cdvw_state~48 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~48 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[23] (
	.clk(clk),
	.d(\v_cdvw_state~48_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[23]~1_combout ),
	.q(\sig_cdvw_state.working_window[23]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[23] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[23] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~47 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[23]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~47 .extended_lut = "off";
defparam \v_cdvw_state~47 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~47 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[22] (
	.clk(clk),
	.d(\v_cdvw_state~47_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[23]~1_combout ),
	.q(\sig_cdvw_state.working_window[22]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[22] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[22] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~46 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[22]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~46 .extended_lut = "off";
defparam \v_cdvw_state~46 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~46 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[21] (
	.clk(clk),
	.d(\v_cdvw_state~46_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[23]~1_combout ),
	.q(\sig_cdvw_state.working_window[21]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[21] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[21] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~45 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[21]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~45 .extended_lut = "off";
defparam \v_cdvw_state~45 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~45 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[20] (
	.clk(clk),
	.d(\v_cdvw_state~45_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[23]~1_combout ),
	.q(\sig_cdvw_state.working_window[20]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[20] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[20] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~44 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[20]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~44 .extended_lut = "off";
defparam \v_cdvw_state~44 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~44 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[19] (
	.clk(clk),
	.d(\v_cdvw_state~44_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[23]~1_combout ),
	.q(\sig_cdvw_state.working_window[19]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[19] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[19] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~43 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[19]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~43 .extended_lut = "off";
defparam \v_cdvw_state~43 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~43 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[18] (
	.clk(clk),
	.d(\v_cdvw_state~43_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[23]~1_combout ),
	.q(\sig_cdvw_state.working_window[18]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[18] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[18] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~42 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[18]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~42 .extended_lut = "off";
defparam \v_cdvw_state~42 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~42 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[17] (
	.clk(clk),
	.d(\v_cdvw_state~42_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[23]~1_combout ),
	.q(\sig_cdvw_state.working_window[17]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[17] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[17] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~41 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[17]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~41 .extended_lut = "off";
defparam \v_cdvw_state~41 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~41 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[16] (
	.clk(clk),
	.d(\v_cdvw_state~41_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[23]~1_combout ),
	.q(\sig_cdvw_state.working_window[16]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[16] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[16] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~40 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[16]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~40 .extended_lut = "off";
defparam \v_cdvw_state~40 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~40 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[15] (
	.clk(clk),
	.d(\v_cdvw_state~40_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[23]~1_combout ),
	.q(\sig_cdvw_state.working_window[15]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[15] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[15] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~39 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~39 .extended_lut = "off";
defparam \v_cdvw_state~39 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~39 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[14] (
	.clk(clk),
	.d(\v_cdvw_state~39_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[23]~1_combout ),
	.q(\sig_cdvw_state.working_window[14]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[14] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[14] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~38 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~38 .extended_lut = "off";
defparam \v_cdvw_state~38 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~38 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[13] (
	.clk(clk),
	.d(\v_cdvw_state~38_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[23]~1_combout ),
	.q(\sig_cdvw_state.working_window[13]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[13] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[13] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~37 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~37 .extended_lut = "off";
defparam \v_cdvw_state~37 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~37 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[12] (
	.clk(clk),
	.d(\v_cdvw_state~37_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[23]~1_combout ),
	.q(\sig_cdvw_state.working_window[12]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[12] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[12] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~36 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~36 .extended_lut = "off";
defparam \v_cdvw_state~36 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~36 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[11] (
	.clk(clk),
	.d(\v_cdvw_state~36_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[23]~1_combout ),
	.q(\sig_cdvw_state.working_window[11]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[11] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[11] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~35 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~35 .extended_lut = "off";
defparam \v_cdvw_state~35 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~35 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[10] (
	.clk(clk),
	.d(\v_cdvw_state~35_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[23]~1_combout ),
	.q(\sig_cdvw_state.working_window[10]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[10] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[10] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~34 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~34 .extended_lut = "off";
defparam \v_cdvw_state~34 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~34 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[9] (
	.clk(clk),
	.d(\v_cdvw_state~34_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[23]~1_combout ),
	.q(\sig_cdvw_state.working_window[9]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[9] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[9] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~33 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~33 .extended_lut = "off";
defparam \v_cdvw_state~33 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~33 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[8] (
	.clk(clk),
	.d(\v_cdvw_state~33_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[23]~1_combout ),
	.q(\sig_cdvw_state.working_window[8]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[8] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[8] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~32 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~32 .extended_lut = "off";
defparam \v_cdvw_state~32 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~32 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[7] (
	.clk(clk),
	.d(\v_cdvw_state~32_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[23]~1_combout ),
	.q(\sig_cdvw_state.working_window[7]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[7] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[7] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~28 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~28 .extended_lut = "off";
defparam \v_cdvw_state~28 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~28 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[6] (
	.clk(clk),
	.d(\v_cdvw_state~28_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[23]~1_combout ),
	.q(\sig_cdvw_state.working_window[6]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[6] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[6] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~27 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~27 .extended_lut = "off";
defparam \v_cdvw_state~27 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~27 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[5] (
	.clk(clk),
	.d(\v_cdvw_state~27_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[23]~1_combout ),
	.q(\sig_cdvw_state.working_window[5]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[5] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[5] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~26 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~26 .extended_lut = "off";
defparam \v_cdvw_state~26 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~26 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[4] (
	.clk(clk),
	.d(\v_cdvw_state~26_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[23]~1_combout ),
	.q(\sig_cdvw_state.working_window[4]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[4] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[4] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~25 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~25 .extended_lut = "off";
defparam \v_cdvw_state~25 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~25 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[3] (
	.clk(clk),
	.d(\v_cdvw_state~25_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[23]~1_combout ),
	.q(\sig_cdvw_state.working_window[3]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[3] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[3] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~24 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~24 .extended_lut = "off";
defparam \v_cdvw_state~24 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~24 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[2] (
	.clk(clk),
	.d(\v_cdvw_state~24_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[23]~1_combout ),
	.q(\sig_cdvw_state.working_window[2]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[2] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[2] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~23 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~23 .extended_lut = "off";
defparam \v_cdvw_state~23 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~23 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[1] (
	.clk(clk),
	.d(\v_cdvw_state~23_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[23]~1_combout ),
	.q(\sig_cdvw_state.working_window[1]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[1] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[1] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~19 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_last_state.s_track~q ),
	.datad(!\sig_cdvw_state.working_window[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~19 .extended_lut = "off";
defparam \v_cdvw_state~19 .lut_mask = 64'h008A008A008A008A;
defparam \v_cdvw_state~19 .shared_arith = "off";

dffeas \sig_cdvw_state.working_window[0] (
	.clk(clk),
	.d(\v_cdvw_state~19_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.working_window[23]~1_combout ),
	.q(\sig_cdvw_state.working_window[0]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.working_window[0] .is_wysiwyg = "true";
defparam \sig_cdvw_state.working_window[0] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~8 (
	.dataa(!\sig_cdvw_state.status.calculating~q ),
	.datab(!\sig_cdvw_state.valid_phase_seen~q ),
	.datac(!\v_cdvw_state~2_combout ),
	.datad(!\sig_cdvw_state.working_window[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~8 .extended_lut = "off";
defparam \v_cdvw_state~8 .lut_mask = 64'h7030703070307030;
defparam \v_cdvw_state~8 .shared_arith = "off";

dffeas \sig_cdvw_state.valid_phase_seen (
	.clk(clk),
	.d(\v_cdvw_state~8_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_cdvw_state.valid_phase_seen~q ),
	.prn(vcc));
defparam \sig_cdvw_state.valid_phase_seen .is_wysiwyg = "true";
defparam \sig_cdvw_state.valid_phase_seen .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~9 (
	.dataa(!\sig_cdvw_state.status.calculating~q ),
	.datab(!\sig_cdvw_state.first_cycle~q ),
	.datac(!\cdvw_proc~1_combout ),
	.datad(!\cdvw_block:sig_cdvw_calc_1t~q ),
	.datae(!\Selector33~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~9 .extended_lut = "off";
defparam \v_cdvw_state~9 .lut_mask = 64'h2020F0202020F020;
defparam \v_cdvw_state~9 .shared_arith = "off";

dffeas \sig_cdvw_state.first_cycle (
	.clk(clk),
	.d(\v_cdvw_state~9_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_cdvw_state.first_cycle~q ),
	.prn(vcc));
defparam \sig_cdvw_state.first_cycle .is_wysiwyg = "true";
defparam \sig_cdvw_state.first_cycle .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~10 (
	.dataa(!\sig_cdvw_state.current_bit[2]~q ),
	.datab(!\cdvw_proc~1_combout ),
	.datac(!\cdvw_block:sig_cdvw_calc_1t~q ),
	.datad(!\Selector33~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~10 .extended_lut = "off";
defparam \v_cdvw_state~10 .lut_mask = 64'h4404440444044404;
defparam \v_cdvw_state~10 .shared_arith = "off";

arriaii_lcell_comb \sig_cdvw_state.first_good_edge[0]~0 (
	.dataa(!\sig_cdvw_state.status.calculating~q ),
	.datab(!\sig_cdvw_state.found_a_good_edge~q ),
	.datac(!\find_centre_of_largest_data_valid_window~2_combout ),
	.datad(!\cdvw_proc~1_combout ),
	.datae(!\cdvw_block:sig_cdvw_calc_1t~q ),
	.dataf(!\Selector33~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_cdvw_state.first_good_edge[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_cdvw_state.first_good_edge[0]~0 .extended_lut = "off";
defparam \sig_cdvw_state.first_good_edge[0]~0 .lut_mask = 64'h04FF04FFFFFF04FF;
defparam \sig_cdvw_state.first_good_edge[0]~0 .shared_arith = "off";

dffeas \sig_cdvw_state.first_good_edge[2] (
	.clk(clk),
	.d(\v_cdvw_state~10_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.first_good_edge[0]~0_combout ),
	.q(\sig_cdvw_state.first_good_edge[2]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.first_good_edge[2] .is_wysiwyg = "true";
defparam \sig_cdvw_state.first_good_edge[2] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~11 (
	.dataa(!\sig_cdvw_state.current_bit[0]~q ),
	.datab(!\cdvw_proc~1_combout ),
	.datac(!\cdvw_block:sig_cdvw_calc_1t~q ),
	.datad(!\Selector33~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~11 .extended_lut = "off";
defparam \v_cdvw_state~11 .lut_mask = 64'h4404440444044404;
defparam \v_cdvw_state~11 .shared_arith = "off";

dffeas \sig_cdvw_state.first_good_edge[0] (
	.clk(clk),
	.d(\v_cdvw_state~11_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.first_good_edge[0]~0_combout ),
	.q(\sig_cdvw_state.first_good_edge[0]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.first_good_edge[0] .is_wysiwyg = "true";
defparam \sig_cdvw_state.first_good_edge[0] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~12 (
	.dataa(!\sig_cdvw_state.current_bit[1]~q ),
	.datab(!\cdvw_proc~1_combout ),
	.datac(!\cdvw_block:sig_cdvw_calc_1t~q ),
	.datad(!\Selector33~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~12 .extended_lut = "off";
defparam \v_cdvw_state~12 .lut_mask = 64'h4404440444044404;
defparam \v_cdvw_state~12 .shared_arith = "off";

dffeas \sig_cdvw_state.first_good_edge[1] (
	.clk(clk),
	.d(\v_cdvw_state~12_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.first_good_edge[0]~0_combout ),
	.q(\sig_cdvw_state.first_good_edge[1]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.first_good_edge[1] .is_wysiwyg = "true";
defparam \sig_cdvw_state.first_good_edge[1] .power_up = "low";

arriaii_lcell_comb \Equal9~0 (
	.dataa(!\sig_cdvw_state.current_bit[0]~q ),
	.datab(!\sig_cdvw_state.current_bit[1]~q ),
	.datac(!\sig_cdvw_state.first_good_edge[0]~q ),
	.datad(!\sig_cdvw_state.first_good_edge[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal9~0 .extended_lut = "off";
defparam \Equal9~0 .lut_mask = 64'h8421842184218421;
defparam \Equal9~0 .shared_arith = "off";

arriaii_lcell_comb \v_cdvw_state~13 (
	.dataa(!\sig_cdvw_state.current_bit[5]~q ),
	.datab(!\cdvw_proc~1_combout ),
	.datac(!\cdvw_block:sig_cdvw_calc_1t~q ),
	.datad(!\Selector33~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~13 .extended_lut = "off";
defparam \v_cdvw_state~13 .lut_mask = 64'h4404440444044404;
defparam \v_cdvw_state~13 .shared_arith = "off";

dffeas \sig_cdvw_state.first_good_edge[5] (
	.clk(clk),
	.d(\v_cdvw_state~13_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.first_good_edge[0]~0_combout ),
	.q(\sig_cdvw_state.first_good_edge[5]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.first_good_edge[5] .is_wysiwyg = "true";
defparam \sig_cdvw_state.first_good_edge[5] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~14 (
	.dataa(!\sig_cdvw_state.current_bit[3]~q ),
	.datab(!\cdvw_proc~1_combout ),
	.datac(!\cdvw_block:sig_cdvw_calc_1t~q ),
	.datad(!\Selector33~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~14 .extended_lut = "off";
defparam \v_cdvw_state~14 .lut_mask = 64'h4404440444044404;
defparam \v_cdvw_state~14 .shared_arith = "off";

dffeas \sig_cdvw_state.first_good_edge[3] (
	.clk(clk),
	.d(\v_cdvw_state~14_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.first_good_edge[0]~0_combout ),
	.q(\sig_cdvw_state.first_good_edge[3]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.first_good_edge[3] .is_wysiwyg = "true";
defparam \sig_cdvw_state.first_good_edge[3] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~15 (
	.dataa(!\sig_cdvw_state.current_bit[4]~q ),
	.datab(!\cdvw_proc~1_combout ),
	.datac(!\cdvw_block:sig_cdvw_calc_1t~q ),
	.datad(!\Selector33~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~15 .extended_lut = "off";
defparam \v_cdvw_state~15 .lut_mask = 64'h4404440444044404;
defparam \v_cdvw_state~15 .shared_arith = "off";

dffeas \sig_cdvw_state.first_good_edge[4] (
	.clk(clk),
	.d(\v_cdvw_state~15_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_cdvw_state.first_good_edge[0]~0_combout ),
	.q(\sig_cdvw_state.first_good_edge[4]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.first_good_edge[4] .is_wysiwyg = "true";
defparam \sig_cdvw_state.first_good_edge[4] .power_up = "low";

arriaii_lcell_comb \Equal9~1 (
	.dataa(!\sig_cdvw_state.current_bit[3]~q ),
	.datab(!\sig_cdvw_state.current_bit[4]~q ),
	.datac(!\sig_cdvw_state.first_good_edge[3]~q ),
	.datad(!\sig_cdvw_state.first_good_edge[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal9~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal9~1 .extended_lut = "off";
defparam \Equal9~1 .lut_mask = 64'h8421842184218421;
defparam \Equal9~1 .shared_arith = "off";

arriaii_lcell_comb \Equal9~2 (
	.dataa(!\sig_cdvw_state.current_bit[2]~q ),
	.datab(!\sig_cdvw_state.current_bit[5]~q ),
	.datac(!\sig_cdvw_state.first_good_edge[2]~q ),
	.datad(!\Equal9~0_combout ),
	.datae(!\sig_cdvw_state.first_good_edge[5]~q ),
	.dataf(!\Equal9~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal9~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal9~2 .extended_lut = "off";
defparam \Equal9~2 .lut_mask = 64'h0000000000840021;
defparam \Equal9~2 .shared_arith = "off";

arriaii_lcell_comb \v_cdvw_state~0 (
	.dataa(!\sig_cdvw_state.invalid_phase_seen~q ),
	.datab(!\sig_cdvw_state.valid_phase_seen~q ),
	.datac(!\find_centre_of_largest_data_valid_window~1_combout ),
	.datad(!\sig_cdvw_state.first_cycle~q ),
	.datae(!\Equal9~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~0 .extended_lut = "off";
defparam \v_cdvw_state~0 .lut_mask = 64'h0E00FE000E00FE00;
defparam \v_cdvw_state~0 .shared_arith = "off";

arriaii_lcell_comb \v_cdvw_state~4 (
	.dataa(!\sig_cdvw_state.status.calculating~q ),
	.datab(!\v_cdvw_state~0_combout ),
	.datac(!\cdvw_proc~1_combout ),
	.datad(!\cdvw_proc~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~4 .extended_lut = "off";
defparam \v_cdvw_state~4 .lut_mask = 64'h40F040F040F040F0;
defparam \v_cdvw_state~4 .shared_arith = "off";

dffeas \sig_cdvw_state.status.calculating (
	.clk(clk),
	.d(\v_cdvw_state~4_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_cdvw_state.status.calculating~q ),
	.prn(vcc));
defparam \sig_cdvw_state.status.calculating .is_wysiwyg = "true";
defparam \sig_cdvw_state.status.calculating .power_up = "low";

arriaii_lcell_comb \Selector128~1 (
	.dataa(!\sig_cdvw_state.status.valid_result~q ),
	.datab(!\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.datac(!\sig_cdvw_state.status.calculating~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector128~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector128~1 .extended_lut = "off";
defparam \Selector128~1 .lut_mask = 64'h2020202020202020;
defparam \Selector128~1 .shared_arith = "off";

arriaii_lcell_comb \sig_trk_state~27 (
	.dataa(!\sig_dgrb_state.s_track~q ),
	.datab(!sig_addr_cmd0cke0),
	.datac(!\Selector128~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_trk_state~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_trk_state~27 .extended_lut = "off";
defparam \sig_trk_state~27 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \sig_trk_state~27 .shared_arith = "off";

dffeas \trk_block:sig_trk_state.s_trk_idle (
	.clk(clk),
	.d(\sig_trk_state~27_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_trk_state.s_trk_idle~q ),
	.prn(vcc));
defparam \trk_block:sig_trk_state.s_trk_idle .is_wysiwyg = "true";
defparam \trk_block:sig_trk_state.s_trk_idle .power_up = "low";

arriaii_lcell_comb \Selector121~0 (
	.dataa(!\shift_in_mmc_seq_value~0_combout ),
	.datab(!\Equal17~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector121~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector121~0 .extended_lut = "off";
defparam \Selector121~0 .lut_mask = 64'h4444444444444444;
defparam \Selector121~0 .shared_arith = "off";

arriaii_lcell_comb \Add10~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_remaining_samples[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add10~1_sumout ),
	.cout(\Add10~2 ),
	.shareout());
defparam \Add10~1 .extended_lut = "off";
defparam \Add10~1 .lut_mask = 64'h00000000000000FF;
defparam \Add10~1 .shared_arith = "off";

arriaii_lcell_comb \Selector126~0 (
	.dataa(!\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.datab(!\trk_block:sig_remaining_samples[0]~q ),
	.datac(!\trk_block:sig_trk_state.s_trk_idle~q ),
	.datad(!\Add10~1_sumout ),
	.datae(!\Selector121~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector126~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector126~0 .extended_lut = "off";
defparam \Selector126~0 .lut_mask = 64'h3131207531312075;
defparam \Selector126~0 .shared_arith = "off";

dffeas \trk_block:sig_remaining_samples[0] (
	.clk(clk),
	.d(\Selector126~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_dgrb_state.s_track~q ),
	.q(\trk_block:sig_remaining_samples[0]~q ),
	.prn(vcc));
defparam \trk_block:sig_remaining_samples[0] .is_wysiwyg = "true";
defparam \trk_block:sig_remaining_samples[0] .power_up = "low";

arriaii_lcell_comb \Add10~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_remaining_samples[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add10~5_sumout ),
	.cout(\Add10~6 ),
	.shareout());
defparam \Add10~5 .extended_lut = "off";
defparam \Add10~5 .lut_mask = 64'h00000000000000FF;
defparam \Add10~5 .shared_arith = "off";

arriaii_lcell_comb \Selector125~0 (
	.dataa(!\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.datab(!\trk_block:sig_remaining_samples[1]~q ),
	.datac(!\trk_block:sig_trk_state.s_trk_idle~q ),
	.datad(!\Add10~5_sumout ),
	.datae(!\Selector121~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector125~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector125~0 .extended_lut = "off";
defparam \Selector125~0 .lut_mask = 64'h3131207531312075;
defparam \Selector125~0 .shared_arith = "off";

dffeas \trk_block:sig_remaining_samples[1] (
	.clk(clk),
	.d(\Selector125~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_dgrb_state.s_track~q ),
	.q(\trk_block:sig_remaining_samples[1]~q ),
	.prn(vcc));
defparam \trk_block:sig_remaining_samples[1] .is_wysiwyg = "true";
defparam \trk_block:sig_remaining_samples[1] .power_up = "low";

arriaii_lcell_comb \Add10~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_remaining_samples[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add10~9_sumout ),
	.cout(\Add10~10 ),
	.shareout());
defparam \Add10~9 .extended_lut = "off";
defparam \Add10~9 .lut_mask = 64'h00000000000000FF;
defparam \Add10~9 .shared_arith = "off";

arriaii_lcell_comb \Selector124~0 (
	.dataa(!\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.datab(!\trk_block:sig_remaining_samples[2]~q ),
	.datac(!\trk_block:sig_trk_state.s_trk_idle~q ),
	.datad(!\Add10~9_sumout ),
	.datae(!\Selector121~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector124~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector124~0 .extended_lut = "off";
defparam \Selector124~0 .lut_mask = 64'h3131207531312075;
defparam \Selector124~0 .shared_arith = "off";

dffeas \trk_block:sig_remaining_samples[2] (
	.clk(clk),
	.d(\Selector124~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_dgrb_state.s_track~q ),
	.q(\trk_block:sig_remaining_samples[2]~q ),
	.prn(vcc));
defparam \trk_block:sig_remaining_samples[2] .is_wysiwyg = "true";
defparam \trk_block:sig_remaining_samples[2] .power_up = "low";

arriaii_lcell_comb \Add10~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_remaining_samples[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add10~13_sumout ),
	.cout(\Add10~14 ),
	.shareout());
defparam \Add10~13 .extended_lut = "off";
defparam \Add10~13 .lut_mask = 64'h00000000000000FF;
defparam \Add10~13 .shared_arith = "off";

arriaii_lcell_comb \Selector123~0 (
	.dataa(!\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.datab(!\trk_block:sig_remaining_samples[3]~q ),
	.datac(!\trk_block:sig_trk_state.s_trk_idle~q ),
	.datad(!\Selector121~0_combout ),
	.datae(!\Add10~13_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector123~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector123~0 .extended_lut = "off";
defparam \Selector123~0 .lut_mask = 64'h3120317531203175;
defparam \Selector123~0 .shared_arith = "off";

dffeas \trk_block:sig_remaining_samples[3] (
	.clk(clk),
	.d(\Selector123~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_dgrb_state.s_track~q ),
	.q(\trk_block:sig_remaining_samples[3]~q ),
	.prn(vcc));
defparam \trk_block:sig_remaining_samples[3] .is_wysiwyg = "true";
defparam \trk_block:sig_remaining_samples[3] .power_up = "low";

arriaii_lcell_comb \Add10~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_remaining_samples[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add10~17_sumout ),
	.cout(\Add10~18 ),
	.shareout());
defparam \Add10~17 .extended_lut = "off";
defparam \Add10~17 .lut_mask = 64'h00000000000000FF;
defparam \Add10~17 .shared_arith = "off";

arriaii_lcell_comb \Selector122~0 (
	.dataa(!\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.datab(!\trk_block:sig_remaining_samples[4]~q ),
	.datac(!\trk_block:sig_trk_state.s_trk_idle~q ),
	.datad(!\Selector121~0_combout ),
	.datae(!\Add10~17_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector122~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector122~0 .extended_lut = "off";
defparam \Selector122~0 .lut_mask = 64'h3120317531203175;
defparam \Selector122~0 .shared_arith = "off";

dffeas \trk_block:sig_remaining_samples[4] (
	.clk(clk),
	.d(\Selector122~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_dgrb_state.s_track~q ),
	.q(\trk_block:sig_remaining_samples[4]~q ),
	.prn(vcc));
defparam \trk_block:sig_remaining_samples[4] .is_wysiwyg = "true";
defparam \trk_block:sig_remaining_samples[4] .power_up = "low";

arriaii_lcell_comb \Add10~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_remaining_samples[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add10~21_sumout ),
	.cout(\Add10~22 ),
	.shareout());
defparam \Add10~21 .extended_lut = "off";
defparam \Add10~21 .lut_mask = 64'h00000000000000FF;
defparam \Add10~21 .shared_arith = "off";

arriaii_lcell_comb \Selector121~1 (
	.dataa(!\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.datab(!\shift_in_mmc_seq_value~0_combout ),
	.datac(!\trk_block:sig_remaining_samples[5]~q ),
	.datad(!\Equal17~1_combout ),
	.datae(!\trk_block:sig_trk_state.s_trk_idle~q ),
	.dataf(!\Add10~21_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector121~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector121~1 .extended_lut = "off";
defparam \Selector121~1 .lut_mask = 64'h0E0EAEAE1F0EBFAE;
defparam \Selector121~1 .shared_arith = "off";

dffeas \trk_block:sig_remaining_samples[5] (
	.clk(clk),
	.d(\Selector121~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_dgrb_state.s_track~q ),
	.q(\trk_block:sig_remaining_samples[5]~q ),
	.prn(vcc));
defparam \trk_block:sig_remaining_samples[5] .is_wysiwyg = "true";
defparam \trk_block:sig_remaining_samples[5] .power_up = "low";

arriaii_lcell_comb \Add10~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_remaining_samples[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add10~25_sumout ),
	.cout(\Add10~26 ),
	.shareout());
defparam \Add10~25 .extended_lut = "off";
defparam \Add10~25 .lut_mask = 64'h00000000000000FF;
defparam \Add10~25 .shared_arith = "off";

arriaii_lcell_comb \Selector120~0 (
	.dataa(!\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.datab(!\trk_block:sig_remaining_samples[6]~q ),
	.datac(!\trk_block:sig_trk_state.s_trk_idle~q ),
	.datad(!\Selector121~0_combout ),
	.datae(!\Add10~25_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector120~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector120~0 .extended_lut = "off";
defparam \Selector120~0 .lut_mask = 64'h3120317531203175;
defparam \Selector120~0 .shared_arith = "off";

dffeas \trk_block:sig_remaining_samples[6] (
	.clk(clk),
	.d(\Selector120~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_dgrb_state.s_track~q ),
	.q(\trk_block:sig_remaining_samples[6]~q ),
	.prn(vcc));
defparam \trk_block:sig_remaining_samples[6] .is_wysiwyg = "true";
defparam \trk_block:sig_remaining_samples[6] .power_up = "low";

arriaii_lcell_comb \Add10~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_remaining_samples[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add10~29_sumout ),
	.cout(),
	.shareout());
defparam \Add10~29 .extended_lut = "off";
defparam \Add10~29 .lut_mask = 64'h00000000000000FF;
defparam \Add10~29 .shared_arith = "off";

arriaii_lcell_comb \Selector119~0 (
	.dataa(!\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.datab(!\trk_block:sig_remaining_samples[7]~q ),
	.datac(!\trk_block:sig_trk_state.s_trk_idle~q ),
	.datad(!\Selector121~0_combout ),
	.datae(!\Add10~29_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector119~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector119~0 .extended_lut = "off";
defparam \Selector119~0 .lut_mask = 64'h3120317531203175;
defparam \Selector119~0 .shared_arith = "off";

dffeas \trk_block:sig_remaining_samples[7] (
	.clk(clk),
	.d(\Selector119~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_dgrb_state.s_track~q ),
	.q(\trk_block:sig_remaining_samples[7]~q ),
	.prn(vcc));
defparam \trk_block:sig_remaining_samples[7] .is_wysiwyg = "true";
defparam \trk_block:sig_remaining_samples[7] .power_up = "low";

arriaii_lcell_comb \Equal17~0 (
	.dataa(!\trk_block:sig_remaining_samples[4]~q ),
	.datab(!\trk_block:sig_remaining_samples[5]~q ),
	.datac(!\trk_block:sig_remaining_samples[7]~q ),
	.datad(!\trk_block:sig_remaining_samples[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal17~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal17~0 .extended_lut = "off";
defparam \Equal17~0 .lut_mask = 64'h8000800080008000;
defparam \Equal17~0 .shared_arith = "off";

arriaii_lcell_comb \Equal17~1 (
	.dataa(!\trk_block:sig_remaining_samples[2]~q ),
	.datab(!\trk_block:sig_remaining_samples[3]~q ),
	.datac(!\Equal17~0_combout ),
	.datad(!\trk_block:sig_remaining_samples[1]~q ),
	.datae(!\trk_block:sig_remaining_samples[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal17~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal17~1 .extended_lut = "off";
defparam \Equal17~1 .lut_mask = 64'h0800000008000000;
defparam \Equal17~1 .shared_arith = "off";

arriaii_lcell_comb \sig_trk_state~14 (
	.dataa(!sig_addr_cmd0cke0),
	.datab(!\trk_block:sig_trk_last_state.s_trk_cdvw_calc~q ),
	.datac(!\trk_block:sig_trk_state.s_trk_cdvw_calc~q ),
	.datad(!\trk_block:sig_trk_state.s_trk_idle~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_trk_state~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_trk_state~14 .extended_lut = "off";
defparam \sig_trk_state~14 .lut_mask = 64'h5400540054005400;
defparam \sig_trk_state~14 .shared_arith = "off";

arriaii_lcell_comb \sig_trk_state~15 (
	.dataa(!\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.datab(!\shift_in_mmc_seq_value~0_combout ),
	.datac(!\Equal17~1_combout ),
	.datad(!\sig_trk_state~14_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_trk_state~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_trk_state~15 .extended_lut = "off";
defparam \sig_trk_state~15 .lut_mask = 64'h00EA00EA00EA00EA;
defparam \sig_trk_state~15 .shared_arith = "off";

arriaii_lcell_comb \Selector88~0 (
	.dataa(!\trk_block:sig_trk_state.s_trk_next_phase~q ),
	.datab(!\sig_phs_shft_end~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector88~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector88~0 .extended_lut = "off";
defparam \Selector88~0 .lut_mask = 64'h1111111111111111;
defparam \Selector88~0 .shared_arith = "off";

arriaii_lcell_comb \sig_trk_state~16 (
	.dataa(!\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.datab(!\sig_cdvw_state.status.calculating~q ),
	.datac(!\sig_trk_state~15_combout ),
	.datad(!\Selector88~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_trk_state~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_trk_state~16 .extended_lut = "off";
defparam \sig_trk_state~16 .lut_mask = 64'h0B010B010B010B01;
defparam \sig_trk_state~16 .shared_arith = "off";

arriaii_lcell_comb \Selector95~0 (
	.dataa(!sig_addr_cmd0cke0),
	.datab(!\sig_cdvw_state.status.valid_result~q ),
	.datac(!\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.datad(!\sig_cdvw_state.status.calculating~q ),
	.datae(!\trk_block:sig_mimic_cdv_found~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector95~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector95~0 .extended_lut = "off";
defparam \Selector95~0 .lut_mask = 64'h03005F5F03005F5F;
defparam \Selector95~0 .shared_arith = "off";

dffeas \trk_block:sig_mimic_cdv_found (
	.clk(clk),
	.d(\Selector95~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_dgrb_state.s_track~q ),
	.q(\trk_block:sig_mimic_cdv_found~q ),
	.prn(vcc));
defparam \trk_block:sig_mimic_cdv_found .is_wysiwyg = "true";
defparam \trk_block:sig_mimic_cdv_found .power_up = "low";

arriaii_lcell_comb \Selector128~2 (
	.dataa(!\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.datab(!\sig_cdvw_state.status.calculating~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector128~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector128~2 .extended_lut = "off";
defparam \Selector128~2 .lut_mask = 64'h4444444444444444;
defparam \Selector128~2 .shared_arith = "off";

arriaii_lcell_comb \Selector88~1 (
	.dataa(!\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.datab(!\shift_in_mmc_seq_value~0_combout ),
	.datac(!\Equal17~1_combout ),
	.datad(!\trk_block:sig_trk_state.s_trk_idle~q ),
	.datae(!\Selector88~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector88~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector88~1 .extended_lut = "off";
defparam \Selector88~1 .lut_mask = 64'h40FFFFFF40FFFFFF;
defparam \Selector88~1 .shared_arith = "off";

dffeas \trk_block:sig_trk_state.s_trk_mimic_sample (
	.clk(clk),
	.d(\Selector88~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_track~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.prn(vcc));
defparam \trk_block:sig_trk_state.s_trk_mimic_sample .is_wysiwyg = "true";
defparam \trk_block:sig_trk_state.s_trk_mimic_sample .power_up = "low";

arriaii_lcell_comb \sig_trk_state~21 (
	.dataa(!\trk_block:sig_trk_state.s_trk_next_phase~q ),
	.datab(!\sig_phs_shft_end~q ),
	.datac(!\trk_block:sig_trk_last_state.s_trk_cdvw_drift~q ),
	.datad(!\trk_block:sig_trk_state.s_trk_cdvw_drift~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_trk_state~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_trk_state~21 .extended_lut = "off";
defparam \sig_trk_state~21 .lut_mask = 64'h110F110F110F110F;
defparam \sig_trk_state~21 .shared_arith = "off";

arriaii_lcell_comb \sig_trk_state~22 (
	.dataa(!\sig_cdvw_state.status.valid_result~q ),
	.datab(!\Selector128~2_combout ),
	.datac(!\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.datad(!\sig_trk_state~15_combout ),
	.datae(!\sig_trk_state~21_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_trk_state~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_trk_state~22 .extended_lut = "off";
defparam \sig_trk_state~22 .lut_mask = 64'h11DD111D11DD111D;
defparam \sig_trk_state~22 .shared_arith = "off";

arriaii_lcell_comb \sig_trk_state~25 (
	.dataa(!\Selector128~2_combout ),
	.datab(!\trk_block:sig_trk_state.s_trk_cdvw_drift~q ),
	.datac(!\trk_block:sig_mimic_cdv_found~q ),
	.datad(!\sig_trk_state~17_combout ),
	.datae(!\sig_trk_state~22_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_trk_state~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_trk_state~25 .extended_lut = "off";
defparam \sig_trk_state~25 .lut_mask = 64'h0000002700000027;
defparam \sig_trk_state~25 .shared_arith = "off";

dffeas \trk_block:sig_trk_state.s_trk_cdvw_drift (
	.clk(clk),
	.d(\sig_trk_state~25_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_trk_state.s_trk_cdvw_drift~q ),
	.prn(vcc));
defparam \trk_block:sig_trk_state.s_trk_cdvw_drift .is_wysiwyg = "true";
defparam \trk_block:sig_trk_state.s_trk_cdvw_drift .power_up = "low";

arriaii_lcell_comb \sig_trk_last_state~0 (
	.dataa(!\sig_dgrb_state.s_track~q ),
	.datab(!\trk_block:sig_trk_state.s_trk_cdvw_drift~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_trk_last_state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_trk_last_state~0 .extended_lut = "off";
defparam \sig_trk_last_state~0 .lut_mask = 64'h1111111111111111;
defparam \sig_trk_last_state~0 .shared_arith = "off";

dffeas \trk_block:sig_trk_last_state.s_trk_cdvw_drift (
	.clk(clk),
	.d(\sig_trk_last_state~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_trk_last_state.s_trk_cdvw_drift~q ),
	.prn(vcc));
defparam \trk_block:sig_trk_last_state.s_trk_cdvw_drift .is_wysiwyg = "true";
defparam \trk_block:sig_trk_last_state.s_trk_cdvw_drift .power_up = "low";

arriaii_lcell_comb \trk_block:sig_req_rsc_shift[5]~0 (
	.dataa(!\sig_dgrb_state.s_track~q ),
	.datab(!\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.datac(!sig_addr_cmd0cke0),
	.datad(!\trk_block:sig_trk_last_state.s_trk_cdvw_drift~q ),
	.datae(!\trk_block:sig_trk_state.s_trk_cdvw_drift~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\trk_block:sig_req_rsc_shift[5]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \trk_block:sig_req_rsc_shift[5]~0 .extended_lut = "off";
defparam \trk_block:sig_req_rsc_shift[5]~0 .lut_mask = 64'h5151005551510055;
defparam \trk_block:sig_req_rsc_shift[5]~0 .shared_arith = "off";

arriaii_lcell_comb \sig_req_rsc_shift~2 (
	.dataa(!\trk_block:sig_trk_last_state.s_trk_adjust_resync~q ),
	.datab(!\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.datac(!\trk_block:sig_mimic_cdv_found~q ),
	.datad(!\trk_block:sig_req_rsc_shift[5]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_req_rsc_shift~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_req_rsc_shift~2 .extended_lut = "off";
defparam \sig_req_rsc_shift~2 .lut_mask = 64'h0F010F010F010F01;
defparam \sig_req_rsc_shift~2 .shared_arith = "off";

arriaii_lcell_comb \trk_block:sig_mimic_cdv[5]~0 (
	.dataa(!\sig_dgrb_state.s_track~q ),
	.datab(!\sig_cdvw_state.status.valid_result~q ),
	.datac(!\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\trk_block:sig_mimic_cdv[5]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \trk_block:sig_mimic_cdv[5]~0 .extended_lut = "off";
defparam \trk_block:sig_mimic_cdv[5]~0 .lut_mask = 64'h0101010101010101;
defparam \trk_block:sig_mimic_cdv[5]~0 .shared_arith = "off";

dffeas \trk_block:sig_mimic_cdv[0] (
	.clk(clk),
	.d(\sig_cdvw_state.largest_window_centre[0]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\trk_block:sig_mimic_cdv[5]~0_combout ),
	.q(\trk_block:sig_mimic_cdv[0]~q ),
	.prn(vcc));
defparam \trk_block:sig_mimic_cdv[0] .is_wysiwyg = "true";
defparam \trk_block:sig_mimic_cdv[0] .power_up = "low";

arriaii_lcell_comb \Add11~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\trk_block:sig_mimic_cdv[0]~q ),
	.datad(!\sig_cdvw_state.largest_window_centre[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add11~1_sumout ),
	.cout(\Add11~2 ),
	.shareout(\Add11~3 ));
defparam \Add11~1 .extended_lut = "off";
defparam \Add11~1 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add11~1 .shared_arith = "on";

arriaii_lcell_comb \sig_mimic_delta~7 (
	.dataa(!\sig_cdvw_state.status.valid_result~q ),
	.datab(!\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.datac(!\trk_block:sig_mimic_cdv_found~q ),
	.datad(!\Add11~1_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_mimic_delta~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_mimic_delta~7 .extended_lut = "off";
defparam \sig_mimic_delta~7 .lut_mask = 64'h0001000100010001;
defparam \sig_mimic_delta~7 .shared_arith = "off";

arriaii_lcell_comb \sig_mimic_delta~1 (
	.dataa(!\sig_dgrb_state.s_track~q ),
	.datab(!sig_addr_cmd0cke0),
	.datac(!\sig_cdvw_state.status.valid_result~q ),
	.datad(!\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.datae(!\trk_block:sig_mimic_cdv_found~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_mimic_delta~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_mimic_delta~1 .extended_lut = "off";
defparam \sig_mimic_delta~1 .lut_mask = 64'hFFFF4405FFFF4405;
defparam \sig_mimic_delta~1 .shared_arith = "off";

dffeas \trk_block:sig_mimic_delta[0] (
	.clk(clk),
	.d(\sig_mimic_delta~7_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_track~q ),
	.sload(gnd),
	.ena(\sig_mimic_delta~1_combout ),
	.q(\trk_block:sig_mimic_delta[0]~q ),
	.prn(vcc));
defparam \trk_block:sig_mimic_delta[0] .is_wysiwyg = "true";
defparam \trk_block:sig_mimic_delta[0] .power_up = "low";

arriaii_lcell_comb \Add15~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_mimic_delta[0]~q ),
	.datae(gnd),
	.dataf(!\trk_block:sig_req_rsc_shift[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add15~1_sumout ),
	.cout(\Add15~2 ),
	.shareout());
defparam \Add15~1 .extended_lut = "off";
defparam \Add15~1 .lut_mask = 64'h000000FF000000FF;
defparam \Add15~1 .shared_arith = "off";

arriaii_lcell_comb \sig_trk_state~12 (
	.dataa(!\trk_block:sig_trk_last_state.s_trk_cdvw_drift~q ),
	.datab(!\trk_block:sig_trk_state.s_trk_cdvw_drift~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_trk_state~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_trk_state~12 .extended_lut = "off";
defparam \sig_trk_state~12 .lut_mask = 64'h1111111111111111;
defparam \sig_trk_state~12 .shared_arith = "off";

arriaii_lcell_comb \Add18~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_req_rsc_shift[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add18~1_sumout ),
	.cout(\Add18~2 ),
	.shareout());
defparam \Add18~1 .extended_lut = "off";
defparam \Add18~1 .lut_mask = 64'h000000000000FF00;
defparam \Add18~1 .shared_arith = "off";

arriaii_lcell_comb \Add18~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_req_rsc_shift[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add18~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add18~5_sumout ),
	.cout(\Add18~6 ),
	.shareout());
defparam \Add18~5 .extended_lut = "off";
defparam \Add18~5 .lut_mask = 64'h00000000000000FF;
defparam \Add18~5 .shared_arith = "off";

arriaii_lcell_comb \Add16~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_req_rsc_shift[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add16~1_sumout ),
	.cout(\Add16~2 ),
	.shareout());
defparam \Add16~1 .extended_lut = "off";
defparam \Add16~1 .lut_mask = 64'h000000000000FF00;
defparam \Add16~1 .shared_arith = "off";

arriaii_lcell_comb \Add16~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_req_rsc_shift[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add16~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add16~5_sumout ),
	.cout(\Add16~6 ),
	.shareout());
defparam \Add16~5 .extended_lut = "off";
defparam \Add16~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add16~5 .shared_arith = "off";

arriaii_lcell_comb \trk_block:sig_req_rsc_shift[5]~1 (
	.dataa(!\trk_block:sig_trk_last_state.s_trk_adjust_resync~q ),
	.datab(!\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.datac(!\sig_trk_state~11_combout ),
	.datad(!\trk_block:sig_req_rsc_shift[5]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\trk_block:sig_req_rsc_shift[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \trk_block:sig_req_rsc_shift[5]~1 .extended_lut = "off";
defparam \trk_block:sig_req_rsc_shift[5]~1 .lut_mask = 64'h00EC00EC00EC00EC;
defparam \trk_block:sig_req_rsc_shift[5]~1 .shared_arith = "off";

arriaii_lcell_comb \trk_block:sig_req_rsc_shift[5]~2 (
	.dataa(!\trk_block:sig_req_rsc_shift[7]~q ),
	.datab(!\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.datac(!\trk_block:sig_trk_state.s_trk_cdvw_drift~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\trk_block:sig_req_rsc_shift[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \trk_block:sig_req_rsc_shift[5]~2 .extended_lut = "off";
defparam \trk_block:sig_req_rsc_shift[5]~2 .lut_mask = 64'h1D1D1D1D1D1D1D1D;
defparam \trk_block:sig_req_rsc_shift[5]~2 .shared_arith = "off";

arriaii_lcell_comb \trk_block:sig_req_rsc_shift[5]~3 (
	.dataa(!\trk_block:sig_req_rsc_shift[7]~q ),
	.datab(!\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.datac(!\trk_block:sig_trk_state.s_trk_cdvw_drift~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\trk_block:sig_req_rsc_shift[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \trk_block:sig_req_rsc_shift[5]~3 .extended_lut = "off";
defparam \trk_block:sig_req_rsc_shift[5]~3 .lut_mask = 64'h2E2E2E2E2E2E2E2E;
defparam \trk_block:sig_req_rsc_shift[5]~3 .shared_arith = "off";

arriaii_lcell_comb \sig_req_rsc_shift~5 (
	.dataa(!\Add15~5_sumout ),
	.datab(!\Add18~5_sumout ),
	.datac(!\Add16~5_sumout ),
	.datad(!\trk_block:sig_req_rsc_shift[5]~1_combout ),
	.datae(!\trk_block:sig_req_rsc_shift[5]~2_combout ),
	.dataf(!\trk_block:sig_req_rsc_shift[5]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_req_rsc_shift~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_req_rsc_shift~5 .extended_lut = "off";
defparam \sig_req_rsc_shift~5 .lut_mask = 64'h00000033000F0055;
defparam \sig_req_rsc_shift~5 .shared_arith = "off";

arriaii_lcell_comb \Add18~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_req_rsc_shift[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add18~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add18~9_sumout ),
	.cout(\Add18~10 ),
	.shareout());
defparam \Add18~9 .extended_lut = "off";
defparam \Add18~9 .lut_mask = 64'h00000000000000FF;
defparam \Add18~9 .shared_arith = "off";

arriaii_lcell_comb \Add16~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_req_rsc_shift[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add16~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add16~9_sumout ),
	.cout(\Add16~10 ),
	.shareout());
defparam \Add16~9 .extended_lut = "off";
defparam \Add16~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add16~9 .shared_arith = "off";

arriaii_lcell_comb \sig_req_rsc_shift~6 (
	.dataa(!\Add15~9_sumout ),
	.datab(!\Add18~9_sumout ),
	.datac(!\Add16~9_sumout ),
	.datad(!\trk_block:sig_req_rsc_shift[5]~1_combout ),
	.datae(!\trk_block:sig_req_rsc_shift[5]~2_combout ),
	.dataf(!\trk_block:sig_req_rsc_shift[5]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_req_rsc_shift~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_req_rsc_shift~6 .extended_lut = "off";
defparam \sig_req_rsc_shift~6 .lut_mask = 64'h00000033000F0055;
defparam \sig_req_rsc_shift~6 .shared_arith = "off";

dffeas \trk_block:sig_req_rsc_shift[2] (
	.clk(clk),
	.d(\sig_req_rsc_shift~6_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\trk_block:sig_req_rsc_shift[5]~4_combout ),
	.q(\trk_block:sig_req_rsc_shift[2]~q ),
	.prn(vcc));
defparam \trk_block:sig_req_rsc_shift[2] .is_wysiwyg = "true";
defparam \trk_block:sig_req_rsc_shift[2] .power_up = "low";

arriaii_lcell_comb \Add18~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_req_rsc_shift[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add18~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add18~13_sumout ),
	.cout(\Add18~14 ),
	.shareout());
defparam \Add18~13 .extended_lut = "off";
defparam \Add18~13 .lut_mask = 64'h00000000000000FF;
defparam \Add18~13 .shared_arith = "off";

arriaii_lcell_comb \Add16~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_req_rsc_shift[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add16~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add16~13_sumout ),
	.cout(\Add16~14 ),
	.shareout());
defparam \Add16~13 .extended_lut = "off";
defparam \Add16~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add16~13 .shared_arith = "off";

arriaii_lcell_comb \sig_req_rsc_shift~7 (
	.dataa(!\Add15~13_sumout ),
	.datab(!\Add18~13_sumout ),
	.datac(!\Add16~13_sumout ),
	.datad(!\trk_block:sig_req_rsc_shift[5]~1_combout ),
	.datae(!\trk_block:sig_req_rsc_shift[5]~2_combout ),
	.dataf(!\trk_block:sig_req_rsc_shift[5]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_req_rsc_shift~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_req_rsc_shift~7 .extended_lut = "off";
defparam \sig_req_rsc_shift~7 .lut_mask = 64'h00000033000F0055;
defparam \sig_req_rsc_shift~7 .shared_arith = "off";

dffeas \trk_block:sig_req_rsc_shift[3] (
	.clk(clk),
	.d(\sig_req_rsc_shift~7_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\trk_block:sig_req_rsc_shift[5]~4_combout ),
	.q(\trk_block:sig_req_rsc_shift[3]~q ),
	.prn(vcc));
defparam \trk_block:sig_req_rsc_shift[3] .is_wysiwyg = "true";
defparam \trk_block:sig_req_rsc_shift[3] .power_up = "low";

arriaii_lcell_comb \Add18~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_req_rsc_shift[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add18~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add18~17_sumout ),
	.cout(\Add18~18 ),
	.shareout());
defparam \Add18~17 .extended_lut = "off";
defparam \Add18~17 .lut_mask = 64'h00000000000000FF;
defparam \Add18~17 .shared_arith = "off";

arriaii_lcell_comb \Add16~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_req_rsc_shift[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add16~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add16~17_sumout ),
	.cout(\Add16~18 ),
	.shareout());
defparam \Add16~17 .extended_lut = "off";
defparam \Add16~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add16~17 .shared_arith = "off";

arriaii_lcell_comb \sig_req_rsc_shift~8 (
	.dataa(!\Add15~17_sumout ),
	.datab(!\Add18~17_sumout ),
	.datac(!\Add16~17_sumout ),
	.datad(!\trk_block:sig_req_rsc_shift[5]~1_combout ),
	.datae(!\trk_block:sig_req_rsc_shift[5]~2_combout ),
	.dataf(!\trk_block:sig_req_rsc_shift[5]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_req_rsc_shift~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_req_rsc_shift~8 .extended_lut = "off";
defparam \sig_req_rsc_shift~8 .lut_mask = 64'h00000033000F0055;
defparam \sig_req_rsc_shift~8 .shared_arith = "off";

dffeas \trk_block:sig_req_rsc_shift[4] (
	.clk(clk),
	.d(\sig_req_rsc_shift~8_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\trk_block:sig_req_rsc_shift[5]~4_combout ),
	.q(\trk_block:sig_req_rsc_shift[4]~q ),
	.prn(vcc));
defparam \trk_block:sig_req_rsc_shift[4] .is_wysiwyg = "true";
defparam \trk_block:sig_req_rsc_shift[4] .power_up = "low";

arriaii_lcell_comb \trk_block:sig_req_rsc_shift[5]~5 (
	.dataa(!\trk_block:sig_req_rsc_shift[7]~q ),
	.datab(!\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.datac(!\trk_block:sig_req_rsc_shift[5]~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\trk_block:sig_req_rsc_shift[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \trk_block:sig_req_rsc_shift[5]~5 .extended_lut = "off";
defparam \trk_block:sig_req_rsc_shift[5]~5 .lut_mask = 64'hF2F2F2F2F2F2F2F2;
defparam \trk_block:sig_req_rsc_shift[5]~5 .shared_arith = "off";

dffeas \trk_block:sig_mimic_cdv[4] (
	.clk(clk),
	.d(\sig_cdvw_state.largest_window_centre[4]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\trk_block:sig_mimic_cdv[5]~0_combout ),
	.q(\trk_block:sig_mimic_cdv[4]~q ),
	.prn(vcc));
defparam \trk_block:sig_mimic_cdv[4] .is_wysiwyg = "true";
defparam \trk_block:sig_mimic_cdv[4] .power_up = "low";

dffeas \trk_block:sig_mimic_cdv[3] (
	.clk(clk),
	.d(\sig_cdvw_state.largest_window_centre[3]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\trk_block:sig_mimic_cdv[5]~0_combout ),
	.q(\trk_block:sig_mimic_cdv[3]~q ),
	.prn(vcc));
defparam \trk_block:sig_mimic_cdv[3] .is_wysiwyg = "true";
defparam \trk_block:sig_mimic_cdv[3] .power_up = "low";

dffeas \trk_block:sig_mimic_cdv[2] (
	.clk(clk),
	.d(\sig_cdvw_state.largest_window_centre[2]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\trk_block:sig_mimic_cdv[5]~0_combout ),
	.q(\trk_block:sig_mimic_cdv[2]~q ),
	.prn(vcc));
defparam \trk_block:sig_mimic_cdv[2] .is_wysiwyg = "true";
defparam \trk_block:sig_mimic_cdv[2] .power_up = "low";

dffeas \trk_block:sig_mimic_cdv[1] (
	.clk(clk),
	.d(\sig_cdvw_state.largest_window_centre[1]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\trk_block:sig_mimic_cdv[5]~0_combout ),
	.q(\trk_block:sig_mimic_cdv[1]~q ),
	.prn(vcc));
defparam \trk_block:sig_mimic_cdv[1] .is_wysiwyg = "true";
defparam \trk_block:sig_mimic_cdv[1] .power_up = "low";

arriaii_lcell_comb \Add11~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\trk_block:sig_mimic_cdv[1]~q ),
	.datad(!\sig_cdvw_state.largest_window_centre[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add11~2 ),
	.sharein(\Add11~3 ),
	.combout(),
	.sumout(\Add11~5_sumout ),
	.cout(\Add11~6 ),
	.shareout(\Add11~7 ));
defparam \Add11~5 .extended_lut = "off";
defparam \Add11~5 .lut_mask = 64'h00000F000000F00F;
defparam \Add11~5 .shared_arith = "on";

arriaii_lcell_comb \Add11~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\trk_block:sig_mimic_cdv[2]~q ),
	.datad(!\sig_cdvw_state.largest_window_centre[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add11~6 ),
	.sharein(\Add11~7 ),
	.combout(),
	.sumout(\Add11~9_sumout ),
	.cout(\Add11~10 ),
	.shareout(\Add11~11 ));
defparam \Add11~9 .extended_lut = "off";
defparam \Add11~9 .lut_mask = 64'h00000F000000F00F;
defparam \Add11~9 .shared_arith = "on";

arriaii_lcell_comb \Add11~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\trk_block:sig_mimic_cdv[3]~q ),
	.datad(!\sig_cdvw_state.largest_window_centre[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add11~10 ),
	.sharein(\Add11~11 ),
	.combout(),
	.sumout(\Add11~13_sumout ),
	.cout(\Add11~14 ),
	.shareout(\Add11~15 ));
defparam \Add11~13 .extended_lut = "off";
defparam \Add11~13 .lut_mask = 64'h00000F000000F00F;
defparam \Add11~13 .shared_arith = "on";

arriaii_lcell_comb \Add11~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\trk_block:sig_mimic_cdv[4]~q ),
	.datad(!\sig_cdvw_state.largest_window_centre[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add11~14 ),
	.sharein(\Add11~15 ),
	.combout(),
	.sumout(\Add11~17_sumout ),
	.cout(\Add11~18 ),
	.shareout(\Add11~19 ));
defparam \Add11~17 .extended_lut = "off";
defparam \Add11~17 .lut_mask = 64'h00000F000000F00F;
defparam \Add11~17 .shared_arith = "on";

arriaii_lcell_comb \sig_mimic_delta~3 (
	.dataa(!\sig_cdvw_state.status.valid_result~q ),
	.datab(!\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.datac(!\trk_block:sig_mimic_cdv_found~q ),
	.datad(!\Add11~17_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_mimic_delta~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_mimic_delta~3 .extended_lut = "off";
defparam \sig_mimic_delta~3 .lut_mask = 64'h0001000100010001;
defparam \sig_mimic_delta~3 .shared_arith = "off";

dffeas \trk_block:sig_mimic_delta[4] (
	.clk(clk),
	.d(\sig_mimic_delta~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_track~q ),
	.sload(gnd),
	.ena(\sig_mimic_delta~1_combout ),
	.q(\trk_block:sig_mimic_delta[4]~q ),
	.prn(vcc));
defparam \trk_block:sig_mimic_delta[4] .is_wysiwyg = "true";
defparam \trk_block:sig_mimic_delta[4] .power_up = "low";

arriaii_lcell_comb \sig_mimic_delta~4 (
	.dataa(!\sig_cdvw_state.status.valid_result~q ),
	.datab(!\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.datac(!\trk_block:sig_mimic_cdv_found~q ),
	.datad(!\Add11~13_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_mimic_delta~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_mimic_delta~4 .extended_lut = "off";
defparam \sig_mimic_delta~4 .lut_mask = 64'h0001000100010001;
defparam \sig_mimic_delta~4 .shared_arith = "off";

dffeas \trk_block:sig_mimic_delta[3] (
	.clk(clk),
	.d(\sig_mimic_delta~4_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_track~q ),
	.sload(gnd),
	.ena(\sig_mimic_delta~1_combout ),
	.q(\trk_block:sig_mimic_delta[3]~q ),
	.prn(vcc));
defparam \trk_block:sig_mimic_delta[3] .is_wysiwyg = "true";
defparam \trk_block:sig_mimic_delta[3] .power_up = "low";

arriaii_lcell_comb \sig_mimic_delta~5 (
	.dataa(!\sig_cdvw_state.status.valid_result~q ),
	.datab(!\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.datac(!\trk_block:sig_mimic_cdv_found~q ),
	.datad(!\Add11~9_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_mimic_delta~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_mimic_delta~5 .extended_lut = "off";
defparam \sig_mimic_delta~5 .lut_mask = 64'h0001000100010001;
defparam \sig_mimic_delta~5 .shared_arith = "off";

dffeas \trk_block:sig_mimic_delta[2] (
	.clk(clk),
	.d(\sig_mimic_delta~5_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_track~q ),
	.sload(gnd),
	.ena(\sig_mimic_delta~1_combout ),
	.q(\trk_block:sig_mimic_delta[2]~q ),
	.prn(vcc));
defparam \trk_block:sig_mimic_delta[2] .is_wysiwyg = "true";
defparam \trk_block:sig_mimic_delta[2] .power_up = "low";

arriaii_lcell_comb \sig_mimic_delta~6 (
	.dataa(!\sig_cdvw_state.status.valid_result~q ),
	.datab(!\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.datac(!\trk_block:sig_mimic_cdv_found~q ),
	.datad(!\Add11~5_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_mimic_delta~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_mimic_delta~6 .extended_lut = "off";
defparam \sig_mimic_delta~6 .lut_mask = 64'h0001000100010001;
defparam \sig_mimic_delta~6 .shared_arith = "off";

dffeas \trk_block:sig_mimic_delta[1] (
	.clk(clk),
	.d(\sig_mimic_delta~6_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_track~q ),
	.sload(gnd),
	.ena(\sig_mimic_delta~1_combout ),
	.q(\trk_block:sig_mimic_delta[1]~q ),
	.prn(vcc));
defparam \trk_block:sig_mimic_delta[1] .is_wysiwyg = "true";
defparam \trk_block:sig_mimic_delta[1] .power_up = "low";

arriaii_lcell_comb \Add12~5 (
	.dataa(!\trk_block:sig_mimic_delta[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_mimic_delta[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add12~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~5_sumout ),
	.cout(\Add12~6 ),
	.shareout());
defparam \Add12~5 .extended_lut = "off";
defparam \Add12~5 .lut_mask = 64'h0000FFFF0000AA55;
defparam \Add12~5 .shared_arith = "off";

arriaii_lcell_comb \Add12~9 (
	.dataa(!\trk_block:sig_mimic_delta[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_mimic_delta[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add12~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~9_sumout ),
	.cout(\Add12~10 ),
	.shareout());
defparam \Add12~9 .extended_lut = "off";
defparam \Add12~9 .lut_mask = 64'h0000FFFF0000AA55;
defparam \Add12~9 .shared_arith = "off";

arriaii_lcell_comb \Add12~17 (
	.dataa(!\trk_block:sig_mimic_delta[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_mimic_delta[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add12~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~17_sumout ),
	.cout(\Add12~18 ),
	.shareout());
defparam \Add12~17 .extended_lut = "off";
defparam \Add12~17 .lut_mask = 64'h0000FFFF0000AA55;
defparam \Add12~17 .shared_arith = "off";

dffeas \trk_block:sig_mimic_cdv[5] (
	.clk(clk),
	.d(\sig_cdvw_state.largest_window_centre[5]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\trk_block:sig_mimic_cdv[5]~0_combout ),
	.q(\trk_block:sig_mimic_cdv[5]~q ),
	.prn(vcc));
defparam \trk_block:sig_mimic_cdv[5] .is_wysiwyg = "true";
defparam \trk_block:sig_mimic_cdv[5] .power_up = "low";

arriaii_lcell_comb \Add11~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\trk_block:sig_mimic_cdv[5]~q ),
	.datad(!\sig_cdvw_state.largest_window_centre[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add11~18 ),
	.sharein(\Add11~19 ),
	.combout(),
	.sumout(\Add11~21_sumout ),
	.cout(\Add11~22 ),
	.shareout(\Add11~23 ));
defparam \Add11~21 .extended_lut = "off";
defparam \Add11~21 .lut_mask = 64'h00000F000000F00F;
defparam \Add11~21 .shared_arith = "on";

arriaii_lcell_comb \sig_mimic_delta~2 (
	.dataa(!\sig_dgrb_state.s_track~q ),
	.datab(!\sig_cdvw_state.status.valid_result~q ),
	.datac(!\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.datad(!\trk_block:sig_mimic_cdv_found~q ),
	.datae(!\Add11~21_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_mimic_delta~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_mimic_delta~2 .extended_lut = "off";
defparam \sig_mimic_delta~2 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \sig_mimic_delta~2 .shared_arith = "off";

dffeas \trk_block:sig_mimic_delta[5] (
	.clk(clk),
	.d(\sig_mimic_delta~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_mimic_delta~1_combout ),
	.q(\trk_block:sig_mimic_delta[5]~q ),
	.prn(vcc));
defparam \trk_block:sig_mimic_delta[5] .is_wysiwyg = "true";
defparam \trk_block:sig_mimic_delta[5] .power_up = "low";

arriaii_lcell_comb \Add12~21 (
	.dataa(!\trk_block:sig_mimic_delta[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_mimic_delta[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add12~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~21_sumout ),
	.cout(\Add12~22 ),
	.shareout());
defparam \Add12~21 .extended_lut = "off";
defparam \Add12~21 .lut_mask = 64'h0000FFFF000055AA;
defparam \Add12~21 .shared_arith = "off";

arriaii_lcell_comb \Add12~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add12~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add12~25_sumout ),
	.cout(),
	.shareout());
defparam \Add12~25 .extended_lut = "off";
defparam \Add12~25 .lut_mask = 64'h0000FFFF00000000;
defparam \Add12~25 .shared_arith = "off";

arriaii_lcell_comb \LessThan8~0 (
	.dataa(!\Add12~1_sumout ),
	.datab(!\Add12~5_sumout ),
	.datac(!\Add12~9_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan8~0 .extended_lut = "off";
defparam \LessThan8~0 .lut_mask = 64'h8080808080808080;
defparam \LessThan8~0 .shared_arith = "off";

arriaii_lcell_comb \LessThan8~1 (
	.dataa(!\Add12~13_sumout ),
	.datab(!\Add12~17_sumout ),
	.datac(!\Add12~21_sumout ),
	.datad(!\Add12~25_sumout ),
	.datae(!\LessThan8~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan8~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan8~1 .extended_lut = "off";
defparam \LessThan8~1 .lut_mask = 64'h3FFF1FFF3FFF1FFF;
defparam \LessThan8~1 .shared_arith = "off";

dffeas \trk_block:sig_large_drift_seen (
	.clk(clk),
	.d(\LessThan8~1_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_track~q ),
	.sload(!\trk_block:sig_trk_state.s_trk_cdvw_drift~q ),
	.ena(vcc),
	.q(\trk_block:sig_large_drift_seen~q ),
	.prn(vcc));
defparam \trk_block:sig_large_drift_seen .is_wysiwyg = "true";
defparam \trk_block:sig_large_drift_seen .power_up = "low";

arriaii_lcell_comb \trk_block:sig_req_rsc_shift[5]~6 (
	.dataa(!\trk_block:sig_req_rsc_shift[7]~q ),
	.datab(!\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.datac(!\trk_block:sig_large_drift_seen~q ),
	.datad(!\trk_block:sig_trk_state.s_trk_cdvw_drift~q ),
	.datae(!\trk_block:sig_req_rsc_shift[5]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\trk_block:sig_req_rsc_shift[5]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \trk_block:sig_req_rsc_shift[5]~6 .extended_lut = "off";
defparam \trk_block:sig_req_rsc_shift[5]~6 .lut_mask = 64'hFFFFDD0DFFFFDD0D;
defparam \trk_block:sig_req_rsc_shift[5]~6 .shared_arith = "off";

arriaii_lcell_comb \Add15~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_mimic_delta[5]~q ),
	.datae(gnd),
	.dataf(!\trk_block:sig_req_rsc_shift[5]~q ),
	.datag(gnd),
	.cin(\Add15~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add15~21_sumout ),
	.cout(\Add15~22 ),
	.shareout());
defparam \Add15~21 .extended_lut = "off";
defparam \Add15~21 .lut_mask = 64'h0000FF000000FF00;
defparam \Add15~21 .shared_arith = "off";

arriaii_lcell_comb \Add16~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_req_rsc_shift[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add16~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add16~21_sumout ),
	.cout(\Add16~22 ),
	.shareout());
defparam \Add16~21 .extended_lut = "off";
defparam \Add16~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add16~21 .shared_arith = "off";

arriaii_lcell_comb \sig_req_rsc_shift~12 (
	.dataa(!\Add18~21_sumout ),
	.datab(!\trk_block:sig_req_rsc_shift[5]~2_combout ),
	.datac(!\trk_block:sig_req_rsc_shift[5]~3_combout ),
	.datad(!\trk_block:sig_req_rsc_shift[5]~5_combout ),
	.datae(!\trk_block:sig_req_rsc_shift[5]~6_combout ),
	.dataf(!\Add15~21_sumout ),
	.datag(!\Add16~21_sumout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_req_rsc_shift~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_req_rsc_shift~12 .extended_lut = "on";
defparam \sig_req_rsc_shift~12 .lut_mask = 64'h000F1300FF0F1000;
defparam \sig_req_rsc_shift~12 .shared_arith = "off";

dffeas \trk_block:sig_req_rsc_shift[5] (
	.clk(clk),
	.d(\sig_req_rsc_shift~12_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\trk_block:sig_req_rsc_shift[5]~4_combout ),
	.q(\trk_block:sig_req_rsc_shift[5]~q ),
	.prn(vcc));
defparam \trk_block:sig_req_rsc_shift[5] .is_wysiwyg = "true";
defparam \trk_block:sig_req_rsc_shift[5] .power_up = "low";

arriaii_lcell_comb \Add16~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_req_rsc_shift[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add16~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add16~25_sumout ),
	.cout(\Add16~26 ),
	.shareout());
defparam \Add16~25 .extended_lut = "off";
defparam \Add16~25 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add16~25 .shared_arith = "off";

arriaii_lcell_comb \Add15~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_mimic_delta[6]~q ),
	.datae(gnd),
	.dataf(!\trk_block:sig_req_rsc_shift[6]~q ),
	.datag(gnd),
	.cin(\Add15~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add15~25_sumout ),
	.cout(\Add15~26 ),
	.shareout());
defparam \Add15~25 .extended_lut = "off";
defparam \Add15~25 .lut_mask = 64'h0000FF000000FF00;
defparam \Add15~25 .shared_arith = "off";

arriaii_lcell_comb \Add18~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_req_rsc_shift[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add18~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add18~25_sumout ),
	.cout(\Add18~26 ),
	.shareout());
defparam \Add18~25 .extended_lut = "off";
defparam \Add18~25 .lut_mask = 64'h00000000000000FF;
defparam \Add18~25 .shared_arith = "off";

arriaii_lcell_comb \sig_req_rsc_shift~9 (
	.dataa(!\trk_block:sig_mimic_delta[6]~q ),
	.datab(!\Add15~21_sumout ),
	.datac(!\Add15~25_sumout ),
	.datad(!\Add18~25_sumout ),
	.datae(!\trk_block:sig_req_rsc_shift[5]~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_req_rsc_shift~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_req_rsc_shift~9 .extended_lut = "off";
defparam \sig_req_rsc_shift~9 .lut_mask = 64'h00FF696900FF6969;
defparam \sig_req_rsc_shift~9 .shared_arith = "off";

arriaii_lcell_comb \sig_req_rsc_shift~10 (
	.dataa(!\Add15~25_sumout ),
	.datab(!\Add16~25_sumout ),
	.datac(!\trk_block:sig_req_rsc_shift[5]~2_combout ),
	.datad(!\sig_req_rsc_shift~9_combout ),
	.datae(!\trk_block:sig_req_rsc_shift[5]~5_combout ),
	.dataf(!\trk_block:sig_req_rsc_shift[5]~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_req_rsc_shift~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_req_rsc_shift~10 .extended_lut = "off";
defparam \sig_req_rsc_shift~10 .lut_mask = 64'h55553333000F0000;
defparam \sig_req_rsc_shift~10 .shared_arith = "off";

dffeas \trk_block:sig_req_rsc_shift[6] (
	.clk(clk),
	.d(\sig_req_rsc_shift~10_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\trk_block:sig_req_rsc_shift[5]~4_combout ),
	.q(\trk_block:sig_req_rsc_shift[6]~q ),
	.prn(vcc));
defparam \trk_block:sig_req_rsc_shift[6] .is_wysiwyg = "true";
defparam \trk_block:sig_req_rsc_shift[6] .power_up = "low";

arriaii_lcell_comb \LessThan11~0 (
	.dataa(!\trk_block:sig_req_rsc_shift[3]~q ),
	.datab(!\trk_block:sig_req_rsc_shift[4]~q ),
	.datac(!\trk_block:sig_req_rsc_shift[6]~q ),
	.datad(!\trk_block:sig_req_rsc_shift[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan11~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan11~0 .extended_lut = "off";
defparam \LessThan11~0 .lut_mask = 64'h8000800080008000;
defparam \LessThan11~0 .shared_arith = "off";

arriaii_lcell_comb \trk_block:sig_req_rsc_shift[5]~7 (
	.dataa(!\trk_block:sig_req_rsc_shift[7]~q ),
	.datab(!\trk_block:sig_req_rsc_shift[0]~q ),
	.datac(!\trk_block:sig_req_rsc_shift[1]~q ),
	.datad(!\trk_block:sig_req_rsc_shift[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\trk_block:sig_req_rsc_shift[5]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \trk_block:sig_req_rsc_shift[5]~7 .extended_lut = "off";
defparam \trk_block:sig_req_rsc_shift[5]~7 .lut_mask = 64'h1000100010001000;
defparam \trk_block:sig_req_rsc_shift[5]~7 .shared_arith = "off";

arriaii_lcell_comb \trk_block:sig_req_rsc_shift[5]~4 (
	.dataa(!\trk_block:sig_mimic_cdv_found~q ),
	.datab(!\trk_block:sig_trk_last_state.s_trk_adjust_resync~q ),
	.datac(!\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.datad(!\trk_block:sig_req_rsc_shift[5]~0_combout ),
	.datae(!\LessThan11~0_combout ),
	.dataf(!\trk_block:sig_req_rsc_shift[5]~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\trk_block:sig_req_rsc_shift[5]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \trk_block:sig_req_rsc_shift[5]~4 .extended_lut = "off";
defparam \trk_block:sig_req_rsc_shift[5]~4 .lut_mask = 64'hAAFEAAFEAAFEAAFA;
defparam \trk_block:sig_req_rsc_shift[5]~4 .shared_arith = "off";

dffeas \trk_block:sig_req_rsc_shift[1] (
	.clk(clk),
	.d(\sig_req_rsc_shift~5_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\trk_block:sig_req_rsc_shift[5]~4_combout ),
	.q(\trk_block:sig_req_rsc_shift[1]~q ),
	.prn(vcc));
defparam \trk_block:sig_req_rsc_shift[1] .is_wysiwyg = "true";
defparam \trk_block:sig_req_rsc_shift[1] .power_up = "low";

arriaii_lcell_comb \LessThan11~1 (
	.dataa(!\trk_block:sig_req_rsc_shift[0]~q ),
	.datab(!\trk_block:sig_req_rsc_shift[1]~q ),
	.datac(!\trk_block:sig_req_rsc_shift[2]~q ),
	.datad(!\LessThan11~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan11~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan11~1 .extended_lut = "off";
defparam \LessThan11~1 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \LessThan11~1 .shared_arith = "off";

arriaii_lcell_comb \sig_req_rsc_shift~11 (
	.dataa(!\trk_block:sig_trk_last_state.s_trk_adjust_resync~q ),
	.datab(!\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.datac(!\trk_block:sig_req_rsc_shift[7]~q ),
	.datad(!\LessThan11~1_combout ),
	.datae(!\Add18~1_sumout ),
	.dataf(!\Add16~1_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_req_rsc_shift~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_req_rsc_shift~11 .extended_lut = "off";
defparam \sig_req_rsc_shift~11 .lut_mask = 64'h0000000220202022;
defparam \sig_req_rsc_shift~11 .shared_arith = "off";

arriaii_lcell_comb \sig_req_rsc_shift~4 (
	.dataa(!\sig_dgrb_state.s_track~q ),
	.datab(!\trk_block:sig_req_rsc_shift[0]~q ),
	.datac(!\sig_req_rsc_shift~2_combout ),
	.datad(!\Add15~1_sumout ),
	.datae(!\sig_trk_state~12_combout ),
	.dataf(!\sig_req_rsc_shift~11_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_req_rsc_shift~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_req_rsc_shift~4 .extended_lut = "off";
defparam \sig_req_rsc_shift~4 .lut_mask = 64'hF3F3F3A2A2A2A2A2;
defparam \sig_req_rsc_shift~4 .shared_arith = "off";

dffeas \trk_block:sig_req_rsc_shift[0] (
	.clk(clk),
	.d(\sig_req_rsc_shift~4_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_req_rsc_shift[0]~q ),
	.prn(vcc));
defparam \trk_block:sig_req_rsc_shift[0] .is_wysiwyg = "true";
defparam \trk_block:sig_req_rsc_shift[0] .power_up = "low";

arriaii_lcell_comb \sig_trk_state~11 (
	.dataa(!\trk_block:sig_req_rsc_shift[7]~q ),
	.datab(!\trk_block:sig_req_rsc_shift[0]~q ),
	.datac(!\trk_block:sig_req_rsc_shift[1]~q ),
	.datad(!\trk_block:sig_req_rsc_shift[2]~q ),
	.datae(!\LessThan11~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_trk_state~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_trk_state~11 .extended_lut = "off";
defparam \sig_trk_state~11 .lut_mask = 64'h0000100000001000;
defparam \sig_trk_state~11 .shared_arith = "off";

arriaii_lcell_comb \sig_trk_state~13 (
	.dataa(!\sig_dgrb_state.s_track~q ),
	.datab(!\trk_block:sig_trk_last_state.s_trk_adjust_resync~q ),
	.datac(!\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.datad(!\sig_trk_state~11_combout ),
	.datae(!\sig_phs_shft_end~q ),
	.dataf(!\sig_trk_state~12_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_trk_state~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_trk_state~13 .extended_lut = "off";
defparam \sig_trk_state~13 .lut_mask = 64'h0501000055515050;
defparam \sig_trk_state~13 .shared_arith = "off";

dffeas \trk_block:sig_trk_state.s_trk_adjust_resync (
	.clk(clk),
	.d(\sig_trk_state~13_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.prn(vcc));
defparam \trk_block:sig_trk_state.s_trk_adjust_resync .is_wysiwyg = "true";
defparam \trk_block:sig_trk_state.s_trk_adjust_resync .power_up = "low";

arriaii_lcell_comb \sig_trk_pll_inc_dec_n~1 (
	.dataa(!\sig_dgrb_state.s_track~q ),
	.datab(!\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_trk_pll_inc_dec_n~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_trk_pll_inc_dec_n~1 .extended_lut = "off";
defparam \sig_trk_pll_inc_dec_n~1 .lut_mask = 64'h1111111111111111;
defparam \sig_trk_pll_inc_dec_n~1 .shared_arith = "off";

dffeas \trk_block:sig_trk_last_state.s_trk_adjust_resync (
	.clk(clk),
	.d(\sig_trk_pll_inc_dec_n~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_trk_last_state.s_trk_adjust_resync~q ),
	.prn(vcc));
defparam \trk_block:sig_trk_last_state.s_trk_adjust_resync .is_wysiwyg = "true";
defparam \trk_block:sig_trk_last_state.s_trk_adjust_resync .power_up = "low";

arriaii_lcell_comb \sig_trk_state~17 (
	.dataa(!\sig_dgrb_state.s_track~q ),
	.datab(!\trk_block:sig_trk_last_state.s_trk_adjust_resync~q ),
	.datac(!\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.datad(!\sig_trk_state~11_combout ),
	.datae(!\sig_phs_shft_end~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_trk_state~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_trk_state~17 .extended_lut = "off";
defparam \sig_trk_state~17 .lut_mask = 64'h5551505055515050;
defparam \sig_trk_state~17 .shared_arith = "off";

arriaii_lcell_comb \sig_trk_state~18 (
	.dataa(!\sig_trk_state~12_combout ),
	.datab(!\sig_trk_state~17_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_trk_state~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_trk_state~18 .extended_lut = "off";
defparam \sig_trk_state~18 .lut_mask = 64'h2222222222222222;
defparam \sig_trk_state~18 .shared_arith = "off";

arriaii_lcell_comb \sig_trk_state~26 (
	.dataa(!\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.datab(!\Equal17~1_combout ),
	.datac(!\trk_block:sig_trk_state.s_trk_cdvw_calc~q ),
	.datad(!\sig_trk_state~16_combout ),
	.datae(!\sig_trk_state~18_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_trk_state~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_trk_state~26 .extended_lut = "off";
defparam \sig_trk_state~26 .lut_mask = 64'h0000110F0000110F;
defparam \sig_trk_state~26 .shared_arith = "off";

dffeas \trk_block:sig_trk_state.s_trk_cdvw_calc (
	.clk(clk),
	.d(\sig_trk_state~26_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_trk_state.s_trk_cdvw_calc~q ),
	.prn(vcc));
defparam \trk_block:sig_trk_state.s_trk_cdvw_calc .is_wysiwyg = "true";
defparam \trk_block:sig_trk_state.s_trk_cdvw_calc .power_up = "low";

arriaii_lcell_comb \sig_trk_last_state~1 (
	.dataa(!\sig_dgrb_state.s_track~q ),
	.datab(!\trk_block:sig_trk_state.s_trk_cdvw_calc~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_trk_last_state~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_trk_last_state~1 .extended_lut = "off";
defparam \sig_trk_last_state~1 .lut_mask = 64'h1111111111111111;
defparam \sig_trk_last_state~1 .shared_arith = "off";

dffeas \trk_block:sig_trk_last_state.s_trk_cdvw_calc (
	.clk(clk),
	.d(\sig_trk_last_state~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_trk_last_state.s_trk_cdvw_calc~q ),
	.prn(vcc));
defparam \trk_block:sig_trk_last_state.s_trk_cdvw_calc .is_wysiwyg = "true";
defparam \trk_block:sig_trk_last_state.s_trk_cdvw_calc .power_up = "low";

arriaii_lcell_comb \sig_trk_state~24 (
	.dataa(!\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.datab(!\sig_cdvw_state.status.calculating~q ),
	.datac(!\trk_block:sig_trk_last_state.s_trk_cdvw_calc~q ),
	.datad(!\trk_block:sig_trk_state.s_trk_cdvw_calc~q ),
	.datae(!\sig_trk_state~18_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_trk_state~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_trk_state~24 .extended_lut = "off";
defparam \sig_trk_state~24 .lut_mask = 64'h0000111F0000111F;
defparam \sig_trk_state~24 .shared_arith = "off";

dffeas \trk_block:sig_trk_state.s_trk_cdvw_wait (
	.clk(clk),
	.d(\sig_trk_state~24_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.prn(vcc));
defparam \trk_block:sig_trk_state.s_trk_cdvw_wait .is_wysiwyg = "true";
defparam \trk_block:sig_trk_state.s_trk_cdvw_wait .power_up = "low";

arriaii_lcell_comb \Add11~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add11~22 ),
	.sharein(\Add11~23 ),
	.combout(),
	.sumout(\Add11~25_sumout ),
	.cout(),
	.shareout());
defparam \Add11~25 .extended_lut = "off";
defparam \Add11~25 .lut_mask = 64'h000000000000FFFF;
defparam \Add11~25 .shared_arith = "on";

arriaii_lcell_comb \sig_mimic_delta~0 (
	.dataa(!\sig_dgrb_state.s_track~q ),
	.datab(!\sig_cdvw_state.status.valid_result~q ),
	.datac(!\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.datad(!\trk_block:sig_mimic_cdv_found~q ),
	.datae(!\Add11~25_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_mimic_delta~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_mimic_delta~0 .extended_lut = "off";
defparam \sig_mimic_delta~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \sig_mimic_delta~0 .shared_arith = "off";

dffeas \trk_block:sig_mimic_delta[6] (
	.clk(clk),
	.d(\sig_mimic_delta~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_mimic_delta~1_combout ),
	.q(\trk_block:sig_mimic_delta[6]~q ),
	.prn(vcc));
defparam \trk_block:sig_mimic_delta[6] .is_wysiwyg = "true";
defparam \trk_block:sig_mimic_delta[6] .power_up = "low";

arriaii_lcell_comb \Add15~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_mimic_delta[6]~q ),
	.datae(gnd),
	.dataf(!\trk_block:sig_req_rsc_shift[7]~q ),
	.datag(gnd),
	.cin(\Add15~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add15~29_sumout ),
	.cout(),
	.shareout());
defparam \Add15~29 .extended_lut = "off";
defparam \Add15~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add15~29 .shared_arith = "off";

arriaii_lcell_comb \sig_req_rsc_shift~1 (
	.dataa(!\trk_block:sig_mimic_delta[6]~q ),
	.datab(!\Add15~21_sumout ),
	.datac(!\Add15~25_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_req_rsc_shift~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_req_rsc_shift~1 .extended_lut = "off";
defparam \sig_req_rsc_shift~1 .lut_mask = 64'h4242424242424242;
defparam \sig_req_rsc_shift~1 .shared_arith = "off";

arriaii_lcell_comb \Add16~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_req_rsc_shift[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add16~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add16~29_sumout ),
	.cout(),
	.shareout());
defparam \Add16~29 .extended_lut = "off";
defparam \Add16~29 .lut_mask = 64'h0000FFFF0000FF00;
defparam \Add16~29 .shared_arith = "off";

arriaii_lcell_comb \Add18~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_req_rsc_shift[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add18~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add18~29_sumout ),
	.cout(),
	.shareout());
defparam \Add18~29 .extended_lut = "off";
defparam \Add18~29 .lut_mask = 64'h000000000000FF00;
defparam \Add18~29 .shared_arith = "off";

arriaii_lcell_comb \sig_req_rsc_shift~16 (
	.dataa(!\sig_trk_pll_inc_dec_n~1_combout ),
	.datab(!\trk_block:sig_trk_last_state.s_trk_adjust_resync~q ),
	.datac(!\LessThan11~1_combout ),
	.datad(!\Add16~29_sumout ),
	.datae(!\trk_block:sig_req_rsc_shift[7]~q ),
	.dataf(!\Add18~29_sumout ),
	.datag(!\sig_req_rsc_shift~2_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_req_rsc_shift~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_req_rsc_shift~16 .extended_lut = "on";
defparam \sig_req_rsc_shift~16 .lut_mask = 64'h0F4F00000F4F0404;
defparam \sig_req_rsc_shift~16 .shared_arith = "off";

arriaii_lcell_comb \sig_req_rsc_shift~3 (
	.dataa(!\sig_dgrb_state.s_track~q ),
	.datab(!\Add15~29_sumout ),
	.datac(!\sig_req_rsc_shift~1_combout ),
	.datad(!\trk_block:sig_large_drift_seen~q ),
	.datae(!\sig_trk_state~12_combout ),
	.dataf(!\sig_req_rsc_shift~16_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_req_rsc_shift~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_req_rsc_shift~3 .extended_lut = "off";
defparam \sig_req_rsc_shift~3 .lut_mask = 64'hFFFFEEEB00000000;
defparam \sig_req_rsc_shift~3 .shared_arith = "off";

dffeas \trk_block:sig_req_rsc_shift[7] (
	.clk(clk),
	.d(\sig_req_rsc_shift~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_req_rsc_shift[7]~q ),
	.prn(vcc));
defparam \trk_block:sig_req_rsc_shift[7] .is_wysiwyg = "true";
defparam \trk_block:sig_req_rsc_shift[7] .power_up = "low";

arriaii_lcell_comb \Add17~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_rsc_drift[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~2_sumout ),
	.cout(\Add17~3 ),
	.shareout());
defparam \Add17~2 .extended_lut = "off";
defparam \Add17~2 .lut_mask = 64'h000000000000FF00;
defparam \Add17~2 .shared_arith = "off";

arriaii_lcell_comb \sig_rsc_drift~0 (
	.dataa(!\trk_block:sig_trk_last_state.s_trk_adjust_resync~q ),
	.datab(!\sig_trk_pll_inc_dec_n~1_combout ),
	.datac(!\sig_trk_state~11_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_rsc_drift~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_rsc_drift~0 .extended_lut = "off";
defparam \sig_rsc_drift~0 .lut_mask = 64'h2020202020202020;
defparam \sig_rsc_drift~0 .shared_arith = "off";

arriaii_lcell_comb \sig_rsc_drift~1 (
	.dataa(!\sig_dgrb_state.s_track~q ),
	.datab(!\trk_block:sig_trk_last_state.s_trk_adjust_resync~q ),
	.datac(!\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.datad(!\sig_trk_state~11_combout ),
	.datae(!sig_addr_cmd0cke0),
	.dataf(!\trk_block:sig_mimic_cdv_found~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_rsc_drift~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_rsc_drift~1 .extended_lut = "off";
defparam \sig_rsc_drift~1 .lut_mask = 64'h00000000ABAFFBFF;
defparam \sig_rsc_drift~1 .shared_arith = "off";

arriaii_lcell_comb \sig_rsc_drift~7 (
	.dataa(!\trk_block:sig_rsc_drift[0]~q ),
	.datab(!\Add17~2_sumout ),
	.datac(!\sig_rsc_drift~0_combout ),
	.datad(!\sig_rsc_drift~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_rsc_drift~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_rsc_drift~7 .extended_lut = "off";
defparam \sig_rsc_drift~7 .lut_mask = 64'hFC54FC54FC54FC54;
defparam \sig_rsc_drift~7 .shared_arith = "off";

dffeas \trk_block:sig_rsc_drift[0] (
	.clk(clk),
	.d(\sig_rsc_drift~7_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_rsc_drift[0]~q ),
	.prn(vcc));
defparam \trk_block:sig_rsc_drift[0] .is_wysiwyg = "true";
defparam \trk_block:sig_rsc_drift[0] .power_up = "low";

arriaii_lcell_comb \Add17~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_rsc_drift[1]~q ),
	.datae(gnd),
	.dataf(!\trk_block:sig_req_rsc_shift[7]~q ),
	.datag(gnd),
	.cin(\Add17~3 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~6_sumout ),
	.cout(\Add17~7 ),
	.shareout());
defparam \Add17~6 .extended_lut = "off";
defparam \Add17~6 .lut_mask = 64'h0000FF00000000FF;
defparam \Add17~6 .shared_arith = "off";

arriaii_lcell_comb \sig_rsc_drift~6 (
	.dataa(!\trk_block:sig_rsc_drift[1]~q ),
	.datab(!\Add17~6_sumout ),
	.datac(!\sig_rsc_drift~0_combout ),
	.datad(!\sig_rsc_drift~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_rsc_drift~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_rsc_drift~6 .extended_lut = "off";
defparam \sig_rsc_drift~6 .lut_mask = 64'h0357035703570357;
defparam \sig_rsc_drift~6 .shared_arith = "off";

dffeas \trk_block:sig_rsc_drift[1] (
	.clk(clk),
	.d(\sig_rsc_drift~6_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_rsc_drift[1]~q ),
	.prn(vcc));
defparam \trk_block:sig_rsc_drift[1] .is_wysiwyg = "true";
defparam \trk_block:sig_rsc_drift[1] .power_up = "low";

arriaii_lcell_comb \Selector75~0 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_seek_cdvw~q ),
	.datab(!\sig_cdvw_state.largest_window_centre[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector75~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector75~0 .extended_lut = "off";
defparam \Selector75~0 .lut_mask = 64'h1111111111111111;
defparam \Selector75~0 .shared_arith = "off";

arriaii_lcell_comb \Selector55~0 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_idle~q ),
	.datab(!\sig_rsc_req.s_rsc_reset_cdvw~q ),
	.datac(!\rsc_block:sig_rsc_last_state.s_rsc_idle~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector55~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector55~0 .extended_lut = "off";
defparam \Selector55~0 .lut_mask = 64'h2020202020202020;
defparam \Selector55~0 .shared_arith = "off";

dffeas \rsc_block:sig_rsc_state.s_rsc_reset_cdvw (
	.clk(clk),
	.d(\Selector55~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rsc_state.s_rsc_reset_cdvw~q ),
	.prn(vcc));
defparam \rsc_block:sig_rsc_state.s_rsc_reset_cdvw .is_wysiwyg = "true";
defparam \rsc_block:sig_rsc_state.s_rsc_reset_cdvw .power_up = "low";

arriaii_lcell_comb \Selector71~3 (
	.dataa(!\rsc_block:sig_count[0]~q ),
	.datab(!\rsc_block:sig_count[1]~q ),
	.datac(!\rsc_block:sig_count[2]~q ),
	.datad(!\rsc_block:sig_count[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector71~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector71~3 .extended_lut = "off";
defparam \Selector71~3 .lut_mask = 64'h8000800080008000;
defparam \Selector71~3 .shared_arith = "off";

arriaii_lcell_comb \Selector71~2 (
	.dataa(!\rsc_block:sig_rsc_last_state.s_rsc_seek_cdvw~q ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_seek_cdvw~q ),
	.datac(!\sig_cdvw_state.status.valid_result~q ),
	.datad(!\rsc_block:sig_rsc_state.s_rsc_reset_cdvw~q ),
	.datae(!\Equal14~0_combout ),
	.dataf(!\Selector71~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector71~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector71~2 .extended_lut = "off";
defparam \Selector71~2 .lut_mask = 64'h00CC00CC00CC01CD;
defparam \Selector71~2 .shared_arith = "off";

dffeas \cal_codvw_phase[1] (
	.clk(clk),
	.d(\Selector75~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector71~2_combout ),
	.q(\cal_codvw_phase[1]~q ),
	.prn(vcc));
defparam \cal_codvw_phase[1] .is_wysiwyg = "true";
defparam \cal_codvw_phase[1] .power_up = "low";

arriaii_lcell_comb \Selector76~0 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_seek_cdvw~q ),
	.datab(!\sig_cdvw_state.largest_window_centre[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector76~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector76~0 .extended_lut = "off";
defparam \Selector76~0 .lut_mask = 64'h1111111111111111;
defparam \Selector76~0 .shared_arith = "off";

dffeas \cal_codvw_phase[0] (
	.clk(clk),
	.d(\Selector76~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector71~2_combout ),
	.q(\cal_codvw_phase[0]~q ),
	.prn(vcc));
defparam \cal_codvw_phase[0] .is_wysiwyg = "true";
defparam \cal_codvw_phase[0] .power_up = "low";

arriaii_lcell_comb \Add9~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_rsc_drift[0]~q ),
	.datae(gnd),
	.dataf(!\cal_codvw_phase[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~1_sumout ),
	.cout(\Add9~2 ),
	.shareout());
defparam \Add9~1 .extended_lut = "off";
defparam \Add9~1 .lut_mask = 64'h0000FF000000FF00;
defparam \Add9~1 .shared_arith = "off";

arriaii_lcell_comb \Add9~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_rsc_drift[1]~q ),
	.datae(gnd),
	.dataf(!\cal_codvw_phase[1]~q ),
	.datag(gnd),
	.cin(\Add9~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~5_sumout ),
	.cout(\Add9~6 ),
	.shareout());
defparam \Add9~5 .extended_lut = "off";
defparam \Add9~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add9~5 .shared_arith = "off";

arriaii_lcell_comb \Add17~10 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_rsc_drift[2]~q ),
	.datae(gnd),
	.dataf(!\trk_block:sig_req_rsc_shift[7]~q ),
	.datag(gnd),
	.cin(\Add17~7 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~10_sumout ),
	.cout(\Add17~11 ),
	.shareout());
defparam \Add17~10 .extended_lut = "off";
defparam \Add17~10 .lut_mask = 64'h0000FF00000000FF;
defparam \Add17~10 .shared_arith = "off";

arriaii_lcell_comb \sig_rsc_drift~5 (
	.dataa(!\trk_block:sig_rsc_drift[2]~q ),
	.datab(!\Add17~10_sumout ),
	.datac(!\sig_rsc_drift~0_combout ),
	.datad(!\sig_rsc_drift~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_rsc_drift~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_rsc_drift~5 .extended_lut = "off";
defparam \sig_rsc_drift~5 .lut_mask = 64'h0357035703570357;
defparam \sig_rsc_drift~5 .shared_arith = "off";

dffeas \trk_block:sig_rsc_drift[2] (
	.clk(clk),
	.d(\sig_rsc_drift~5_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_rsc_drift[2]~q ),
	.prn(vcc));
defparam \trk_block:sig_rsc_drift[2] .is_wysiwyg = "true";
defparam \trk_block:sig_rsc_drift[2] .power_up = "low";

arriaii_lcell_comb \Add17~14 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_rsc_drift[3]~q ),
	.datae(gnd),
	.dataf(!\trk_block:sig_req_rsc_shift[7]~q ),
	.datag(gnd),
	.cin(\Add17~11 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~14_sumout ),
	.cout(\Add17~15 ),
	.shareout());
defparam \Add17~14 .extended_lut = "off";
defparam \Add17~14 .lut_mask = 64'h0000FF00000000FF;
defparam \Add17~14 .shared_arith = "off";

arriaii_lcell_comb \sig_rsc_drift~4 (
	.dataa(!\trk_block:sig_rsc_drift[3]~q ),
	.datab(!\Add17~14_sumout ),
	.datac(!\sig_rsc_drift~0_combout ),
	.datad(!\sig_rsc_drift~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_rsc_drift~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_rsc_drift~4 .extended_lut = "off";
defparam \sig_rsc_drift~4 .lut_mask = 64'h0357035703570357;
defparam \sig_rsc_drift~4 .shared_arith = "off";

dffeas \trk_block:sig_rsc_drift[3] (
	.clk(clk),
	.d(\sig_rsc_drift~4_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_rsc_drift[3]~q ),
	.prn(vcc));
defparam \trk_block:sig_rsc_drift[3] .is_wysiwyg = "true";
defparam \trk_block:sig_rsc_drift[3] .power_up = "low";

arriaii_lcell_comb \Add17~18 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_rsc_drift[4]~q ),
	.datae(gnd),
	.dataf(!\trk_block:sig_req_rsc_shift[7]~q ),
	.datag(gnd),
	.cin(\Add17~15 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~18_sumout ),
	.cout(\Add17~19 ),
	.shareout());
defparam \Add17~18 .extended_lut = "off";
defparam \Add17~18 .lut_mask = 64'h0000FF00000000FF;
defparam \Add17~18 .shared_arith = "off";

arriaii_lcell_comb \sig_rsc_drift~3 (
	.dataa(!\trk_block:sig_rsc_drift[4]~q ),
	.datab(!\Add17~18_sumout ),
	.datac(!\sig_rsc_drift~0_combout ),
	.datad(!\sig_rsc_drift~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_rsc_drift~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_rsc_drift~3 .extended_lut = "off";
defparam \sig_rsc_drift~3 .lut_mask = 64'h0357035703570357;
defparam \sig_rsc_drift~3 .shared_arith = "off";

dffeas \trk_block:sig_rsc_drift[4] (
	.clk(clk),
	.d(\sig_rsc_drift~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_rsc_drift[4]~q ),
	.prn(vcc));
defparam \trk_block:sig_rsc_drift[4] .is_wysiwyg = "true";
defparam \trk_block:sig_rsc_drift[4] .power_up = "low";

arriaii_lcell_comb \Add17~22 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_rsc_drift[5]~q ),
	.datae(gnd),
	.dataf(!\trk_block:sig_req_rsc_shift[7]~q ),
	.datag(gnd),
	.cin(\Add17~19 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~22_sumout ),
	.cout(\Add17~23 ),
	.shareout());
defparam \Add17~22 .extended_lut = "off";
defparam \Add17~22 .lut_mask = 64'h0000FF00000000FF;
defparam \Add17~22 .shared_arith = "off";

arriaii_lcell_comb \sig_rsc_drift~8 (
	.dataa(!\trk_block:sig_rsc_drift[5]~q ),
	.datab(!\Add17~22_sumout ),
	.datac(!\sig_rsc_drift~0_combout ),
	.datad(!\sig_rsc_drift~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_rsc_drift~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_rsc_drift~8 .extended_lut = "off";
defparam \sig_rsc_drift~8 .lut_mask = 64'h0357035703570357;
defparam \sig_rsc_drift~8 .shared_arith = "off";

dffeas \trk_block:sig_rsc_drift[5] (
	.clk(clk),
	.d(\sig_rsc_drift~8_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_rsc_drift[5]~q ),
	.prn(vcc));
defparam \trk_block:sig_rsc_drift[5] .is_wysiwyg = "true";
defparam \trk_block:sig_rsc_drift[5] .power_up = "low";

arriaii_lcell_comb \Add17~26 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_rsc_drift[6]~q ),
	.datae(gnd),
	.dataf(!\trk_block:sig_req_rsc_shift[7]~q ),
	.datag(gnd),
	.cin(\Add17~23 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~26_sumout ),
	.cout(\Add17~27 ),
	.shareout());
defparam \Add17~26 .extended_lut = "off";
defparam \Add17~26 .lut_mask = 64'h0000FF00000000FF;
defparam \Add17~26 .shared_arith = "off";

arriaii_lcell_comb \sig_rsc_drift~9 (
	.dataa(!\trk_block:sig_rsc_drift[6]~q ),
	.datab(!\Add17~26_sumout ),
	.datac(!\sig_rsc_drift~0_combout ),
	.datad(!\sig_rsc_drift~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_rsc_drift~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_rsc_drift~9 .extended_lut = "off";
defparam \sig_rsc_drift~9 .lut_mask = 64'h0357035703570357;
defparam \sig_rsc_drift~9 .shared_arith = "off";

dffeas \trk_block:sig_rsc_drift[6] (
	.clk(clk),
	.d(\sig_rsc_drift~9_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_rsc_drift[6]~q ),
	.prn(vcc));
defparam \trk_block:sig_rsc_drift[6] .is_wysiwyg = "true";
defparam \trk_block:sig_rsc_drift[6] .power_up = "low";

arriaii_lcell_comb \Add17~30 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_rsc_drift[7]~q ),
	.datae(gnd),
	.dataf(!\trk_block:sig_req_rsc_shift[7]~q ),
	.datag(gnd),
	.cin(\Add17~27 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~30_sumout ),
	.cout(),
	.shareout());
defparam \Add17~30 .extended_lut = "off";
defparam \Add17~30 .lut_mask = 64'h0000FF000000FF00;
defparam \Add17~30 .shared_arith = "off";

arriaii_lcell_comb \sig_rsc_drift~2 (
	.dataa(!\trk_block:sig_rsc_drift[7]~q ),
	.datab(!\Add17~30_sumout ),
	.datac(!\sig_rsc_drift~0_combout ),
	.datad(!\sig_rsc_drift~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_rsc_drift~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_rsc_drift~2 .extended_lut = "off";
defparam \sig_rsc_drift~2 .lut_mask = 64'hFC54FC54FC54FC54;
defparam \sig_rsc_drift~2 .shared_arith = "off";

dffeas \trk_block:sig_rsc_drift[7] (
	.clk(clk),
	.d(\sig_rsc_drift~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_rsc_drift[7]~q ),
	.prn(vcc));
defparam \trk_block:sig_rsc_drift[7] .is_wysiwyg = "true";
defparam \trk_block:sig_rsc_drift[7] .power_up = "low";

arriaii_lcell_comb \Selector71~1 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_seek_cdvw~q ),
	.datab(!\sig_cdvw_state.largest_window_centre[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector71~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector71~1 .extended_lut = "off";
defparam \Selector71~1 .lut_mask = 64'h1111111111111111;
defparam \Selector71~1 .shared_arith = "off";

dffeas \cal_codvw_phase[5] (
	.clk(clk),
	.d(\Selector71~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector71~2_combout ),
	.q(\cal_codvw_phase[5]~q ),
	.prn(vcc));
defparam \cal_codvw_phase[5] .is_wysiwyg = "true";
defparam \cal_codvw_phase[5] .power_up = "low";

arriaii_lcell_comb \Selector72~0 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_seek_cdvw~q ),
	.datab(!\sig_cdvw_state.largest_window_centre[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector72~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector72~0 .extended_lut = "off";
defparam \Selector72~0 .lut_mask = 64'h1111111111111111;
defparam \Selector72~0 .shared_arith = "off";

dffeas \cal_codvw_phase[4] (
	.clk(clk),
	.d(\Selector72~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector71~2_combout ),
	.q(\cal_codvw_phase[4]~q ),
	.prn(vcc));
defparam \cal_codvw_phase[4] .is_wysiwyg = "true";
defparam \cal_codvw_phase[4] .power_up = "low";

arriaii_lcell_comb \Selector73~0 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_seek_cdvw~q ),
	.datab(!\sig_cdvw_state.largest_window_centre[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector73~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector73~0 .extended_lut = "off";
defparam \Selector73~0 .lut_mask = 64'h1111111111111111;
defparam \Selector73~0 .shared_arith = "off";

dffeas \cal_codvw_phase[3] (
	.clk(clk),
	.d(\Selector73~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector71~2_combout ),
	.q(\cal_codvw_phase[3]~q ),
	.prn(vcc));
defparam \cal_codvw_phase[3] .is_wysiwyg = "true";
defparam \cal_codvw_phase[3] .power_up = "low";

arriaii_lcell_comb \Selector74~0 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_seek_cdvw~q ),
	.datab(!\sig_cdvw_state.largest_window_centre[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector74~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector74~0 .extended_lut = "off";
defparam \Selector74~0 .lut_mask = 64'h1111111111111111;
defparam \Selector74~0 .shared_arith = "off";

dffeas \cal_codvw_phase[2] (
	.clk(clk),
	.d(\Selector74~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector71~2_combout ),
	.q(\cal_codvw_phase[2]~q ),
	.prn(vcc));
defparam \cal_codvw_phase[2] .is_wysiwyg = "true";
defparam \cal_codvw_phase[2] .power_up = "low";

arriaii_lcell_comb \Add9~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_rsc_drift[2]~q ),
	.datae(gnd),
	.dataf(!\cal_codvw_phase[2]~q ),
	.datag(gnd),
	.cin(\Add9~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~9_sumout ),
	.cout(\Add9~10 ),
	.shareout());
defparam \Add9~9 .extended_lut = "off";
defparam \Add9~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add9~9 .shared_arith = "off";

arriaii_lcell_comb \Add9~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_rsc_drift[3]~q ),
	.datae(gnd),
	.dataf(!\cal_codvw_phase[3]~q ),
	.datag(gnd),
	.cin(\Add9~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~13_sumout ),
	.cout(\Add9~14 ),
	.shareout());
defparam \Add9~13 .extended_lut = "off";
defparam \Add9~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add9~13 .shared_arith = "off";

arriaii_lcell_comb \Add9~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_rsc_drift[4]~q ),
	.datae(gnd),
	.dataf(!\cal_codvw_phase[4]~q ),
	.datag(gnd),
	.cin(\Add9~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~17_sumout ),
	.cout(\Add9~18 ),
	.shareout());
defparam \Add9~17 .extended_lut = "off";
defparam \Add9~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add9~17 .shared_arith = "off";

arriaii_lcell_comb \Add9~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_rsc_drift[5]~q ),
	.datae(gnd),
	.dataf(!\cal_codvw_phase[5]~q ),
	.datag(gnd),
	.cin(\Add9~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~21_sumout ),
	.cout(\Add9~22 ),
	.shareout());
defparam \Add9~21 .extended_lut = "off";
defparam \Add9~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add9~21 .shared_arith = "off";

arriaii_lcell_comb \Add9~26 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_rsc_drift[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add9~26_cout ),
	.shareout());
defparam \Add9~26 .extended_lut = "off";
defparam \Add9~26 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add9~26 .shared_arith = "off";

arriaii_lcell_comb \Add9~30 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_rsc_drift[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~26_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add9~30_cout ),
	.shareout());
defparam \Add9~30 .extended_lut = "off";
defparam \Add9~30 .lut_mask = 64'h0000FFFF0000FF00;
defparam \Add9~30 .shared_arith = "off";

arriaii_lcell_comb \Add9~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_rsc_drift[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add9~30_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add9~33_sumout ),
	.cout(),
	.shareout());
defparam \Add9~33 .extended_lut = "off";
defparam \Add9~33 .lut_mask = 64'h0000FFFF0000FF00;
defparam \Add9~33 .shared_arith = "off";

arriaii_lcell_comb \rsc_block:sig_num_phase_shifts[2]~0 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_reset_cdvw~q ),
	.datab(!\Add9~33_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rsc_block:sig_num_phase_shifts[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rsc_block:sig_num_phase_shifts[2]~0 .extended_lut = "off";
defparam \rsc_block:sig_num_phase_shifts[2]~0 .lut_mask = 64'h4444444444444444;
defparam \rsc_block:sig_num_phase_shifts[2]~0 .shared_arith = "off";

dffeas sig_phs_shft_busy(
	.clk(clk),
	.d(\phs_shft_busy_reg:phs_shft_busy_2r~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_phs_shft_busy~q ),
	.prn(vcc));
defparam sig_phs_shft_busy.is_wysiwyg = "true";
defparam sig_phs_shft_busy.power_up = "low";

arriaii_lcell_comb \Selector50~0 (
	.dataa(!\Equal13~0_combout ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_next_phase~q ),
	.datac(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datad(!\rsc_block:sig_chkd_all_dq_pins~q ),
	.datae(!\Selector53~0_combout ),
	.dataf(!\sig_phs_shft_end~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector50~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector50~0 .extended_lut = "off";
defparam \Selector50~0 .lut_mask = 64'h3333333700000005;
defparam \Selector50~0 .shared_arith = "off";

dffeas \rsc_block:sig_rsc_state.s_rsc_next_phase (
	.clk(clk),
	.d(\Selector50~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rsc_state.s_rsc_next_phase~q ),
	.prn(vcc));
defparam \rsc_block:sig_rsc_state.s_rsc_next_phase .is_wysiwyg = "true";
defparam \rsc_block:sig_rsc_state.s_rsc_next_phase .power_up = "low";

arriaii_lcell_comb \WideOr17~0 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_rewind_phase~q ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_next_phase~q ),
	.datac(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datad(!\rsc_block:sig_rsc_state.s_rsc_reset_cdvw~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr17~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr17~0 .extended_lut = "off";
defparam \WideOr17~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \WideOr17~0 .shared_arith = "off";

arriaii_lcell_comb \Selector56~0 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_rewind_phase~q ),
	.datab(!\Equal13~0_combout ),
	.datac(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datad(!\rsc_block:sig_rsc_state.s_rsc_reset_cdvw~q ),
	.datae(!\rsc_block:sig_chkd_all_dq_pins~q ),
	.dataf(!\Selector53~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector56~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector56~0 .extended_lut = "off";
defparam \Selector56~0 .lut_mask = 64'h11FF11FF11FF1DFF;
defparam \Selector56~0 .shared_arith = "off";

dffeas \rsc_block:sig_rsc_state.s_rsc_rewind_phase (
	.clk(clk),
	.d(\Selector56~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rsc_state.s_rsc_rewind_phase~q ),
	.prn(vcc));
defparam \rsc_block:sig_rsc_state.s_rsc_rewind_phase .is_wysiwyg = "true";
defparam \rsc_block:sig_rsc_state.s_rsc_rewind_phase .power_up = "low";

arriaii_lcell_comb \rsc_block:sig_num_phase_shifts[2]~3 (
	.dataa(!\sig_phs_shft_busy_1t~q ),
	.datab(!\sig_phs_shft_busy~q ),
	.datac(!\sig_phs_shft_end~q ),
	.datad(!\WideOr17~0_combout ),
	.datae(!\rsc_block:sig_rsc_state.s_rsc_next_phase~q ),
	.dataf(!\rsc_block:sig_rsc_state.s_rsc_rewind_phase~q ),
	.datag(!\Equal13~0_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rsc_block:sig_num_phase_shifts[2]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rsc_block:sig_num_phase_shifts[2]~3 .extended_lut = "on";
defparam \rsc_block:sig_num_phase_shifts[2]~3 .lut_mask = 64'hFF00FFF0FF0BFFBB;
defparam \rsc_block:sig_num_phase_shifts[2]~3 .shared_arith = "off";

arriaii_lcell_comb \rsc_block:sig_num_phase_shifts[2]~1 (
	.dataa(!\Equal13~0_combout ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datac(!\rsc_block:sig_chkd_all_dq_pins~q ),
	.datad(!\Selector53~0_combout ),
	.datae(!\rsc_block:sig_num_phase_shifts[2]~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rsc_block:sig_num_phase_shifts[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rsc_block:sig_num_phase_shifts[2]~1 .extended_lut = "off";
defparam \rsc_block:sig_num_phase_shifts[2]~1 .lut_mask = 64'hCCCE0000CCCE0000;
defparam \rsc_block:sig_num_phase_shifts[2]~1 .shared_arith = "off";

arriaii_lcell_comb \rsc_block:sig_num_phase_shifts[5]~0 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_rewind_phase~q ),
	.datab(!\Equal13~0_combout ),
	.datac(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rsc_block:sig_num_phase_shifts[5]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rsc_block:sig_num_phase_shifts[5]~0 .extended_lut = "off";
defparam \rsc_block:sig_num_phase_shifts[5]~0 .lut_mask = 64'hB0B0B0B0B0B0B0B0;
defparam \rsc_block:sig_num_phase_shifts[5]~0 .shared_arith = "off";

arriaii_lcell_comb \Add5~6 (
	.dataa(!\rsc_block:sig_num_phase_shifts[1]~q ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_reset_cdvw~q ),
	.datac(!\Add9~5_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add5~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add5~6 .extended_lut = "off";
defparam \Add5~6 .lut_mask = 64'h4747474747474747;
defparam \Add5~6 .shared_arith = "off";

arriaii_lcell_comb \Add5~1 (
	.dataa(!\rsc_block:sig_num_phase_shifts[0]~q ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_reset_cdvw~q ),
	.datac(!\Add9~1_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add5~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add5~1 .extended_lut = "off";
defparam \Add5~1 .lut_mask = 64'h4747474747474747;
defparam \Add5~1 .shared_arith = "off";

arriaii_lcell_comb \Add5~8 (
	.dataa(!\WideOr17~0_combout ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datac(!\rsc_block:sig_rsc_state.s_rsc_rewind_phase~q ),
	.datad(!\Add5~6_combout ),
	.datae(gnd),
	.dataf(!\rsc_block:sig_rsc_state.s_rsc_next_phase~q ),
	.datag(gnd),
	.cin(\Add5~4 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~8_sumout ),
	.cout(\Add5~9 ),
	.shareout());
defparam \Add5~8 .extended_lut = "off";
defparam \Add5~8 .lut_mask = 64'h0000F00000004400;
defparam \Add5~8 .shared_arith = "off";

arriaii_lcell_comb \rsc_block:sig_num_phase_shifts[1]~0 (
	.dataa(!\rsc_block:sig_num_phase_shifts[1]~q ),
	.datab(!\Add9~5_sumout ),
	.datac(!\rsc_block:sig_num_phase_shifts[2]~0_combout ),
	.datad(!\rsc_block:sig_num_phase_shifts[2]~1_combout ),
	.datae(!\rsc_block:sig_num_phase_shifts[5]~0_combout ),
	.dataf(!\Add5~8_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rsc_block:sig_num_phase_shifts[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rsc_block:sig_num_phase_shifts[1]~0 .extended_lut = "off";
defparam \rsc_block:sig_num_phase_shifts[1]~0 .lut_mask = 64'h550055FC5500550C;
defparam \rsc_block:sig_num_phase_shifts[1]~0 .shared_arith = "off";

dffeas \rsc_block:sig_num_phase_shifts[1] (
	.clk(clk),
	.d(\rsc_block:sig_num_phase_shifts[1]~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_num_phase_shifts[1]~q ),
	.prn(vcc));
defparam \rsc_block:sig_num_phase_shifts[1] .is_wysiwyg = "true";
defparam \rsc_block:sig_num_phase_shifts[1] .power_up = "low";

arriaii_lcell_comb \Add5~11 (
	.dataa(!\rsc_block:sig_num_phase_shifts[2]~q ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_reset_cdvw~q ),
	.datac(!\Add9~9_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add5~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add5~11 .extended_lut = "off";
defparam \Add5~11 .lut_mask = 64'h4747474747474747;
defparam \Add5~11 .shared_arith = "off";

arriaii_lcell_comb \Add5~13 (
	.dataa(!\WideOr17~0_combout ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_rewind_phase~q ),
	.datac(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datad(!\Add5~11_combout ),
	.datae(gnd),
	.dataf(!\rsc_block:sig_rsc_state.s_rsc_next_phase~q ),
	.datag(gnd),
	.cin(\Add5~9 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~13_sumout ),
	.cout(\Add5~14 ),
	.shareout());
defparam \Add5~13 .extended_lut = "off";
defparam \Add5~13 .lut_mask = 64'h0000CC0000005000;
defparam \Add5~13 .shared_arith = "off";

arriaii_lcell_comb \rsc_block:sig_num_phase_shifts[2]~2 (
	.dataa(!\rsc_block:sig_num_phase_shifts[2]~q ),
	.datab(!\Add9~9_sumout ),
	.datac(!\rsc_block:sig_num_phase_shifts[2]~0_combout ),
	.datad(!\rsc_block:sig_num_phase_shifts[2]~1_combout ),
	.datae(!\rsc_block:sig_num_phase_shifts[5]~0_combout ),
	.dataf(!\Add5~13_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rsc_block:sig_num_phase_shifts[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rsc_block:sig_num_phase_shifts[2]~2 .extended_lut = "off";
defparam \rsc_block:sig_num_phase_shifts[2]~2 .lut_mask = 64'h550055FC5500550C;
defparam \rsc_block:sig_num_phase_shifts[2]~2 .shared_arith = "off";

dffeas \rsc_block:sig_num_phase_shifts[2] (
	.clk(clk),
	.d(\rsc_block:sig_num_phase_shifts[2]~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_num_phase_shifts[2]~q ),
	.prn(vcc));
defparam \rsc_block:sig_num_phase_shifts[2] .is_wysiwyg = "true";
defparam \rsc_block:sig_num_phase_shifts[2] .power_up = "low";

arriaii_lcell_comb \Add5~16 (
	.dataa(!\rsc_block:sig_num_phase_shifts[3]~q ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_reset_cdvw~q ),
	.datac(!\Add9~13_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add5~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add5~16 .extended_lut = "off";
defparam \Add5~16 .lut_mask = 64'h4747474747474747;
defparam \Add5~16 .shared_arith = "off";

arriaii_lcell_comb \Add5~18 (
	.dataa(!\WideOr17~0_combout ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_rewind_phase~q ),
	.datac(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datad(!\Add5~16_combout ),
	.datae(gnd),
	.dataf(!\rsc_block:sig_rsc_state.s_rsc_next_phase~q ),
	.datag(gnd),
	.cin(\Add5~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~18_sumout ),
	.cout(\Add5~19 ),
	.shareout());
defparam \Add5~18 .extended_lut = "off";
defparam \Add5~18 .lut_mask = 64'h0000CC0000005000;
defparam \Add5~18 .shared_arith = "off";

arriaii_lcell_comb \rsc_block:sig_num_phase_shifts[3]~0 (
	.dataa(!\rsc_block:sig_num_phase_shifts[3]~q ),
	.datab(!\Add9~13_sumout ),
	.datac(!\rsc_block:sig_num_phase_shifts[2]~0_combout ),
	.datad(!\rsc_block:sig_num_phase_shifts[2]~1_combout ),
	.datae(!\rsc_block:sig_num_phase_shifts[5]~0_combout ),
	.dataf(!\Add5~18_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rsc_block:sig_num_phase_shifts[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rsc_block:sig_num_phase_shifts[3]~0 .extended_lut = "off";
defparam \rsc_block:sig_num_phase_shifts[3]~0 .lut_mask = 64'h550055FC5500550C;
defparam \rsc_block:sig_num_phase_shifts[3]~0 .shared_arith = "off";

dffeas \rsc_block:sig_num_phase_shifts[3] (
	.clk(clk),
	.d(\rsc_block:sig_num_phase_shifts[3]~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_num_phase_shifts[3]~q ),
	.prn(vcc));
defparam \rsc_block:sig_num_phase_shifts[3] .is_wysiwyg = "true";
defparam \rsc_block:sig_num_phase_shifts[3] .power_up = "low";

arriaii_lcell_comb \Add5~21 (
	.dataa(!\rsc_block:sig_num_phase_shifts[5]~q ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_reset_cdvw~q ),
	.datac(!\Add9~21_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add5~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add5~21 .extended_lut = "off";
defparam \Add5~21 .lut_mask = 64'h4747474747474747;
defparam \Add5~21 .shared_arith = "off";

arriaii_lcell_comb \Add5~22 (
	.dataa(!\rsc_block:sig_num_phase_shifts[4]~q ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_reset_cdvw~q ),
	.datac(!\Add9~17_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add5~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add5~22 .extended_lut = "off";
defparam \Add5~22 .lut_mask = 64'h4747474747474747;
defparam \Add5~22 .shared_arith = "off";

arriaii_lcell_comb \Add5~24 (
	.dataa(!\WideOr17~0_combout ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_rewind_phase~q ),
	.datac(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datad(!\Add5~22_combout ),
	.datae(gnd),
	.dataf(!\rsc_block:sig_rsc_state.s_rsc_next_phase~q ),
	.datag(gnd),
	.cin(\Add5~19 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~24_sumout ),
	.cout(\Add5~25 ),
	.shareout());
defparam \Add5~24 .extended_lut = "off";
defparam \Add5~24 .lut_mask = 64'h0000CC0000005000;
defparam \Add5~24 .shared_arith = "off";

arriaii_lcell_comb \Add5~28 (
	.dataa(!\WideOr17~0_combout ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_rewind_phase~q ),
	.datac(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datad(!\Add5~21_combout ),
	.datae(gnd),
	.dataf(!\rsc_block:sig_rsc_state.s_rsc_next_phase~q ),
	.datag(gnd),
	.cin(\Add5~25 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add5~28_sumout ),
	.cout(),
	.shareout());
defparam \Add5~28 .extended_lut = "off";
defparam \Add5~28 .lut_mask = 64'h0000CC0000005000;
defparam \Add5~28 .shared_arith = "off";

arriaii_lcell_comb \rsc_block:sig_num_phase_shifts[5]~1 (
	.dataa(!\rsc_block:sig_num_phase_shifts[5]~q ),
	.datab(!\Add9~21_sumout ),
	.datac(!\rsc_block:sig_num_phase_shifts[2]~0_combout ),
	.datad(!\rsc_block:sig_num_phase_shifts[2]~1_combout ),
	.datae(!\rsc_block:sig_num_phase_shifts[5]~0_combout ),
	.dataf(!\Add5~28_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rsc_block:sig_num_phase_shifts[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rsc_block:sig_num_phase_shifts[5]~1 .extended_lut = "off";
defparam \rsc_block:sig_num_phase_shifts[5]~1 .lut_mask = 64'h550055FC5500550C;
defparam \rsc_block:sig_num_phase_shifts[5]~1 .shared_arith = "off";

dffeas \rsc_block:sig_num_phase_shifts[5] (
	.clk(clk),
	.d(\rsc_block:sig_num_phase_shifts[5]~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_num_phase_shifts[5]~q ),
	.prn(vcc));
defparam \rsc_block:sig_num_phase_shifts[5] .is_wysiwyg = "true";
defparam \rsc_block:sig_num_phase_shifts[5] .power_up = "low";

arriaii_lcell_comb \rsc_block:sig_num_phase_shifts[4]~0 (
	.dataa(!\rsc_block:sig_num_phase_shifts[4]~q ),
	.datab(!\Add9~17_sumout ),
	.datac(!\rsc_block:sig_num_phase_shifts[2]~0_combout ),
	.datad(!\rsc_block:sig_num_phase_shifts[2]~1_combout ),
	.datae(!\rsc_block:sig_num_phase_shifts[5]~0_combout ),
	.dataf(!\Add5~24_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rsc_block:sig_num_phase_shifts[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rsc_block:sig_num_phase_shifts[4]~0 .extended_lut = "off";
defparam \rsc_block:sig_num_phase_shifts[4]~0 .lut_mask = 64'h550055FC5500550C;
defparam \rsc_block:sig_num_phase_shifts[4]~0 .shared_arith = "off";

dffeas \rsc_block:sig_num_phase_shifts[4] (
	.clk(clk),
	.d(\rsc_block:sig_num_phase_shifts[4]~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_num_phase_shifts[4]~q ),
	.prn(vcc));
defparam \rsc_block:sig_num_phase_shifts[4] .is_wysiwyg = "true";
defparam \rsc_block:sig_num_phase_shifts[4] .power_up = "low";

arriaii_lcell_comb \Equal13~0 (
	.dataa(!\rsc_block:sig_num_phase_shifts[0]~q ),
	.datab(!\rsc_block:sig_num_phase_shifts[1]~q ),
	.datac(!\rsc_block:sig_num_phase_shifts[2]~q ),
	.datad(!\rsc_block:sig_num_phase_shifts[3]~q ),
	.datae(!\rsc_block:sig_num_phase_shifts[5]~q ),
	.dataf(!\rsc_block:sig_num_phase_shifts[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal13~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal13~0 .extended_lut = "off";
defparam \Equal13~0 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \Equal13~0 .shared_arith = "off";

arriaii_lcell_comb \Selector71~0 (
	.dataa(!\rsc_block:sig_rsc_last_state.s_rsc_seek_cdvw~q ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_seek_cdvw~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector71~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector71~0 .extended_lut = "off";
defparam \Selector71~0 .lut_mask = 64'h1111111111111111;
defparam \Selector71~0 .shared_arith = "off";

arriaii_lcell_comb \Selector85~0 (
	.dataa(!\sig_dgrb_state.s_read_mtp~q ),
	.datab(!\sig_cdvw_state.status.valid_result~q ),
	.datac(!\sig_cdvw_state.status.calculating~q ),
	.datad(!\rsc_block:sig_rsc_state.s_rsc_cdvw_wait~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector85~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector85~0 .extended_lut = "off";
defparam \Selector85~0 .lut_mask = 64'h00D000D000D000D0;
defparam \Selector85~0 .shared_arith = "off";

arriaii_lcell_comb \Selector85~1 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_rewind_phase~q ),
	.datab(!\Equal13~0_combout ),
	.datac(!\Equal14~1_combout ),
	.datad(!\Selector71~0_combout ),
	.datae(!\Selector85~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector85~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector85~1 .extended_lut = "off";
defparam \Selector85~1 .lut_mask = 64'h444FFFFF444FFFFF;
defparam \Selector85~1 .shared_arith = "off";

dffeas sig_rsc_ack(
	.clk(clk),
	.d(\Selector85~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_rsc_ack~q ),
	.prn(vcc));
defparam sig_rsc_ack.is_wysiwyg = "true";
defparam sig_rsc_ack.power_up = "low";

arriaii_lcell_comb \sig_rsc_req~16 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_rsc_ack~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_rsc_req~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_rsc_req~16 .extended_lut = "off";
defparam \sig_rsc_req~16 .lut_mask = 64'h4444444444444444;
defparam \sig_rsc_req~16 .shared_arith = "off";

dffeas \sig_rsc_req.s_rsc_reset_cdvw (
	.clk(clk),
	.d(\sig_rsc_req~16_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_rsc_req.s_rsc_reset_cdvw~q ),
	.prn(vcc));
defparam \sig_rsc_req.s_rsc_reset_cdvw .is_wysiwyg = "true";
defparam \sig_rsc_req.s_rsc_reset_cdvw .power_up = "low";

arriaii_lcell_comb \sig_rsc_req~17 (
	.dataa(!\sig_dgrb_state.s_seek_cdvw~q ),
	.datab(!\sig_rsc_ack~q ),
	.datac(!\sig_dgrb_state.s_read_mtp~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_rsc_req~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_rsc_req~17 .extended_lut = "off";
defparam \sig_rsc_req~17 .lut_mask = 64'h4C4C4C4C4C4C4C4C;
defparam \sig_rsc_req~17 .shared_arith = "off";

dffeas \sig_rsc_req.s_rsc_cdvw_calc (
	.clk(clk),
	.d(\sig_rsc_req~17_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_rsc_req.s_rsc_cdvw_calc~q ),
	.prn(vcc));
defparam \sig_rsc_req.s_rsc_cdvw_calc .is_wysiwyg = "true";
defparam \sig_rsc_req.s_rsc_cdvw_calc .power_up = "low";

arriaii_lcell_comb \Selector49~0 (
	.dataa(!\Selector85~1_combout ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_idle~q ),
	.datac(!\sig_rsc_req.s_rsc_reset_cdvw~q ),
	.datad(!\rsc_block:sig_rsc_last_state.s_rsc_idle~q ),
	.datae(!\sig_rsc_req.s_rsc_cdvw_calc~q ),
	.dataf(!\sig_rsc_req.s_rsc_test_phase~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector49~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector49~0 .extended_lut = "off";
defparam \Selector49~0 .lut_mask = 64'h2A22AA22AA22AA22;
defparam \Selector49~0 .shared_arith = "off";

dffeas \rsc_block:sig_rsc_state.s_rsc_idle (
	.clk(clk),
	.d(\Selector49~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rsc_state.s_rsc_idle~q ),
	.prn(vcc));
defparam \rsc_block:sig_rsc_state.s_rsc_idle .is_wysiwyg = "true";
defparam \rsc_block:sig_rsc_state.s_rsc_idle .power_up = "low";

dffeas \rsc_block:sig_rsc_last_state.s_rsc_idle (
	.clk(clk),
	.d(\rsc_block:sig_rsc_state.s_rsc_idle~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rsc_last_state.s_rsc_idle~q ),
	.prn(vcc));
defparam \rsc_block:sig_rsc_last_state.s_rsc_idle .is_wysiwyg = "true";
defparam \rsc_block:sig_rsc_last_state.s_rsc_idle .power_up = "low";

arriaii_lcell_comb \Selector57~0 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_idle~q ),
	.datab(!\rsc_block:sig_rsc_last_state.s_rsc_idle~q ),
	.datac(!\sig_rsc_req.s_rsc_cdvw_calc~q ),
	.datad(!\sig_rsc_cdvw_calc~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector57~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector57~0 .extended_lut = "off";
defparam \Selector57~0 .lut_mask = 64'h08FF08FF08FF08FF;
defparam \Selector57~0 .shared_arith = "off";

dffeas \rsc_block:sig_rsc_state.s_rsc_cdvw_calc (
	.clk(clk),
	.d(\Selector57~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rsc_block:sig_rsc_state.s_rsc_cdvw_calc~q ),
	.prn(vcc));
defparam \rsc_block:sig_rsc_state.s_rsc_cdvw_calc .is_wysiwyg = "true";
defparam \rsc_block:sig_rsc_state.s_rsc_cdvw_calc .power_up = "low";

arriaii_lcell_comb \sig_rsc_cdvw_calc~0 (
	.dataa(!\rsc_block:sig_rsc_last_state.s_rsc_cdvw_calc~q ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_cdvw_calc~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_rsc_cdvw_calc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_rsc_cdvw_calc~0 .extended_lut = "off";
defparam \sig_rsc_cdvw_calc~0 .lut_mask = 64'h2222222222222222;
defparam \sig_rsc_cdvw_calc~0 .shared_arith = "off";

dffeas sig_rsc_cdvw_calc(
	.clk(clk),
	.d(\sig_rsc_cdvw_calc~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_rsc_cdvw_calc~q ),
	.prn(vcc));
defparam sig_rsc_cdvw_calc.is_wysiwyg = "true";
defparam sig_rsc_cdvw_calc.power_up = "low";

arriaii_lcell_comb \sig_trk_cdvw_calc~0 (
	.dataa(!\trk_block:sig_trk_last_state.s_trk_cdvw_calc~q ),
	.datab(!\trk_block:sig_trk_state.s_trk_cdvw_calc~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_trk_cdvw_calc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_trk_cdvw_calc~0 .extended_lut = "off";
defparam \sig_trk_cdvw_calc~0 .lut_mask = 64'h2222222222222222;
defparam \sig_trk_cdvw_calc~0 .shared_arith = "off";

dffeas sig_trk_cdvw_calc(
	.clk(clk),
	.d(\sig_trk_cdvw_calc~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_track~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_trk_cdvw_calc~q ),
	.prn(vcc));
defparam sig_trk_cdvw_calc.is_wysiwyg = "true";
defparam sig_trk_cdvw_calc.power_up = "low";

arriaii_lcell_comb \Selector33~0 (
	.dataa(!\sig_dgrb_state.s_seek_cdvw~q ),
	.datab(!\sig_dgrb_state.s_test_phases~q ),
	.datac(!\sig_dgrb_state.s_track~q ),
	.datad(!\sig_dgrb_state.s_read_mtp~q ),
	.datae(!\sig_rsc_cdvw_calc~q ),
	.dataf(!\sig_trk_cdvw_calc~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector33~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector33~0 .extended_lut = "off";
defparam \Selector33~0 .lut_mask = 64'h000077FF0F0F7FFF;
defparam \Selector33~0 .shared_arith = "off";

arriaii_lcell_comb \sig_cdvw_state.current_bit[5]~1 (
	.dataa(!\sig_dgrb_state.s_track~q ),
	.datab(!\sig_cdvw_state.current_bit[0]~q ),
	.datac(!\sig_cdvw_state.current_bit[5]~q ),
	.datad(!\sig_cdvw_state.current_bit[2]~q ),
	.datae(!\sig_cdvw_state.current_bit[3]~q ),
	.dataf(!\sig_cdvw_state.current_bit[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_cdvw_state.current_bit[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_cdvw_state.current_bit[5]~1 .extended_lut = "off";
defparam \sig_cdvw_state.current_bit[5]~1 .lut_mask = 64'h0505050505050517;
defparam \sig_cdvw_state.current_bit[5]~1 .shared_arith = "off";

arriaii_lcell_comb \sig_cdvw_state.current_bit[5]~2 (
	.dataa(!\sig_cdvw_state.current_bit[5]~q ),
	.datab(!\Selector33~0_combout ),
	.datac(!\sig_cdvw_state.current_bit[5]~1_combout ),
	.datad(!\cdvw_block:sig_cdvw_calc_1t~q ),
	.datae(!\sig_cdvw_state.current_bit[1]~q ),
	.dataf(!\cdvw_proc~1_combout ),
	.datag(!\sig_dgrb_state.s_track~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_cdvw_state.current_bit[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_cdvw_state.current_bit[5]~2 .extended_lut = "on";
defparam \sig_cdvw_state.current_bit[5]~2 .lut_mask = 64'h37053F0FFFFFFFFF;
defparam \sig_cdvw_state.current_bit[5]~2 .shared_arith = "off";

dffeas \sig_cdvw_state.current_bit[0] (
	.clk(clk),
	.d(\Add4~1_sumout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_bit[5]~2_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.current_bit[5]~0_combout ),
	.q(\sig_cdvw_state.current_bit[0]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_bit[0] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_bit[0] .power_up = "low";

dffeas \sig_cdvw_state.current_bit[1] (
	.clk(clk),
	.d(\Add4~5_sumout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.current_bit[5]~2_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.current_bit[5]~0_combout ),
	.q(\sig_cdvw_state.current_bit[1]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.current_bit[1] .is_wysiwyg = "true";
defparam \sig_cdvw_state.current_bit[1] .power_up = "low";

arriaii_lcell_comb \find_centre_of_largest_data_valid_window~0 (
	.dataa(!\sig_cdvw_state.current_bit[3]~q ),
	.datab(!\sig_cdvw_state.current_bit[4]~q ),
	.datac(!\sig_cdvw_state.found_a_good_edge~q ),
	.datad(!\sig_cdvw_state.current_bit[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\find_centre_of_largest_data_valid_window~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \find_centre_of_largest_data_valid_window~0 .extended_lut = "off";
defparam \find_centre_of_largest_data_valid_window~0 .lut_mask = 64'h8000800080008000;
defparam \find_centre_of_largest_data_valid_window~0 .shared_arith = "off";

arriaii_lcell_comb \find_centre_of_largest_data_valid_window~1 (
	.dataa(!\sig_cdvw_state.current_bit[0]~q ),
	.datab(!\sig_cdvw_state.current_bit[1]~q ),
	.datac(!\sig_cdvw_state.current_bit[2]~q ),
	.datad(!\find_centre_of_largest_data_valid_window~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\find_centre_of_largest_data_valid_window~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \find_centre_of_largest_data_valid_window~1 .extended_lut = "off";
defparam \find_centre_of_largest_data_valid_window~1 .lut_mask = 64'h0080008000800080;
defparam \find_centre_of_largest_data_valid_window~1 .shared_arith = "off";

arriaii_lcell_comb \v_cdvw_state~1 (
	.dataa(!\sig_cdvw_state.status.calculating~q ),
	.datab(!\v_cdvw_state~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~1 .extended_lut = "off";
defparam \v_cdvw_state~1 .lut_mask = 64'h1111111111111111;
defparam \v_cdvw_state~1 .shared_arith = "off";

dffeas \sig_cdvw_state.largest_window_size[1] (
	.clk(clk),
	.d(\sig_cdvw_state.current_window_size[1]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\v_cdvw_state~2_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.largest_window_centre[1]~0_combout ),
	.q(\sig_cdvw_state.largest_window_size[1]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.largest_window_size[1] .is_wysiwyg = "true";
defparam \sig_cdvw_state.largest_window_size[1] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~16 (
	.dataa(!\sig_cdvw_state.largest_window_size[2]~q ),
	.datab(!\sig_cdvw_state.current_window_size[2]~q ),
	.datac(!\sig_cdvw_state.largest_window_size[1]~q ),
	.datad(!\sig_cdvw_state.current_window_size[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~16 .extended_lut = "off";
defparam \v_cdvw_state~16 .lut_mask = 64'h9009900990099009;
defparam \v_cdvw_state~16 .shared_arith = "off";

arriaii_lcell_comb \v_cdvw_state~17 (
	.dataa(!\sig_cdvw_state.largest_window_size[0]~q ),
	.datab(!\sig_cdvw_state.current_window_size[0]~q ),
	.datac(!\sig_cdvw_state.largest_window_size[3]~q ),
	.datad(!\sig_cdvw_state.current_window_size[3]~q ),
	.datae(!\LessThan3~1_combout ),
	.dataf(!\v_cdvw_state~16_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~17 .extended_lut = "off";
defparam \v_cdvw_state~17 .lut_mask = 64'h0000000000009009;
defparam \v_cdvw_state~17 .shared_arith = "off";

arriaii_lcell_comb \v_cdvw_state~18 (
	.dataa(!\sig_cdvw_state.multiple_eq_windows~q ),
	.datab(!\v_cdvw_state~2_combout ),
	.datac(!\v_cdvw_state~5_combout ),
	.datad(!\LessThan3~3_combout ),
	.datae(!\v_cdvw_state~17_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~18 .extended_lut = "off";
defparam \v_cdvw_state~18 .lut_mask = 64'h4044404C4044404C;
defparam \v_cdvw_state~18 .shared_arith = "off";

dffeas \sig_cdvw_state.multiple_eq_windows (
	.clk(clk),
	.d(\v_cdvw_state~18_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_cdvw_state.multiple_eq_windows~q ),
	.prn(vcc));
defparam \sig_cdvw_state.multiple_eq_windows .is_wysiwyg = "true";
defparam \sig_cdvw_state.multiple_eq_windows .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~3 (
	.dataa(!\sig_cdvw_state.status.valid_result~q ),
	.datab(!\find_centre_of_largest_data_valid_window~1_combout ),
	.datac(!\v_cdvw_state~1_combout ),
	.datad(!\sig_cdvw_state.multiple_eq_windows~q ),
	.datae(!\v_cdvw_state~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~3 .extended_lut = "off";
defparam \v_cdvw_state~3 .lut_mask = 64'h5C5000005C500000;
defparam \v_cdvw_state~3 .shared_arith = "off";

dffeas \sig_cdvw_state.status.valid_result (
	.clk(clk),
	.d(\v_cdvw_state~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_cdvw_state.status.valid_result~q ),
	.prn(vcc));
defparam \sig_cdvw_state.status.valid_result .is_wysiwyg = "true";
defparam \sig_cdvw_state.status.valid_result .power_up = "low";

arriaii_lcell_comb \Selector128~0 (
	.dataa(!\trk_block:sig_trk_state.s_trk_complete~q ),
	.datab(!\sig_cdvw_state.status.valid_result~q ),
	.datac(!\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.datad(!\sig_cdvw_state.status.calculating~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector128~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector128~0 .extended_lut = "off";
defparam \Selector128~0 .lut_mask = 64'h5D555D555D555D55;
defparam \Selector128~0 .shared_arith = "off";

dffeas sig_trk_ack(
	.clk(clk),
	.d(\Selector128~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_track~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_trk_ack~q ),
	.prn(vcc));
defparam sig_trk_ack.is_wysiwyg = "true";
defparam sig_trk_ack.power_up = "low";

dffeas \tp_match_block:sig_rdata_valid_1t (
	.clk(clk),
	.d(rdata_valid[0]),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_valid_1t~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_valid_1t .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_valid_1t .power_up = "low";

dffeas \tp_match_block:sig_rdata_valid_2t (
	.clk(clk),
	.d(\tp_match_block:sig_rdata_valid_1t~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tp_match_block:sig_rdata_valid_2t~q ),
	.prn(vcc));
defparam \tp_match_block:sig_rdata_valid_2t .is_wysiwyg = "true";
defparam \tp_match_block:sig_rdata_valid_2t .power_up = "low";

arriaii_lcell_comb \poa_match_proc~0 (
	.dataa(!\tp_match_block:sig_rdata_valid_1t~q ),
	.datab(!\tp_match_block:sig_rdata_valid_2t~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\poa_match_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \poa_match_proc~0 .extended_lut = "off";
defparam \poa_match_proc~0 .lut_mask = 64'h2222222222222222;
defparam \poa_match_proc~0 .shared_arith = "off";

dffeas sig_poa_match_en(
	.clk(clk),
	.d(\poa_match_proc~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_poa_match_en~q ),
	.prn(vcc));
defparam sig_poa_match_en.is_wysiwyg = "true";
defparam sig_poa_match_en.power_up = "low";

arriaii_lcell_comb \Equal16~0 (
	.dataa(!\Equal15~0_combout ),
	.datab(!\tp_match_block:sig_rdata_current_pin[10]~q ),
	.datac(!\tp_match_block:sig_rdata_current_pin[11]~q ),
	.datad(!\tp_match_block:sig_rdata_current_pin[15]~q ),
	.datae(!\tp_match_block:sig_rdata_current_pin[14]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal16~0 .extended_lut = "off";
defparam \Equal16~0 .lut_mask = 64'h0000000100000001;
defparam \Equal16~0 .shared_arith = "off";

dffeas sig_poa_match(
	.clk(clk),
	.d(\Equal16~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_poa_match~q ),
	.prn(vcc));
defparam sig_poa_match.is_wysiwyg = "true";
defparam sig_poa_match.power_up = "low";

arriaii_lcell_comb \sig_poa_state~0 (
	.dataa(!\sig_dgrb_state.s_poa_cal~q ),
	.datab(!\poa_block:sig_poa_state~q ),
	.datac(!\sig_poa_match_en~q ),
	.datad(!\sig_poa_match~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_poa_state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_poa_state~0 .extended_lut = "off";
defparam \sig_poa_state~0 .lut_mask = 64'h1115111511151115;
defparam \sig_poa_state~0 .shared_arith = "off";

dffeas \poa_block:sig_poa_state (
	.clk(clk),
	.d(\sig_poa_state~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\poa_block:sig_poa_state~q ),
	.prn(vcc));
defparam \poa_block:sig_poa_state .is_wysiwyg = "true";
defparam \poa_block:sig_poa_state .power_up = "low";

arriaii_lcell_comb \sig_poa_ack~0 (
	.dataa(!\sig_dgrb_state.s_poa_cal~q ),
	.datab(!\poa_block:sig_poa_state~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_poa_ack~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_poa_ack~0 .extended_lut = "off";
defparam \sig_poa_ack~0 .lut_mask = 64'h1111111111111111;
defparam \sig_poa_ack~0 .shared_arith = "off";

dffeas sig_poa_ack(
	.clk(clk),
	.d(\sig_poa_ack~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_poa_ack~q ),
	.prn(vcc));
defparam sig_poa_ack.is_wysiwyg = "true";
defparam sig_poa_ack.power_up = "low";

arriaii_lcell_comb \sig_dgrb_state~34 (
	.dataa(!\sig_dgrb_state.s_adv_wd_lat~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_trk_ack~q ),
	.datad(!\sig_poa_ack~q ),
	.datae(!\sig_dgrb_state.s_adv_rd_lat~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~34 .extended_lut = "off";
defparam \sig_dgrb_state~34 .lut_mask = 64'h028A0000028A0000;
defparam \sig_dgrb_state~34 .shared_arith = "off";

arriaii_lcell_comb \sig_dgrb_state~35 (
	.dataa(!\sig_dimm_driving_dq~q ),
	.datab(!\sig_dgrb_state.s_adv_wd_lat~q ),
	.datac(!rdata_valid[0]),
	.datad(!seq_rdata_valid_1),
	.datae(!\sig_dgrb_state.s_adv_rd_lat~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~35 .extended_lut = "off";
defparam \sig_dgrb_state~35 .lut_mask = 64'h02220FFF02220FFF;
defparam \sig_dgrb_state~35 .shared_arith = "off";

dffeas \ctrl_dgrb_r.command.cmd_poa (
	.clk(clk),
	.d(\ctrl_dgrb.command.cmd_poa ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_dgrb_r.command.cmd_poa~q ),
	.prn(vcc));
defparam \ctrl_dgrb_r.command.cmd_poa .is_wysiwyg = "true";
defparam \ctrl_dgrb_r.command.cmd_poa .power_up = "low";

arriaii_lcell_comb \sig_dgrb_state~60 (
	.dataa(!\sig_dgrb_state.s_wait_admin~q ),
	.datab(!\sig_dgrb_state.s_poa_cal~q ),
	.datac(!\sig_dgrb_state~45_combout ),
	.datad(!\ctrl_dgrb_r.command.cmd_poa~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~60_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~60 .extended_lut = "off";
defparam \sig_dgrb_state~60 .lut_mask = 64'h0207020702070207;
defparam \sig_dgrb_state~60 .shared_arith = "off";

dffeas \sig_dgrb_state.s_poa_cal (
	.clk(clk),
	.d(\sig_dgrb_state~60_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgrb_state.s_poa_cal~q ),
	.prn(vcc));
defparam \sig_dgrb_state.s_poa_cal .is_wysiwyg = "true";
defparam \sig_dgrb_state.s_poa_cal .power_up = "low";

arriaii_lcell_comb \sig_dgrb_state~36 (
	.dataa(!\sig_dgrb_state.s_adv_wd_lat~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_state.s_adv_rd_lat~q ),
	.datad(!\sig_dgrb_state.s_poa_cal~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~36 .extended_lut = "off";
defparam \sig_dgrb_state~36 .lut_mask = 64'h8000800080008000;
defparam \sig_dgrb_state~36 .shared_arith = "off";

arriaii_lcell_comb \sig_dgrb_state~37 (
	.dataa(!\sig_dgrb_state.s_rdata_valid_align~q ),
	.datab(!\sig_dgrb_state~34_combout ),
	.datac(!\sig_dgrb_state~35_combout ),
	.datad(!\sig_dgrb_state~36_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~37 .extended_lut = "off";
defparam \sig_dgrb_state~37 .lut_mask = 64'h2A002A002A002A00;
defparam \sig_dgrb_state~37 .shared_arith = "off";

arriaii_lcell_comb \sig_dgrb_state~67 (
	.dataa(!\sig_dgrb_state~38_combout ),
	.datab(!\sig_dimm_driving_dq~q ),
	.datac(!sig_doing_rd_4),
	.datad(!\sig_dgrb_state.s_rdata_valid_align~q ),
	.datae(!\sig_dgrb_state.s_adv_rd_lat_setup~q ),
	.dataf(!\v_aligned~0_combout ),
	.datag(!\sig_dgrb_state~37_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~67_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~67 .extended_lut = "on";
defparam \sig_dgrb_state~67 .lut_mask = 64'h5F5F5D555FFF5DFF;
defparam \sig_dgrb_state~67 .shared_arith = "off";

arriaii_lcell_comb \sig_dgrb_state~39 (
	.dataa(!\sig_dimm_driving_dq~q ),
	.datab(!rdata_valid[0]),
	.datac(!seq_rdata_valid_1),
	.datad(!\sig_dgrb_state.s_adv_rd_lat~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~39 .extended_lut = "off";
defparam \sig_dgrb_state~39 .lut_mask = 64'h2AAA2AAA2AAA2AAA;
defparam \sig_dgrb_state~39 .shared_arith = "off";

arriaii_lcell_comb \sig_dgrb_state~40 (
	.dataa(!\sig_dimm_driving_dq~q ),
	.datab(!\sig_dgrb_state.s_rdata_valid_align~q ),
	.datac(!\sig_dgrb_state.s_idle~q ),
	.datad(!\sig_dgrb_state~39_combout ),
	.datae(!ac_muxctrl_broadcast_rcommand_req),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~40 .extended_lut = "off";
defparam \sig_dgrb_state~40 .lut_mask = 64'h3330131033301310;
defparam \sig_dgrb_state~40 .shared_arith = "off";

dffeas \sig_dgrb_last_state.s_adv_rd_lat_setup (
	.clk(clk),
	.d(\sig_dgrb_state.s_adv_rd_lat_setup~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgrb_last_state.s_adv_rd_lat_setup~q ),
	.prn(vcc));
defparam \sig_dgrb_last_state.s_adv_rd_lat_setup .is_wysiwyg = "true";
defparam \sig_dgrb_last_state.s_adv_rd_lat_setup .power_up = "low";

arriaii_lcell_comb \sig_dgrb_state~41 (
	.dataa(!\sig_dgrb_last_state.s_adv_wd_lat~q ),
	.datab(!\sig_dgrb_state.s_adv_wd_lat~q ),
	.datac(!\sig_dgrb_state.s_wait_admin~q ),
	.datad(!\sig_dgrb_state.s_release_admin~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~41 .extended_lut = "off";
defparam \sig_dgrb_state~41 .lut_mask = 64'hD000D000D000D000;
defparam \sig_dgrb_state~41 .shared_arith = "off";

arriaii_lcell_comb \sig_dgrb_state~42 (
	.dataa(!\sig_dimm_driving_dq~q ),
	.datab(!\sig_dgrb_state.s_idle~q ),
	.datac(!\sig_dgrb_state.s_adv_rd_lat~q ),
	.datad(!ac_muxctrl_broadcast_rcommand_req),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~42 .extended_lut = "off";
defparam \sig_dgrb_state~42 .lut_mask = 64'hCD01CD01CD01CD01;
defparam \sig_dgrb_state~42 .shared_arith = "off";

arriaii_lcell_comb \sig_dgrb_state~43 (
	.dataa(!\sig_dgrb_state.s_adv_rd_lat_setup~q ),
	.datab(!\sig_dgrb_state~40_combout ),
	.datac(!\sig_dgrb_last_state.s_adv_rd_lat_setup~q ),
	.datad(!\sig_dgrb_state~41_combout ),
	.datae(!\sig_dgrb_state~42_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~43 .extended_lut = "off";
defparam \sig_dgrb_state~43 .lut_mask = 64'h008C0000008C0000;
defparam \sig_dgrb_state~43 .shared_arith = "off";

arriaii_lcell_comb \sig_dgrb_state~44 (
	.dataa(!\sig_dimm_driving_dq~q ),
	.datab(!dgb_ac_access_gnt_r),
	.datac(!\sig_dgrb_state.s_release_admin~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~44 .extended_lut = "off";
defparam \sig_dgrb_state~44 .lut_mask = 64'h0404040404040404;
defparam \sig_dgrb_state~44 .shared_arith = "off";

arriaii_lcell_comb \sig_dgrb_state~45 (
	.dataa(!WideOr2),
	.datab(!\sig_dgrb_state.s_idle~q ),
	.datac(!\sig_dgrb_state~67_combout ),
	.datad(!\sig_dgrb_state~43_combout ),
	.datae(!\dgrb_state_proc~0_combout ),
	.dataf(!\sig_dgrb_state~44_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~45 .extended_lut = "off";
defparam \sig_dgrb_state~45 .lut_mask = 64'hFFB8000000000000;
defparam \sig_dgrb_state~45 .shared_arith = "off";

dffeas \ctrl_dgrb_r.command.cmd_rrp_sweep (
	.clk(clk),
	.d(\ctrl_dgrb.command.cmd_rrp_sweep ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_dgrb_r.command.cmd_rrp_sweep~q ),
	.prn(vcc));
defparam \ctrl_dgrb_r.command.cmd_rrp_sweep .is_wysiwyg = "true";
defparam \ctrl_dgrb_r.command.cmd_rrp_sweep .power_up = "low";

arriaii_lcell_comb \sig_dgrb_state~50 (
	.dataa(!\sig_dgrb_state.s_test_phases~q ),
	.datab(!\sig_dgrb_state.s_wait_admin~q ),
	.datac(!\sig_dgrb_state~45_combout ),
	.datad(!\ctrl_dgrb_r.command.cmd_rrp_sweep~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~50_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~50 .extended_lut = "off";
defparam \sig_dgrb_state~50 .lut_mask = 64'h0407040704070407;
defparam \sig_dgrb_state~50 .shared_arith = "off";

dffeas \sig_dgrb_state.s_test_phases (
	.clk(clk),
	.d(\sig_dgrb_state~50_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgrb_state.s_test_phases~q ),
	.prn(vcc));
defparam \sig_dgrb_state.s_test_phases .is_wysiwyg = "true";
defparam \sig_dgrb_state.s_test_phases .power_up = "low";

arriaii_lcell_comb \Selector25~0 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_dgrb_state.s_wait_admin~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector25~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector25~0 .extended_lut = "off";
defparam \Selector25~0 .lut_mask = 64'h8080808080808080;
defparam \Selector25~0 .shared_arith = "off";

arriaii_lcell_comb \Selector25~1 (
	.dataa(!\sig_dgrb_state.s_seek_cdvw~q ),
	.datab(!\sig_dgrb_state.s_test_phases~q ),
	.datac(!\sig_rsc_ack~q ),
	.datad(!\sig_dgrb_state.s_read_mtp~q ),
	.datae(!\Selector25~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector25~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector25~1 .extended_lut = "off";
defparam \Selector25~1 .lut_mask = 64'h0000A8000000A800;
defparam \Selector25~1 .shared_arith = "off";

arriaii_lcell_comb \sig_rsc_ac_access_req~0 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_flush_datapath~q ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_test_dq~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_rsc_ac_access_req~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_rsc_ac_access_req~0 .extended_lut = "off";
defparam \sig_rsc_ac_access_req~0 .lut_mask = 64'h7777777777777777;
defparam \sig_rsc_ac_access_req~0 .shared_arith = "off";

dffeas sig_rsc_ac_access_req(
	.clk(clk),
	.d(\sig_rsc_ac_access_req~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_rsc_ac_access_req~q ),
	.prn(vcc));
defparam sig_rsc_ac_access_req.is_wysiwyg = "true";
defparam sig_rsc_ac_access_req.power_up = "low";

arriaii_lcell_comb \Selector21~0 (
	.dataa(!\sig_ac_req.s_ac_idle~q ),
	.datab(!\sig_dgrb_state.s_idle~q ),
	.datac(!\sig_dgrb_state.s_release_admin~q ),
	.datad(!\Selector25~1_combout ),
	.datae(!\sig_rsc_ac_access_req~q ),
	.dataf(!\Selector23~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector21~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector21~0 .extended_lut = "off";
defparam \Selector21~0 .lut_mask = 64'h1030103000001030;
defparam \Selector21~0 .shared_arith = "off";

dffeas \sig_ac_req.s_ac_idle (
	.clk(clk),
	.d(\Selector21~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_ac_req.s_ac_idle~q ),
	.prn(vcc));
defparam \sig_ac_req.s_ac_idle .is_wysiwyg = "true";
defparam \sig_ac_req.s_ac_idle .power_up = "low";

arriaii_lcell_comb \sig_addr_cmd_state~5 (
	.dataa(!\Equal21~0_combout ),
	.datab(!\ac_block:sig_addr_cmd_state.s_ac_idle~q ),
	.datac(!\ac_block:sig_addr_cmd_state.s_ac_relax~q ),
	.datad(!\ac_block:sig_addr_cmd_last_state.s_ac_relax~q ),
	.datae(!\sig_ac_req.s_ac_idle~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_addr_cmd_state~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_addr_cmd_state~5 .extended_lut = "off";
defparam \sig_addr_cmd_state~5 .lut_mask = 64'h3332FFFA3332FFFA;
defparam \sig_addr_cmd_state~5 .shared_arith = "off";

dffeas \ac_block:sig_addr_cmd_state.s_ac_idle (
	.clk(clk),
	.d(\sig_addr_cmd_state~5_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_block:sig_addr_cmd_state.s_ac_idle~q ),
	.prn(vcc));
defparam \ac_block:sig_addr_cmd_state.s_ac_idle .is_wysiwyg = "true";
defparam \ac_block:sig_addr_cmd_state.s_ac_idle .power_up = "low";

arriaii_lcell_comb \Selector25~2 (
	.dataa(!\sig_ac_req.s_ac_read_poa_mtp~q ),
	.datab(!\sig_dgrb_state.s_poa_cal~q ),
	.datac(!\Selector25~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector25~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector25~2 .extended_lut = "off";
defparam \Selector25~2 .lut_mask = 64'h7373737373737373;
defparam \Selector25~2 .shared_arith = "off";

dffeas \sig_ac_req.s_ac_read_poa_mtp (
	.clk(clk),
	.d(\Selector25~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_ac_req.s_ac_read_poa_mtp~q ),
	.prn(vcc));
defparam \sig_ac_req.s_ac_read_poa_mtp .is_wysiwyg = "true";
defparam \sig_ac_req.s_ac_read_poa_mtp .power_up = "low";

arriaii_lcell_comb \Selector26~0 (
	.dataa(!\sig_dgrb_state.s_adv_wd_lat~q ),
	.datab(!\sig_ac_req.s_ac_read_wd_lat~q ),
	.datac(!\Selector25~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector26~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector26~0 .extended_lut = "off";
defparam \Selector26~0 .lut_mask = 64'h7575757575757575;
defparam \Selector26~0 .shared_arith = "off";

dffeas \sig_ac_req.s_ac_read_wd_lat (
	.clk(clk),
	.d(\Selector26~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_ac_req.s_ac_read_wd_lat~q ),
	.prn(vcc));
defparam \sig_ac_req.s_ac_read_wd_lat .is_wysiwyg = "true";
defparam \sig_ac_req.s_ac_read_wd_lat .power_up = "low";

arriaii_lcell_comb \ac_proc~0 (
	.dataa(!\ac_block:sig_addr_cmd_state.s_ac_read_wd_lat~q ),
	.datab(!\ac_block:sig_addr_cmd_state.s_ac_relax~q ),
	.datac(!\sig_ac_req.s_ac_read_wd_lat~q ),
	.datad(!\sig_ac_req.s_ac_idle~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_proc~0 .extended_lut = "off";
defparam \ac_proc~0 .lut_mask = 64'h0084008400840084;
defparam \ac_proc~0 .shared_arith = "off";

arriaii_lcell_comb \sig_addr_cmd_state~0 (
	.dataa(!\Equal21~0_combout ),
	.datab(!\ac_block:sig_addr_cmd_state.s_ac_relax~q ),
	.datac(!\ac_block:sig_addr_cmd_last_state.s_ac_relax~q ),
	.datad(!\ac_proc~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_addr_cmd_state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_addr_cmd_state~0 .extended_lut = "off";
defparam \sig_addr_cmd_state~0 .lut_mask = 64'hFE00FE00FE00FE00;
defparam \sig_addr_cmd_state~0 .shared_arith = "off";

arriaii_lcell_comb \sig_addr_cmd_state~4 (
	.dataa(!\sig_ac_req.s_ac_read_rdv~q ),
	.datab(!\sig_addr_cmd_state~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_addr_cmd_state~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_addr_cmd_state~4 .extended_lut = "off";
defparam \sig_addr_cmd_state~4 .lut_mask = 64'h1111111111111111;
defparam \sig_addr_cmd_state~4 .shared_arith = "off";

dffeas \ac_block:sig_addr_cmd_state.s_ac_read_rdv (
	.clk(clk),
	.d(\sig_addr_cmd_state~4_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ),
	.prn(vcc));
defparam \ac_block:sig_addr_cmd_state.s_ac_read_rdv .is_wysiwyg = "true";
defparam \ac_block:sig_addr_cmd_state.s_ac_read_rdv .power_up = "low";

arriaii_lcell_comb \Selector24~0 (
	.dataa(!\sig_dgrb_state.s_rdata_valid_align~q ),
	.datab(!\sig_ac_req.s_ac_read_rdv~q ),
	.datac(!\sig_dgrb_state.s_adv_rd_lat_setup~q ),
	.datad(!\sig_dgrb_state.s_adv_rd_lat~q ),
	.datae(!\Selector25~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector24~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector24~0 .extended_lut = "off";
defparam \Selector24~0 .lut_mask = 64'h7FFF5FFF7FFF5FFF;
defparam \Selector24~0 .shared_arith = "off";

dffeas \sig_ac_req.s_ac_read_rdv (
	.clk(clk),
	.d(\Selector24~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_ac_req.s_ac_read_rdv~q ),
	.prn(vcc));
defparam \sig_ac_req.s_ac_read_rdv .is_wysiwyg = "true";
defparam \sig_ac_req.s_ac_read_rdv .power_up = "low";

arriaii_lcell_comb \Selector23~1 (
	.dataa(!\sig_ac_req.s_ac_read_mtp~q ),
	.datab(!\Selector25~1_combout ),
	.datac(!\sig_rsc_ac_access_req~q ),
	.datad(!\Selector23~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector23~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector23~1 .extended_lut = "off";
defparam \Selector23~1 .lut_mask = 64'h444F444F444F444F;
defparam \Selector23~1 .shared_arith = "off";

dffeas \sig_ac_req.s_ac_read_mtp (
	.clk(clk),
	.d(\Selector23~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_ac_req.s_ac_read_mtp~q ),
	.prn(vcc));
defparam \sig_ac_req.s_ac_read_mtp .is_wysiwyg = "true";
defparam \sig_ac_req.s_ac_read_mtp .power_up = "low";

arriaii_lcell_comb \ac_proc~1 (
	.dataa(!\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.datab(!\ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ),
	.datac(!\sig_ac_req.s_ac_read_rdv~q ),
	.datad(!\sig_ac_req.s_ac_read_mtp~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_proc~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_proc~1 .extended_lut = "off";
defparam \ac_proc~1 .lut_mask = 64'h8241824182418241;
defparam \ac_proc~1 .shared_arith = "off";

arriaii_lcell_comb \ac_proc~2 (
	.dataa(!\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.datab(!\ac_block:sig_addr_cmd_state.s_ac_idle~q ),
	.datac(!\sig_ac_req.s_ac_read_poa_mtp~q ),
	.datad(!\ac_proc~0_combout ),
	.datae(!\ac_proc~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_proc~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_proc~2 .extended_lut = "off";
defparam \ac_proc~2 .lut_mask = 64'h3333331233333312;
defparam \ac_proc~2 .shared_arith = "off";

arriaii_lcell_comb \sig_addr_cmd_state~6 (
	.dataa(!\Equal21~0_combout ),
	.datab(!\ac_block:sig_addr_cmd_state.s_ac_relax~q ),
	.datac(!\ac_block:sig_addr_cmd_last_state.s_ac_relax~q ),
	.datad(!\ac_proc~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_addr_cmd_state~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_addr_cmd_state~6 .extended_lut = "off";
defparam \sig_addr_cmd_state~6 .lut_mask = 64'h00FE00FE00FE00FE;
defparam \sig_addr_cmd_state~6 .shared_arith = "off";

dffeas \ac_block:sig_addr_cmd_state.s_ac_relax (
	.clk(clk),
	.d(\sig_addr_cmd_state~6_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_block:sig_addr_cmd_state.s_ac_relax~q ),
	.prn(vcc));
defparam \ac_block:sig_addr_cmd_state.s_ac_relax .is_wysiwyg = "true";
defparam \ac_block:sig_addr_cmd_state.s_ac_relax .power_up = "low";

arriaii_lcell_comb \Add22~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\ac_block:sig_setup[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add22~1_sumout ),
	.cout(\Add22~2 ),
	.shareout());
defparam \Add22~1 .extended_lut = "off";
defparam \Add22~1 .lut_mask = 64'h000000000000FF00;
defparam \Add22~1 .shared_arith = "off";

arriaii_lcell_comb \sig_setup~0 (
	.dataa(!dgb_ac_access_gnt_r),
	.datab(!\Add22~1_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_setup~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_setup~0 .extended_lut = "off";
defparam \sig_setup~0 .lut_mask = 64'h4444444444444444;
defparam \sig_setup~0 .shared_arith = "off";

arriaii_lcell_comb \ac_block:sig_setup[4]~0 (
	.dataa(!\dimm_driving_dq_proc~0_combout ),
	.datab(!\Selector141~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_block:sig_setup[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_block:sig_setup[4]~0 .extended_lut = "off";
defparam \ac_block:sig_setup[4]~0 .lut_mask = 64'h4444444444444444;
defparam \ac_block:sig_setup[4]~0 .shared_arith = "off";

dffeas \ac_block:sig_setup[0] (
	.clk(clk),
	.d(\sig_setup~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ac_block:sig_setup[4]~0_combout ),
	.q(\ac_block:sig_setup[0]~q ),
	.prn(vcc));
defparam \ac_block:sig_setup[0] .is_wysiwyg = "true";
defparam \ac_block:sig_setup[0] .power_up = "low";

arriaii_lcell_comb \Add22~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\ac_block:sig_setup[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add22~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add22~5_sumout ),
	.cout(\Add22~6 ),
	.shareout());
defparam \Add22~5 .extended_lut = "off";
defparam \Add22~5 .lut_mask = 64'h000000000000FF00;
defparam \Add22~5 .shared_arith = "off";

arriaii_lcell_comb \sig_setup~1 (
	.dataa(!dgb_ac_access_gnt_r),
	.datab(!\Add22~5_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_setup~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_setup~1 .extended_lut = "off";
defparam \sig_setup~1 .lut_mask = 64'h4444444444444444;
defparam \sig_setup~1 .shared_arith = "off";

dffeas \ac_block:sig_setup[1] (
	.clk(clk),
	.d(\sig_setup~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ac_block:sig_setup[4]~0_combout ),
	.q(\ac_block:sig_setup[1]~q ),
	.prn(vcc));
defparam \ac_block:sig_setup[1] .is_wysiwyg = "true";
defparam \ac_block:sig_setup[1] .power_up = "low";

arriaii_lcell_comb \Add22~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\ac_block:sig_setup[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add22~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add22~9_sumout ),
	.cout(\Add22~10 ),
	.shareout());
defparam \Add22~9 .extended_lut = "off";
defparam \Add22~9 .lut_mask = 64'h000000000000FF00;
defparam \Add22~9 .shared_arith = "off";

arriaii_lcell_comb \sig_setup~2 (
	.dataa(!dgb_ac_access_gnt_r),
	.datab(!\Add22~9_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_setup~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_setup~2 .extended_lut = "off";
defparam \sig_setup~2 .lut_mask = 64'h4444444444444444;
defparam \sig_setup~2 .shared_arith = "off";

dffeas \ac_block:sig_setup[2] (
	.clk(clk),
	.d(\sig_setup~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ac_block:sig_setup[4]~0_combout ),
	.q(\ac_block:sig_setup[2]~q ),
	.prn(vcc));
defparam \ac_block:sig_setup[2] .is_wysiwyg = "true";
defparam \ac_block:sig_setup[2] .power_up = "low";

arriaii_lcell_comb \Add22~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\ac_block:sig_setup[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add22~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add22~13_sumout ),
	.cout(\Add22~14 ),
	.shareout());
defparam \Add22~13 .extended_lut = "off";
defparam \Add22~13 .lut_mask = 64'h000000000000FF00;
defparam \Add22~13 .shared_arith = "off";

arriaii_lcell_comb \sig_setup~3 (
	.dataa(!dgb_ac_access_gnt_r),
	.datab(!\Add22~13_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_setup~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_setup~3 .extended_lut = "off";
defparam \sig_setup~3 .lut_mask = 64'h4444444444444444;
defparam \sig_setup~3 .shared_arith = "off";

dffeas \ac_block:sig_setup[3] (
	.clk(clk),
	.d(\sig_setup~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ac_block:sig_setup[4]~0_combout ),
	.q(\ac_block:sig_setup[3]~q ),
	.prn(vcc));
defparam \ac_block:sig_setup[3] .is_wysiwyg = "true";
defparam \ac_block:sig_setup[3] .power_up = "low";

arriaii_lcell_comb \Add22~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\ac_block:sig_setup[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add22~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add22~17_sumout ),
	.cout(),
	.shareout());
defparam \Add22~17 .extended_lut = "off";
defparam \Add22~17 .lut_mask = 64'h000000000000FF00;
defparam \Add22~17 .shared_arith = "off";

arriaii_lcell_comb \sig_setup~4 (
	.dataa(!dgb_ac_access_gnt_r),
	.datab(!\Add22~17_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_setup~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_setup~4 .extended_lut = "off";
defparam \sig_setup~4 .lut_mask = 64'h4444444444444444;
defparam \sig_setup~4 .shared_arith = "off";

dffeas \ac_block:sig_setup[4] (
	.clk(clk),
	.d(\sig_setup~4_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ac_block:sig_setup[4]~0_combout ),
	.q(\ac_block:sig_setup[4]~q ),
	.prn(vcc));
defparam \ac_block:sig_setup[4] .is_wysiwyg = "true";
defparam \ac_block:sig_setup[4] .power_up = "low";

arriaii_lcell_comb \Selector141~0 (
	.dataa(!dgb_ac_access_gnt_r),
	.datab(!\ac_block:sig_setup[0]~q ),
	.datac(!\ac_block:sig_setup[1]~q ),
	.datad(!\ac_block:sig_setup[2]~q ),
	.datae(!\ac_block:sig_setup[3]~q ),
	.dataf(!\ac_block:sig_setup[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector141~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector141~0 .extended_lut = "off";
defparam \Selector141~0 .lut_mask = 64'h0000000000000001;
defparam \Selector141~0 .shared_arith = "off";

arriaii_lcell_comb \Selector141~1 (
	.dataa(!\ac_block:sig_addr_cmd_state.s_ac_idle~q ),
	.datab(!\ac_block:sig_addr_cmd_state.s_ac_relax~q ),
	.datac(!\Selector141~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector141~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector141~1 .extended_lut = "off";
defparam \Selector141~1 .lut_mask = 64'hC8C8C8C8C8C8C8C8;
defparam \Selector141~1 .shared_arith = "off";

dffeas sig_dimm_driving_dq(
	.clk(clk),
	.d(\Selector141~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dimm_driving_dq~q ),
	.prn(vcc));
defparam sig_dimm_driving_dq.is_wysiwyg = "true";
defparam sig_dimm_driving_dq.power_up = "low";

arriaii_lcell_comb \sig_dgrb_state~58 (
	.dataa(!sig_doing_rd_4),
	.datab(!\sig_dimm_driving_dq~q ),
	.datac(!\sig_dgrb_state.s_adv_rd_lat_setup~q ),
	.datad(!\sig_dgrb_last_state.s_adv_rd_lat_setup~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~58_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~58 .extended_lut = "off";
defparam \sig_dgrb_state~58 .lut_mask = 64'h0004000400040004;
defparam \sig_dgrb_state~58 .shared_arith = "off";

arriaii_lcell_comb \sig_dgrb_state~59 (
	.dataa(!\sig_dimm_driving_dq~q ),
	.datab(!rdata_valid[0]),
	.datac(!seq_rdata_valid_1),
	.datad(!\sig_dgrb_state.s_adv_rd_lat~q ),
	.datae(!\dgrb_state_proc~0_combout ),
	.dataf(!\sig_dgrb_state~58_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~59_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~59 .extended_lut = "off";
defparam \sig_dgrb_state~59 .lut_mask = 64'h00D50000FFFF0000;
defparam \sig_dgrb_state~59 .shared_arith = "off";

dffeas \sig_dgrb_state.s_adv_rd_lat (
	.clk(clk),
	.d(\sig_dgrb_state~59_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgrb_state.s_adv_rd_lat~q ),
	.prn(vcc));
defparam \sig_dgrb_state.s_adv_rd_lat .is_wysiwyg = "true";
defparam \sig_dgrb_state.s_adv_rd_lat .power_up = "low";

dffeas \ctrl_dgrb_r.command.cmd_rrp_reset (
	.clk(clk),
	.d(\ctrl_dgrb.command.cmd_rrp_reset ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_dgrb_r.command.cmd_rrp_reset~q ),
	.prn(vcc));
defparam \ctrl_dgrb_r.command.cmd_rrp_reset .is_wysiwyg = "true";
defparam \ctrl_dgrb_r.command.cmd_rrp_reset .power_up = "low";

arriaii_lcell_comb \sig_dgrb_state~49 (
	.dataa(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datab(!\sig_dgrb_state.s_wait_admin~q ),
	.datac(!\sig_dgrb_state~45_combout ),
	.datad(!\ctrl_dgrb_r.command.cmd_rrp_reset~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~49 .extended_lut = "off";
defparam \sig_dgrb_state~49 .lut_mask = 64'h0407040704070407;
defparam \sig_dgrb_state~49 .shared_arith = "off";

dffeas \sig_dgrb_state.s_reset_cdvw (
	.clk(clk),
	.d(\sig_dgrb_state~49_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgrb_state.s_reset_cdvw~q ),
	.prn(vcc));
defparam \sig_dgrb_state.s_reset_cdvw .is_wysiwyg = "true";
defparam \sig_dgrb_state.s_reset_cdvw .power_up = "low";

arriaii_lcell_comb \sig_dgrb_state~38 (
	.dataa(!\sig_dgrb_state.s_seek_cdvw~q ),
	.datab(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datac(!\sig_dgrb_state.s_test_phases~q ),
	.datad(!\sig_rsc_ack~q ),
	.datae(!\sig_dgrb_state.s_read_mtp~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~38 .extended_lut = "off";
defparam \sig_dgrb_state~38 .lut_mask = 64'h007F00FF007F00FF;
defparam \sig_dgrb_state~38 .shared_arith = "off";

arriaii_lcell_comb \sig_dgrb_state~62 (
	.dataa(!\v_aligned~0_combout ),
	.datab(!\sig_dgrb_state.s_rdata_valid_align~q ),
	.datac(!\sig_dgrb_state~38_combout ),
	.datad(!\sig_dgrb_state~39_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~62_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~62 .extended_lut = "off";
defparam \sig_dgrb_state~62 .lut_mask = 64'h0C1F0C1F0C1F0C1F;
defparam \sig_dgrb_state~62 .shared_arith = "off";

arriaii_lcell_comb \sig_dgrb_state~63 (
	.dataa(!\sig_dgrb_last_state.s_adv_wd_lat~q ),
	.datab(!\sig_dgrb_state.s_adv_wd_lat~q ),
	.datac(!\sig_dgrb_state.s_idle~q ),
	.datad(!\sig_dgrb_state.s_adv_rd_lat_setup~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~63_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~63 .extended_lut = "off";
defparam \sig_dgrb_state~63 .lut_mask = 64'h0D000D000D000D00;
defparam \sig_dgrb_state~63 .shared_arith = "off";

arriaii_lcell_comb \sig_dgrb_state~64 (
	.dataa(!\sig_dimm_driving_dq~q ),
	.datab(!\sig_dgrb_state.s_adv_rd_lat~q ),
	.datac(!\sig_dgrb_state~37_combout ),
	.datad(!\sig_dgrb_state~62_combout ),
	.datae(!\sig_dgrb_state~63_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~64_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~64 .extended_lut = "off";
defparam \sig_dgrb_state~64 .lut_mask = 64'h00000EEE00000EEE;
defparam \sig_dgrb_state~64 .shared_arith = "off";

arriaii_lcell_comb \sig_dgrb_state~65 (
	.dataa(!\sig_dgrb_state.s_wait_admin~q ),
	.datab(!\sig_dgrb_state~44_combout ),
	.datac(!\sig_dgrb_state~58_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~65_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~65 .extended_lut = "off";
defparam \sig_dgrb_state~65 .lut_mask = 64'h8080808080808080;
defparam \sig_dgrb_state~65 .shared_arith = "off";

arriaii_lcell_comb \sig_dgrb_state~66 (
	.dataa(!\sig_dgrb_state.s_release_admin~q ),
	.datab(!\dgrb_state_proc~0_combout ),
	.datac(!\sig_dgrb_state~56_combout ),
	.datad(!\sig_dgrb_state~64_combout ),
	.datae(!\sig_dgrb_state~65_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~66_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~66 .extended_lut = "off";
defparam \sig_dgrb_state~66 .lut_mask = 64'h333373F3333373F3;
defparam \sig_dgrb_state~66 .shared_arith = "off";

dffeas \sig_dgrb_state.s_release_admin (
	.clk(clk),
	.d(\sig_dgrb_state~66_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgrb_state.s_release_admin~q ),
	.prn(vcc));
defparam \sig_dgrb_state.s_release_admin .is_wysiwyg = "true";
defparam \sig_dgrb_state.s_release_admin .power_up = "low";

arriaii_lcell_comb \dgrb_state_proc~0 (
	.dataa(!curr_cmdcmd_idle),
	.datab(!\sig_dgrb_state.s_idle~q ),
	.datac(!\sig_dgrb_state.s_release_admin~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dgrb_state_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dgrb_state_proc~0 .extended_lut = "off";
defparam \dgrb_state_proc~0 .lut_mask = 64'h2020202020202020;
defparam \dgrb_state_proc~0 .shared_arith = "off";

arriaii_lcell_comb \sig_dgrb_state~52 (
	.dataa(!\sig_dgrb_state.s_wait_admin~q ),
	.datab(!\ctrl_dgrb_r.command.cmd_read_mtp~q ),
	.datac(!\ctrl_dgrb_r.command.cmd_rrp_reset~q ),
	.datad(!\ctrl_dgrb_r.command.cmd_rrp_sweep~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~52 .extended_lut = "off";
defparam \sig_dgrb_state~52 .lut_mask = 64'h4000400040004000;
defparam \sig_dgrb_state~52 .shared_arith = "off";

arriaii_lcell_comb \sig_dgrb_state~53 (
	.dataa(!\ctrl_dgrb_r.command.cmd_prep_adv_wr_lat~q ),
	.datab(!\ctrl_dgrb_r.command.cmd_tr_due~q ),
	.datac(!\ctrl_dgrb_r.command.cmd_poa~q ),
	.datad(!\ctrl_dgrb_r.command.cmd_prep_adv_rd_lat~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~53_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~53 .extended_lut = "off";
defparam \sig_dgrb_state~53 .lut_mask = 64'h8000800080008000;
defparam \sig_dgrb_state~53 .shared_arith = "off";

arriaii_lcell_comb \sig_dgrb_state~54 (
	.dataa(!\sig_dgrb_state~44_combout ),
	.datab(!\ctrl_dgrb_r.command.cmd_rdv~q ),
	.datac(!\ctrl_dgrb_r.command.cmd_rrp_seek~q ),
	.datad(!\sig_dgrb_state~52_combout ),
	.datae(!\sig_dgrb_state~53_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~54_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~54 .extended_lut = "off";
defparam \sig_dgrb_state~54 .lut_mask = 64'hAAAAAA2AAAAAAA2A;
defparam \sig_dgrb_state~54 .shared_arith = "off";

arriaii_lcell_comb \sig_dgrb_state~55 (
	.dataa(!WideOr2),
	.datab(!\sig_dgrb_state.s_idle~q ),
	.datac(!\sig_dgrb_state.s_wait_admin~q ),
	.datad(!ac_muxctrl_broadcast_rcommand_req),
	.datae(!\dgrb_state_proc~0_combout ),
	.dataf(!\sig_dgrb_state~54_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~55_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~55 .extended_lut = "off";
defparam \sig_dgrb_state~55 .lut_mask = 64'h0000FFFF3F7FFFFF;
defparam \sig_dgrb_state~55 .shared_arith = "off";

dffeas \sig_dgrb_state.s_idle (
	.clk(clk),
	.d(\sig_dgrb_state~55_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgrb_state.s_idle~q ),
	.prn(vcc));
defparam \sig_dgrb_state.s_idle .is_wysiwyg = "true";
defparam \sig_dgrb_state.s_idle .power_up = "low";

arriaii_lcell_comb \sig_dgrb_state~56 (
	.dataa(!curr_ctrlcommand_ack),
	.datab(!curr_cmdcmd_idle),
	.datac(!WideOr0),
	.datad(!\sig_dgrb_state.s_idle~q ),
	.datae(!ac_muxctrl_broadcast_rcommand_req),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~56_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~56 .extended_lut = "off";
defparam \sig_dgrb_state~56 .lut_mask = 64'h0000010000000100;
defparam \sig_dgrb_state~56 .shared_arith = "off";

dffeas \sig_dgrb_state.s_wait_admin (
	.clk(clk),
	.d(\sig_dgrb_state~56_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgrb_state.s_wait_admin~q ),
	.prn(vcc));
defparam \sig_dgrb_state.s_wait_admin .is_wysiwyg = "true";
defparam \sig_dgrb_state.s_wait_admin .power_up = "low";

dffeas \ctrl_dgrb_r.command.cmd_prep_adv_wr_lat (
	.clk(clk),
	.d(\ctrl_dgrb.command.cmd_prep_adv_wr_lat ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_dgrb_r.command.cmd_prep_adv_wr_lat~q ),
	.prn(vcc));
defparam \ctrl_dgrb_r.command.cmd_prep_adv_wr_lat .is_wysiwyg = "true";
defparam \ctrl_dgrb_r.command.cmd_prep_adv_wr_lat .power_up = "low";

arriaii_lcell_comb \sig_dgrb_state~46 (
	.dataa(!\sig_dgrb_state.s_adv_wd_lat~q ),
	.datab(!\sig_dgrb_state.s_wait_admin~q ),
	.datac(!\ctrl_dgrb_r.command.cmd_prep_adv_wr_lat~q ),
	.datad(!\sig_dgrb_state~45_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_dgrb_state~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_dgrb_state~46 .extended_lut = "off";
defparam \sig_dgrb_state~46 .lut_mask = 64'h0047004700470047;
defparam \sig_dgrb_state~46 .shared_arith = "off";

dffeas \sig_dgrb_state.s_adv_wd_lat (
	.clk(clk),
	.d(\sig_dgrb_state~46_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgrb_state.s_adv_wd_lat~q ),
	.prn(vcc));
defparam \sig_dgrb_state.s_adv_wd_lat .is_wysiwyg = "true";
defparam \sig_dgrb_state.s_adv_wd_lat .power_up = "low";

dffeas \sig_dgrb_last_state.s_adv_wd_lat (
	.clk(clk),
	.d(\sig_dgrb_state.s_adv_wd_lat~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgrb_last_state.s_adv_wd_lat~q ),
	.prn(vcc));
defparam \sig_dgrb_last_state.s_adv_wd_lat .is_wysiwyg = "true";
defparam \sig_dgrb_last_state.s_adv_wd_lat .power_up = "low";

arriaii_lcell_comb \sig_wd_lat~1 (
	.dataa(!q_b_2),
	.datab(!\sig_dgrb_last_state.s_adv_wd_lat~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_wd_lat~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_wd_lat~1 .extended_lut = "off";
defparam \sig_wd_lat~1 .lut_mask = 64'h1111111111111111;
defparam \sig_wd_lat~1 .shared_arith = "off";

arriaii_lcell_comb \dgrb_main_block:sig_wd_lat[1]~0 (
	.dataa(!\sig_dimm_driving_dq~q ),
	.datab(!\sig_dgrb_last_state.s_adv_wd_lat~q ),
	.datac(!\sig_dgrb_state.s_adv_wd_lat~q ),
	.datad(!rdata_valid[0]),
	.datae(!seq_rdata_valid_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dgrb_main_block:sig_wd_lat[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dgrb_main_block:sig_wd_lat[1]~0 .extended_lut = "off";
defparam \dgrb_main_block:sig_wd_lat[1]~0 .lut_mask = 64'h0C0E0E0E0C0E0E0E;
defparam \dgrb_main_block:sig_wd_lat[1]~0 .shared_arith = "off";

dffeas \dgrb_main_block:sig_wd_lat[2] (
	.clk(clk),
	.d(\sig_wd_lat~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dgrb_main_block:sig_wd_lat[1]~0_combout ),
	.q(\dgrb_main_block:sig_wd_lat[2]~q ),
	.prn(vcc));
defparam \dgrb_main_block:sig_wd_lat[2] .is_wysiwyg = "true";
defparam \dgrb_main_block:sig_wd_lat[2] .power_up = "low";

arriaii_lcell_comb \wd_lat[2]~0 (
	.dataa(!\dgrb_main_block:sig_wd_lat[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wd_lat[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wd_lat[2]~0 .extended_lut = "off";
defparam \wd_lat[2]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \wd_lat[2]~0 .shared_arith = "off";

arriaii_lcell_comb \sig_wd_lat~2 (
	.dataa(!q_b_1),
	.datab(!\sig_dgrb_last_state.s_adv_wd_lat~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_wd_lat~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_wd_lat~2 .extended_lut = "off";
defparam \sig_wd_lat~2 .lut_mask = 64'h1111111111111111;
defparam \sig_wd_lat~2 .shared_arith = "off";

dffeas \dgrb_main_block:sig_wd_lat[1] (
	.clk(clk),
	.d(\sig_wd_lat~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dgrb_main_block:sig_wd_lat[1]~0_combout ),
	.q(\dgrb_main_block:sig_wd_lat[1]~q ),
	.prn(vcc));
defparam \dgrb_main_block:sig_wd_lat[1] .is_wysiwyg = "true";
defparam \dgrb_main_block:sig_wd_lat[1] .power_up = "low";

arriaii_lcell_comb \sig_wd_lat~3 (
	.dataa(!q_b_0),
	.datab(!\sig_dgrb_last_state.s_adv_wd_lat~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_wd_lat~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_wd_lat~3 .extended_lut = "off";
defparam \sig_wd_lat~3 .lut_mask = 64'h1111111111111111;
defparam \sig_wd_lat~3 .shared_arith = "off";

dffeas \dgrb_main_block:sig_wd_lat[0] (
	.clk(clk),
	.d(\sig_wd_lat~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dgrb_main_block:sig_wd_lat[1]~0_combout ),
	.q(\dgrb_main_block:sig_wd_lat[0]~q ),
	.prn(vcc));
defparam \dgrb_main_block:sig_wd_lat[0] .is_wysiwyg = "true";
defparam \dgrb_main_block:sig_wd_lat[0] .power_up = "low";

arriaii_lcell_comb \wd_lat[0]~1 (
	.dataa(!\dgrb_main_block:sig_wd_lat[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wd_lat[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wd_lat[0]~1 .extended_lut = "off";
defparam \wd_lat[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \wd_lat[0]~1 .shared_arith = "off";

arriaii_lcell_comb \sig_wd_lat~4 (
	.dataa(!q_b_3),
	.datab(!\sig_dgrb_last_state.s_adv_wd_lat~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_wd_lat~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_wd_lat~4 .extended_lut = "off";
defparam \sig_wd_lat~4 .lut_mask = 64'h1111111111111111;
defparam \sig_wd_lat~4 .shared_arith = "off";

dffeas \dgrb_main_block:sig_wd_lat[3] (
	.clk(clk),
	.d(\sig_wd_lat~4_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dgrb_main_block:sig_wd_lat[1]~0_combout ),
	.q(\dgrb_main_block:sig_wd_lat[3]~q ),
	.prn(vcc));
defparam \dgrb_main_block:sig_wd_lat[3] .is_wysiwyg = "true";
defparam \dgrb_main_block:sig_wd_lat[3] .power_up = "low";

arriaii_lcell_comb \sig_wd_lat~5 (
	.dataa(!q_b_4),
	.datab(!\sig_dgrb_last_state.s_adv_wd_lat~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_wd_lat~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_wd_lat~5 .extended_lut = "off";
defparam \sig_wd_lat~5 .lut_mask = 64'h1111111111111111;
defparam \sig_wd_lat~5 .shared_arith = "off";

dffeas \dgrb_main_block:sig_wd_lat[4] (
	.clk(clk),
	.d(\sig_wd_lat~5_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dgrb_main_block:sig_wd_lat[1]~0_combout ),
	.q(\dgrb_main_block:sig_wd_lat[4]~q ),
	.prn(vcc));
defparam \dgrb_main_block:sig_wd_lat[4] .is_wysiwyg = "true";
defparam \dgrb_main_block:sig_wd_lat[4] .power_up = "low";

arriaii_lcell_comb \sig_burst_count~0 (
	.dataa(!\ac_block:sig_burst_count[0]~q ),
	.datab(!\ac_block:sig_addr_cmd_state.s_ac_idle~q ),
	.datac(!\ac_block:sig_addr_cmd_state.s_ac_relax~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_burst_count~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_burst_count~0 .extended_lut = "off";
defparam \sig_burst_count~0 .lut_mask = 64'h2020202020202020;
defparam \sig_burst_count~0 .shared_arith = "off";

dffeas \ac_block:sig_burst_count[0] (
	.clk(clk),
	.d(\sig_burst_count~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_block:sig_burst_count[0]~q ),
	.prn(vcc));
defparam \ac_block:sig_burst_count[0] .is_wysiwyg = "true";
defparam \ac_block:sig_burst_count[0] .power_up = "low";

arriaii_lcell_comb \sig_addr_cmd_state~1 (
	.dataa(!\sig_ac_req.s_ac_read_wd_lat~q ),
	.datab(!\sig_addr_cmd_state~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_addr_cmd_state~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_addr_cmd_state~1 .extended_lut = "off";
defparam \sig_addr_cmd_state~1 .lut_mask = 64'h1111111111111111;
defparam \sig_addr_cmd_state~1 .shared_arith = "off";

dffeas \ac_block:sig_addr_cmd_state.s_ac_read_wd_lat (
	.clk(clk),
	.d(\sig_addr_cmd_state~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_block:sig_addr_cmd_state.s_ac_read_wd_lat~q ),
	.prn(vcc));
defparam \ac_block:sig_addr_cmd_state.s_ac_read_wd_lat .is_wysiwyg = "true";
defparam \ac_block:sig_addr_cmd_state.s_ac_read_wd_lat .power_up = "low";

dffeas \ac_block:sig_addr_cmd_last_state.s_ac_read_wd_lat (
	.clk(clk),
	.d(\ac_block:sig_addr_cmd_state.s_ac_read_wd_lat~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_block:sig_addr_cmd_last_state.s_ac_read_wd_lat~q ),
	.prn(vcc));
defparam \ac_block:sig_addr_cmd_last_state.s_ac_read_wd_lat .is_wysiwyg = "true";
defparam \ac_block:sig_addr_cmd_last_state.s_ac_read_wd_lat .power_up = "low";

arriaii_lcell_comb \Selector188~0 (
	.dataa(!\ac_block:sig_addr_cmd_state.s_ac_read_wd_lat~q ),
	.datab(!\sig_dimm_driving_dq~q ),
	.datac(!\ac_block:sig_addr_cmd_last_state.s_ac_read_wd_lat~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector188~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector188~0 .extended_lut = "off";
defparam \Selector188~0 .lut_mask = 64'h0404040404040404;
defparam \Selector188~0 .shared_arith = "off";

arriaii_lcell_comb \sig_addr_cmd_state~2 (
	.dataa(!\sig_ac_req.s_ac_read_poa_mtp~q ),
	.datab(!\sig_addr_cmd_state~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_addr_cmd_state~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_addr_cmd_state~2 .extended_lut = "off";
defparam \sig_addr_cmd_state~2 .lut_mask = 64'h1111111111111111;
defparam \sig_addr_cmd_state~2 .shared_arith = "off";

dffeas \ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp (
	.clk(clk),
	.d(\sig_addr_cmd_state~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.prn(vcc));
defparam \ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp .is_wysiwyg = "true";
defparam \ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp .power_up = "low";

arriaii_lcell_comb \ac_block:sig_count[7]~0 (
	.dataa(!\ac_block:sig_addr_cmd_state.s_ac_relax~q ),
	.datab(!\ac_block:sig_addr_cmd_last_state.s_ac_relax~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_block:sig_count[7]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_block:sig_count[7]~0 .extended_lut = "off";
defparam \ac_block:sig_count[7]~0 .lut_mask = 64'h4444444444444444;
defparam \ac_block:sig_count[7]~0 .shared_arith = "off";

arriaii_lcell_comb \Selector153~0 (
	.dataa(!\ac_block:sig_addr_cmd_last_state.s_ac_read_poa_mtp~q ),
	.datab(!\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector153~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector153~0 .extended_lut = "off";
defparam \Selector153~0 .lut_mask = 64'h1111111111111111;
defparam \Selector153~0 .shared_arith = "off";

arriaii_lcell_comb \sig_addr_cmd_state~3 (
	.dataa(!\sig_ac_req.s_ac_read_mtp~q ),
	.datab(!\sig_addr_cmd_state~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_addr_cmd_state~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_addr_cmd_state~3 .extended_lut = "off";
defparam \sig_addr_cmd_state~3 .lut_mask = 64'h1111111111111111;
defparam \sig_addr_cmd_state~3 .shared_arith = "off";

dffeas \ac_block:sig_addr_cmd_state.s_ac_read_mtp (
	.clk(clk),
	.d(\sig_addr_cmd_state~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.prn(vcc));
defparam \ac_block:sig_addr_cmd_state.s_ac_read_mtp .is_wysiwyg = "true";
defparam \ac_block:sig_addr_cmd_state.s_ac_read_mtp .power_up = "low";

dffeas \ac_block:sig_addr_cmd_last_state.s_ac_read_mtp (
	.clk(clk),
	.d(\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_block:sig_addr_cmd_last_state.s_ac_read_mtp~q ),
	.prn(vcc));
defparam \ac_block:sig_addr_cmd_last_state.s_ac_read_mtp .is_wysiwyg = "true";
defparam \ac_block:sig_addr_cmd_last_state.s_ac_read_mtp .power_up = "low";

dffeas \ac_block:sig_addr_cmd_last_state.s_ac_read_rdv (
	.clk(clk),
	.d(\ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_block:sig_addr_cmd_last_state.s_ac_read_rdv~q ),
	.prn(vcc));
defparam \ac_block:sig_addr_cmd_last_state.s_ac_read_rdv .is_wysiwyg = "true";
defparam \ac_block:sig_addr_cmd_last_state.s_ac_read_rdv .power_up = "low";

arriaii_lcell_comb \ac_block:sig_count[7]~1 (
	.dataa(!\Equal21~0_combout ),
	.datab(!\Selector153~0_combout ),
	.datac(!\ac_block:sig_addr_cmd_last_state.s_ac_read_mtp~q ),
	.datad(!\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.datae(!\ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ),
	.dataf(!\ac_block:sig_addr_cmd_last_state.s_ac_read_rdv~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_block:sig_count[7]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_block:sig_count[7]~1 .extended_lut = "off";
defparam \ac_block:sig_count[7]~1 .lut_mask = 64'hEE0A0000EE0AAAAA;
defparam \ac_block:sig_count[7]~1 .shared_arith = "off";

arriaii_lcell_comb \Selector182~0 (
	.dataa(!\Equal21~0_combout ),
	.datab(!\ac_block:sig_addr_cmd_last_state.s_ac_read_mtp~q ),
	.datac(!\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.datad(!\ac_block:sig_count[7]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector182~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector182~0 .extended_lut = "off";
defparam \Selector182~0 .lut_mask = 64'hF200F200F200F200;
defparam \Selector182~0 .shared_arith = "off";

arriaii_lcell_comb \Selector186~0 (
	.dataa(!\ac_block:sig_addr_cmd_last_state.s_ac_read_poa_mtp~q ),
	.datab(!\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.datac(!\ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ),
	.datad(!\ac_block:sig_addr_cmd_last_state.s_ac_read_rdv~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector186~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector186~0 .extended_lut = "off";
defparam \Selector186~0 .lut_mask = 64'h2F222F222F222F22;
defparam \Selector186~0 .shared_arith = "off";

arriaii_lcell_comb \Add24~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\ac_block:sig_count[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add24~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~13_sumout ),
	.cout(\Add24~14 ),
	.shareout());
defparam \Add24~13 .extended_lut = "off";
defparam \Add24~13 .lut_mask = 64'h00000000000000FF;
defparam \Add24~13 .shared_arith = "off";

arriaii_lcell_comb \Add24~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\ac_block:sig_count[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add24~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~17_sumout ),
	.cout(\Add24~18 ),
	.shareout());
defparam \Add24~17 .extended_lut = "off";
defparam \Add24~17 .lut_mask = 64'h00000000000000FF;
defparam \Add24~17 .shared_arith = "off";

dffeas \ac_block:sig_addr_cmd_last_state.s_ac_read_poa_mtp (
	.clk(clk),
	.d(\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_block:sig_addr_cmd_last_state.s_ac_read_poa_mtp~q ),
	.prn(vcc));
defparam \ac_block:sig_addr_cmd_last_state.s_ac_read_poa_mtp .is_wysiwyg = "true";
defparam \ac_block:sig_addr_cmd_last_state.s_ac_read_poa_mtp .power_up = "low";

arriaii_lcell_comb \Selector153~1 (
	.dataa(!\ac_block:sig_burst_count[0]~q ),
	.datab(!dgb_ac_access_gnt_r),
	.datac(!\ac_block:sig_addr_cmd_last_state.s_ac_read_poa_mtp~q ),
	.datad(!\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector153~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector153~1 .extended_lut = "off";
defparam \Selector153~1 .lut_mask = 64'h0002000200020002;
defparam \Selector153~1 .shared_arith = "off";

arriaii_lcell_comb \Selector183~0 (
	.dataa(!\ac_block:sig_burst_count[0]~q ),
	.datab(!\ac_block:sig_addr_cmd_last_state.s_ac_read_mtp~q ),
	.datac(!\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector183~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector183~0 .extended_lut = "off";
defparam \Selector183~0 .lut_mask = 64'h0202020202020202;
defparam \Selector183~0 .shared_arith = "off";

arriaii_lcell_comb \Selector183~1 (
	.dataa(!\Equal21~0_combout ),
	.datab(!\ac_block:sig_addr_cmd_state.s_ac_relax~q ),
	.datac(!\Selector153~1_combout ),
	.datad(!\Selector183~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector183~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector183~1 .extended_lut = "off";
defparam \Selector183~1 .lut_mask = 64'h2AAA2AAA2AAA2AAA;
defparam \Selector183~1 .shared_arith = "off";

arriaii_lcell_comb \Selector183~2 (
	.dataa(!\ac_block:sig_burst_count[0]~q ),
	.datab(!\ac_block:sig_addr_cmd_state.s_ac_read_wd_lat~q ),
	.datac(!dgb_ac_access_gnt_r),
	.datad(!\Selector153~0_combout ),
	.datae(!\ac_block:sig_addr_cmd_state.s_ac_idle~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector183~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector183~2 .extended_lut = "off";
defparam \Selector183~2 .lut_mask = 64'h0000CC080000CC08;
defparam \Selector183~2 .shared_arith = "off";

arriaii_lcell_comb \Selector183~3 (
	.dataa(!\ac_block:sig_burst_count[0]~q ),
	.datab(!\ac_block:sig_addr_cmd_last_state.s_ac_read_mtp~q ),
	.datac(!\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.datad(!\ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ),
	.datae(!\Selector183~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector183~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector183~3 .extended_lut = "off";
defparam \Selector183~3 .lut_mask = 64'h0000FEAA0000FEAA;
defparam \Selector183~3 .shared_arith = "off";

arriaii_lcell_comb \Selector183~4 (
	.dataa(!\ac_block:sig_count[4]~q ),
	.datab(!\ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ),
	.datac(!\ac_block:sig_addr_cmd_last_state.s_ac_read_rdv~q ),
	.datad(!\ac_block:sig_count[7]~0_combout ),
	.datae(!\Selector183~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector183~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector183~4 .extended_lut = "off";
defparam \Selector183~4 .lut_mask = 64'h8A00CF008A00CF00;
defparam \Selector183~4 .shared_arith = "off";

arriaii_lcell_comb \Selector183~5 (
	.dataa(!\ac_block:sig_burst_count[0]~q ),
	.datab(!\ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ),
	.datac(!\Add24~17_sumout ),
	.datad(!\Selector183~1_combout ),
	.datae(!\Selector183~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector183~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector183~5 .extended_lut = "off";
defparam \Selector183~5 .lut_mask = 64'hFFFF020FFFFF020F;
defparam \Selector183~5 .shared_arith = "off";

dffeas \ac_block:sig_count[4] (
	.clk(clk),
	.d(\Selector183~5_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_block:sig_count[4]~q ),
	.prn(vcc));
defparam \ac_block:sig_count[4] .is_wysiwyg = "true";
defparam \ac_block:sig_count[4] .power_up = "low";

arriaii_lcell_comb \Add24~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\ac_block:sig_count[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add24~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~21_sumout ),
	.cout(\Add24~22 ),
	.shareout());
defparam \Add24~21 .extended_lut = "off";
defparam \Add24~21 .lut_mask = 64'h00000000000000FF;
defparam \Add24~21 .shared_arith = "off";

arriaii_lcell_comb \Selector182~1 (
	.dataa(!\ac_block:sig_count[5]~0_combout ),
	.datab(!\Selector182~0_combout ),
	.datac(!\Selector186~0_combout ),
	.datad(!\Add24~21_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector182~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector182~1 .extended_lut = "off";
defparam \Selector182~1 .lut_mask = 64'h1F3F1F3F1F3F1F3F;
defparam \Selector182~1 .shared_arith = "off";

arriaii_lcell_comb \ac_block:sig_count[5]~3 (
	.dataa(!\ac_block:sig_burst_count[0]~q ),
	.datab(!dgb_ac_access_gnt_r),
	.datac(!\ac_block:sig_addr_cmd_last_state.s_ac_read_poa_mtp~q ),
	.datad(!\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_block:sig_count[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_block:sig_count[5]~3 .extended_lut = "off";
defparam \ac_block:sig_count[5]~3 .lut_mask = 64'h00F200F200F200F2;
defparam \ac_block:sig_count[5]~3 .shared_arith = "off";

arriaii_lcell_comb \ac_block:sig_count[5]~4 (
	.dataa(!\ac_block:sig_count[1]~q ),
	.datab(!\ac_block:sig_count[5]~q ),
	.datac(!\ac_block:sig_count[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_block:sig_count[5]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_block:sig_count[5]~4 .extended_lut = "off";
defparam \ac_block:sig_count[5]~4 .lut_mask = 64'h8080808080808080;
defparam \ac_block:sig_count[5]~4 .shared_arith = "off";

arriaii_lcell_comb \ac_block:sig_count[5]~5 (
	.dataa(!\ac_block:sig_burst_count[0]~q ),
	.datab(!\ac_block:sig_addr_cmd_last_state.s_ac_read_mtp~q ),
	.datac(!\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.datad(!\ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ),
	.datae(!\ac_block:sig_addr_cmd_last_state.s_ac_read_rdv~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_block:sig_count[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_block:sig_count[5]~5 .extended_lut = "off";
defparam \ac_block:sig_count[5]~5 .lut_mask = 64'hF100F151F100F151;
defparam \ac_block:sig_count[5]~5 .shared_arith = "off";

arriaii_lcell_comb \ac_block:sig_count[5]~0 (
	.dataa(!\Equal21~0_combout ),
	.datab(!\Selector153~0_combout ),
	.datac(!\ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ),
	.datad(!\ac_block:sig_addr_cmd_last_state.s_ac_read_rdv~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_block:sig_count[5]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_block:sig_count[5]~0 .extended_lut = "off";
defparam \ac_block:sig_count[5]~0 .lut_mask = 64'h1115111511151115;
defparam \ac_block:sig_count[5]~0 .shared_arith = "off";

arriaii_lcell_comb \Selector187~0 (
	.dataa(!\Add24~1_sumout ),
	.datab(!\ac_block:sig_count[5]~0_combout ),
	.datac(!\Selector182~0_combout ),
	.datad(!\Selector186~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector187~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector187~0 .extended_lut = "off";
defparam \Selector187~0 .lut_mask = 64'hF400F400F400F400;
defparam \Selector187~0 .shared_arith = "off";

dffeas \ac_block:sig_count[0] (
	.clk(clk),
	.d(\Selector187~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ac_block:sig_count[5]~1_combout ),
	.q(\ac_block:sig_count[0]~q ),
	.prn(vcc));
defparam \ac_block:sig_count[0] .is_wysiwyg = "true";
defparam \ac_block:sig_count[0] .power_up = "low";

arriaii_lcell_comb \ac_block:sig_count[7]~4 (
	.dataa(!\ac_block:sig_addr_cmd_last_state.s_ac_relax~q ),
	.datab(!\ac_block:sig_count[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_block:sig_count[7]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_block:sig_count[7]~4 .extended_lut = "off";
defparam \ac_block:sig_count[7]~4 .lut_mask = 64'h4444444444444444;
defparam \ac_block:sig_count[7]~4 .shared_arith = "off";

arriaii_lcell_comb \ac_block:sig_count[5]~1 (
	.dataa(!\ac_block:sig_addr_cmd_state.s_ac_relax~q ),
	.datab(!\Selector189~0_combout ),
	.datac(!\ac_block:sig_count[5]~3_combout ),
	.datad(!\ac_block:sig_count[5]~4_combout ),
	.datae(!\ac_block:sig_count[5]~5_combout ),
	.dataf(!\ac_block:sig_count[7]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_block:sig_count[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_block:sig_count[5]~1 .extended_lut = "off";
defparam \ac_block:sig_count[5]~1 .lut_mask = 64'hFFFF5F5FFFFF5F4F;
defparam \ac_block:sig_count[5]~1 .shared_arith = "off";

dffeas \ac_block:sig_count[5] (
	.clk(clk),
	.d(\Selector182~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ac_block:sig_count[5]~1_combout ),
	.q(\ac_block:sig_count[5]~q ),
	.prn(vcc));
defparam \ac_block:sig_count[5] .is_wysiwyg = "true";
defparam \ac_block:sig_count[5] .power_up = "low";

arriaii_lcell_comb \Equal21~1 (
	.dataa(!\Selector189~0_combout ),
	.datab(!\ac_block:sig_count[1]~q ),
	.datac(!\ac_block:sig_count[5]~q ),
	.datad(!\ac_block:sig_count[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal21~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal21~1 .extended_lut = "off";
defparam \Equal21~1 .lut_mask = 64'h4000400040004000;
defparam \Equal21~1 .shared_arith = "off";

arriaii_lcell_comb \ac_block:sig_count[5]~2 (
	.dataa(!\ac_block:sig_count[0]~q ),
	.datab(!\Equal21~1_combout ),
	.datac(!\ac_block:sig_addr_cmd_last_state.s_ac_read_mtp~q ),
	.datad(!\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_block:sig_count[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_block:sig_count[5]~2 .extended_lut = "off";
defparam \ac_block:sig_count[5]~2 .lut_mask = 64'h00F200F200F200F2;
defparam \ac_block:sig_count[5]~2 .shared_arith = "off";

arriaii_lcell_comb \Add24~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\ac_block:sig_count[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add24~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~5_sumout ),
	.cout(\Add24~6 ),
	.shareout());
defparam \Add24~5 .extended_lut = "off";
defparam \Add24~5 .lut_mask = 64'h00000000000000FF;
defparam \Add24~5 .shared_arith = "off";

arriaii_lcell_comb \Selector186~1 (
	.dataa(!\ac_block:sig_count[5]~0_combout ),
	.datab(!\ac_block:sig_count[7]~0_combout ),
	.datac(!\ac_block:sig_count[5]~2_combout ),
	.datad(!\Selector186~0_combout ),
	.datae(!\Add24~5_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector186~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector186~1 .extended_lut = "off";
defparam \Selector186~1 .lut_mask = 64'h70FFF0FF70FFF0FF;
defparam \Selector186~1 .shared_arith = "off";

dffeas \ac_block:sig_count[1] (
	.clk(clk),
	.d(\Selector186~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ac_block:sig_count[5]~1_combout ),
	.q(\ac_block:sig_count[1]~q ),
	.prn(vcc));
defparam \ac_block:sig_count[1] .is_wysiwyg = "true";
defparam \ac_block:sig_count[1] .power_up = "low";

arriaii_lcell_comb \Add24~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\ac_block:sig_count[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add24~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~9_sumout ),
	.cout(\Add24~10 ),
	.shareout());
defparam \Add24~9 .extended_lut = "off";
defparam \Add24~9 .lut_mask = 64'h00000000000000FF;
defparam \Add24~9 .shared_arith = "off";

arriaii_lcell_comb \Selector185~0 (
	.dataa(!\ac_block:sig_addr_cmd_last_state.s_ac_read_poa_mtp~q ),
	.datab(!\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.datac(!\ac_block:sig_count[7]~0_combout ),
	.datad(!\Add24~9_sumout ),
	.datae(!\ac_block:sig_count[7]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector185~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector185~0 .extended_lut = "off";
defparam \Selector185~0 .lut_mask = 64'h0D0D0DDD0D0D0DDD;
defparam \Selector185~0 .shared_arith = "off";

arriaii_lcell_comb \ac_block:sig_count[7]~3 (
	.dataa(!\ac_block:sig_burst_count[0]~q ),
	.datab(!\ac_block:sig_addr_cmd_last_state.s_ac_read_mtp~q ),
	.datac(!\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.datad(!\ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ),
	.datae(!\ac_block:sig_addr_cmd_last_state.s_ac_read_rdv~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_block:sig_count[7]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_block:sig_count[7]~3 .extended_lut = "off";
defparam \ac_block:sig_count[7]~3 .lut_mask = 64'hF100F155F100F155;
defparam \ac_block:sig_count[7]~3 .shared_arith = "off";

arriaii_lcell_comb \ac_block:sig_count[7]~2 (
	.dataa(!\ac_block:sig_addr_cmd_state.s_ac_relax~q ),
	.datab(!\Selector189~0_combout ),
	.datac(!\ac_block:sig_count[5]~3_combout ),
	.datad(!\ac_block:sig_count[5]~4_combout ),
	.datae(!\ac_block:sig_count[7]~3_combout ),
	.dataf(!\ac_block:sig_count[7]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_block:sig_count[7]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_block:sig_count[7]~2 .extended_lut = "off";
defparam \ac_block:sig_count[7]~2 .lut_mask = 64'hFFFF5F5FFFFF5F4F;
defparam \ac_block:sig_count[7]~2 .shared_arith = "off";

dffeas \ac_block:sig_count[2] (
	.clk(clk),
	.d(\Selector185~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ac_block:sig_count[7]~2_combout ),
	.q(\ac_block:sig_count[2]~q ),
	.prn(vcc));
defparam \ac_block:sig_count[2] .is_wysiwyg = "true";
defparam \ac_block:sig_count[2] .power_up = "low";

arriaii_lcell_comb \Selector184~0 (
	.dataa(!\ac_block:sig_addr_cmd_last_state.s_ac_read_poa_mtp~q ),
	.datab(!\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.datac(!\ac_block:sig_count[7]~0_combout ),
	.datad(!\ac_block:sig_count[7]~1_combout ),
	.datae(!\Add24~13_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector184~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector184~0 .extended_lut = "off";
defparam \Selector184~0 .lut_mask = 64'h0D0D0DDD0D0D0DDD;
defparam \Selector184~0 .shared_arith = "off";

dffeas \ac_block:sig_count[3] (
	.clk(clk),
	.d(\Selector184~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ac_block:sig_count[7]~2_combout ),
	.q(\ac_block:sig_count[3]~q ),
	.prn(vcc));
defparam \ac_block:sig_count[3] .is_wysiwyg = "true";
defparam \ac_block:sig_count[3] .power_up = "low";

arriaii_lcell_comb \Add24~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\ac_block:sig_count[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add24~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~25_sumout ),
	.cout(\Add24~26 ),
	.shareout());
defparam \Add24~25 .extended_lut = "off";
defparam \Add24~25 .lut_mask = 64'h00000000000000FF;
defparam \Add24~25 .shared_arith = "off";

arriaii_lcell_comb \Selector181~0 (
	.dataa(!\ac_block:sig_addr_cmd_last_state.s_ac_read_poa_mtp~q ),
	.datab(!\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.datac(!\ac_block:sig_count[7]~0_combout ),
	.datad(!\ac_block:sig_count[7]~1_combout ),
	.datae(!\Add24~25_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector181~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector181~0 .extended_lut = "off";
defparam \Selector181~0 .lut_mask = 64'h000000D0000000D0;
defparam \Selector181~0 .shared_arith = "off";

dffeas \ac_block:sig_count[6] (
	.clk(clk),
	.d(\Selector181~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ac_block:sig_count[7]~2_combout ),
	.q(\ac_block:sig_count[6]~q ),
	.prn(vcc));
defparam \ac_block:sig_count[6] .is_wysiwyg = "true";
defparam \ac_block:sig_count[6] .power_up = "low";

arriaii_lcell_comb \Add24~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\ac_block:sig_count[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add24~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add24~29_sumout ),
	.cout(),
	.shareout());
defparam \Add24~29 .extended_lut = "off";
defparam \Add24~29 .lut_mask = 64'h00000000000000FF;
defparam \Add24~29 .shared_arith = "off";

arriaii_lcell_comb \Selector180~0 (
	.dataa(!\ac_block:sig_addr_cmd_last_state.s_ac_read_poa_mtp~q ),
	.datab(!\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.datac(!\ac_block:sig_count[7]~0_combout ),
	.datad(!\ac_block:sig_count[7]~1_combout ),
	.datae(!\Add24~29_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector180~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector180~0 .extended_lut = "off";
defparam \Selector180~0 .lut_mask = 64'h000000D0000000D0;
defparam \Selector180~0 .shared_arith = "off";

dffeas \ac_block:sig_count[7] (
	.clk(clk),
	.d(\Selector180~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ac_block:sig_count[7]~2_combout ),
	.q(\ac_block:sig_count[7]~q ),
	.prn(vcc));
defparam \ac_block:sig_count[7] .is_wysiwyg = "true";
defparam \ac_block:sig_count[7] .power_up = "low";

arriaii_lcell_comb \Selector189~0 (
	.dataa(!\ac_block:sig_count[2]~q ),
	.datab(!\ac_block:sig_count[3]~q ),
	.datac(!\ac_block:sig_count[7]~q ),
	.datad(!\ac_block:sig_count[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector189~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector189~0 .extended_lut = "off";
defparam \Selector189~0 .lut_mask = 64'h8000800080008000;
defparam \Selector189~0 .shared_arith = "off";

arriaii_lcell_comb \Equal21~0 (
	.dataa(!\ac_block:sig_count[0]~q ),
	.datab(!\Selector189~0_combout ),
	.datac(!\ac_block:sig_count[1]~q ),
	.datad(!\ac_block:sig_count[5]~q ),
	.datae(!\ac_block:sig_count[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal21~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal21~0 .extended_lut = "off";
defparam \Equal21~0 .lut_mask = 64'h2000000020000000;
defparam \Equal21~0 .shared_arith = "off";

arriaii_lcell_comb \sig_doing_rd_count~0 (
	.dataa(!\ac_block:sig_burst_count[0]~q ),
	.datab(!\Equal21~0_combout ),
	.datac(!dgb_ac_access_gnt_r),
	.datad(!\ac_block:sig_addr_cmd_last_state.s_ac_read_poa_mtp~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_doing_rd_count~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_doing_rd_count~0 .extended_lut = "off";
defparam \sig_doing_rd_count~0 .lut_mask = 64'h0002000200020002;
defparam \sig_doing_rd_count~0 .shared_arith = "off";

dffeas \ac_block:sig_doing_rd_count (
	.clk(clk),
	.d(\sig_doing_rd_count~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\ac_block:sig_doing_rd_count~q ),
	.prn(vcc));
defparam \ac_block:sig_doing_rd_count .is_wysiwyg = "true";
defparam \ac_block:sig_doing_rd_count .power_up = "low";

arriaii_lcell_comb \Selector188~1 (
	.dataa(!\ac_block:sig_addr_cmd_state.s_ac_read_wd_lat~q ),
	.datab(!\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.datac(!\ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector188~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector188~1 .extended_lut = "off";
defparam \Selector188~1 .lut_mask = 64'h8080808080808080;
defparam \Selector188~1 .shared_arith = "off";

arriaii_lcell_comb \dimm_driving_dq_proc~0 (
	.dataa(!\ac_block:sig_addr_cmd_state.s_ac_idle~q ),
	.datab(!\ac_block:sig_addr_cmd_state.s_ac_relax~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dimm_driving_dq_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dimm_driving_dq_proc~0 .extended_lut = "off";
defparam \dimm_driving_dq_proc~0 .lut_mask = 64'h4444444444444444;
defparam \dimm_driving_dq_proc~0 .shared_arith = "off";

arriaii_lcell_comb \Selector188~2 (
	.dataa(!\ac_block:sig_addr_cmd_last_state.s_ac_read_mtp~q ),
	.datab(!\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.datac(!\ac_block:sig_doing_rd_count~q ),
	.datad(!\Selector188~1_combout ),
	.datae(!\dimm_driving_dq_proc~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector188~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector188~2 .extended_lut = "off";
defparam \Selector188~2 .lut_mask = 64'hE0E0E0ECE0E0E0EC;
defparam \Selector188~2 .shared_arith = "off";

arriaii_lcell_comb \Selector188~3 (
	.dataa(!\ac_block:sig_burst_count[0]~q ),
	.datab(!\Selector188~0_combout ),
	.datac(!\Equal21~0_combout ),
	.datad(!dgb_ac_access_gnt_r),
	.datae(!\Selector153~0_combout ),
	.dataf(!\Selector188~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector188~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector188~3 .extended_lut = "off";
defparam \Selector188~3 .lut_mask = 64'hFFFFFFFF2222222A;
defparam \Selector188~3 .shared_arith = "off";

arriaii_lcell_comb \seq_rdata_valid_lat_dec~0 (
	.dataa(!\sig_dimm_driving_dq~q ),
	.datab(!rdata_valid[0]),
	.datac(!seq_rdata_valid_1),
	.datad(!\v_aligned~0_combout ),
	.datae(!\sig_dgrb_state.s_rdata_valid_align~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_rdata_valid_lat_dec~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_rdata_valid_lat_dec~0 .extended_lut = "off";
defparam \seq_rdata_valid_lat_dec~0 .lut_mask = 64'h00002A0000002A00;
defparam \seq_rdata_valid_lat_dec~0 .shared_arith = "off";

arriaii_lcell_comb \Selector189~1 (
	.dataa(!\ac_block:sig_burst_count[0]~q ),
	.datab(!\ac_block:sig_count[0]~q ),
	.datac(!\ac_block:sig_count[1]~q ),
	.datad(!\ac_block:sig_count[5]~q ),
	.datae(!\ac_block:sig_count[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector189~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector189~1 .extended_lut = "off";
defparam \Selector189~1 .lut_mask = 64'h0000000400000004;
defparam \Selector189~1 .shared_arith = "off";

arriaii_lcell_comb \Selector189~2 (
	.dataa(!\Selector189~0_combout ),
	.datab(!\ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ),
	.datac(!\Selector188~3_combout ),
	.datad(!\Selector189~1_combout ),
	.datae(!\ac_block:sig_addr_cmd_last_state.s_ac_read_rdv~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector189~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector189~2 .extended_lut = "off";
defparam \Selector189~2 .lut_mask = 64'h0F0F0F1F0F0F0F1F;
defparam \Selector189~2 .shared_arith = "off";

arriaii_lcell_comb \dgrb_ctrl_ac_nt_good~0 (
	.dataa(!q_b_12),
	.datab(!q_b_76),
	.datac(!q_b_13),
	.datad(!q_b_77),
	.datae(!q_b_14),
	.dataf(!q_b_78),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dgrb_ctrl_ac_nt_good~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dgrb_ctrl_ac_nt_good~0 .extended_lut = "off";
defparam \dgrb_ctrl_ac_nt_good~0 .lut_mask = 64'h9009000000009009;
defparam \dgrb_ctrl_ac_nt_good~0 .shared_arith = "off";

arriaii_lcell_comb \dgrb_ctrl_ac_nt_good~1 (
	.dataa(!q_b_9),
	.datab(!q_b_73),
	.datac(!q_b_10),
	.datad(!q_b_74),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dgrb_ctrl_ac_nt_good~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dgrb_ctrl_ac_nt_good~1 .extended_lut = "off";
defparam \dgrb_ctrl_ac_nt_good~1 .lut_mask = 64'h9009900990099009;
defparam \dgrb_ctrl_ac_nt_good~1 .shared_arith = "off";

arriaii_lcell_comb \dgrb_ctrl_ac_nt_good~2 (
	.dataa(!q_b_6),
	.datab(!q_b_70),
	.datac(!q_b_7),
	.datad(!q_b_71),
	.datae(!q_b_8),
	.dataf(!q_b_72),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dgrb_ctrl_ac_nt_good~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dgrb_ctrl_ac_nt_good~2 .extended_lut = "off";
defparam \dgrb_ctrl_ac_nt_good~2 .lut_mask = 64'h9009000000009009;
defparam \dgrb_ctrl_ac_nt_good~2 .shared_arith = "off";

arriaii_lcell_comb \dgrb_ctrl_ac_nt_good~3 (
	.dataa(!q_b_0),
	.datab(!q_b_64),
	.datac(!q_b_1),
	.datad(!q_b_65),
	.datae(!q_b_2),
	.dataf(!q_b_66),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dgrb_ctrl_ac_nt_good~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dgrb_ctrl_ac_nt_good~3 .extended_lut = "off";
defparam \dgrb_ctrl_ac_nt_good~3 .lut_mask = 64'h9009000000009009;
defparam \dgrb_ctrl_ac_nt_good~3 .shared_arith = "off";

arriaii_lcell_comb \dgrb_ctrl_ac_nt_good~4 (
	.dataa(!q_b_3),
	.datab(!q_b_67),
	.datac(!q_b_4),
	.datad(!q_b_68),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dgrb_ctrl_ac_nt_good~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dgrb_ctrl_ac_nt_good~4 .extended_lut = "off";
defparam \dgrb_ctrl_ac_nt_good~4 .lut_mask = 64'h9009900990099009;
defparam \dgrb_ctrl_ac_nt_good~4 .shared_arith = "off";

arriaii_lcell_comb \dgrb_ctrl_ac_nt_good~5 (
	.dataa(!q_b_5),
	.datab(!q_b_69),
	.datac(!\dgrb_ctrl_ac_nt_good~2_combout ),
	.datad(!\dgrb_ctrl_ac_nt_good~3_combout ),
	.datae(!\dgrb_ctrl_ac_nt_good~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dgrb_ctrl_ac_nt_good~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dgrb_ctrl_ac_nt_good~5 .extended_lut = "off";
defparam \dgrb_ctrl_ac_nt_good~5 .lut_mask = 64'h0000000900000009;
defparam \dgrb_ctrl_ac_nt_good~5 .shared_arith = "off";

arriaii_lcell_comb \dgrb_ctrl_ac_nt_good~6 (
	.dataa(!q_b_11),
	.datab(!q_b_75),
	.datac(!\dgrb_ctrl_ac_nt_good~0_combout ),
	.datad(!\dgrb_ctrl_ac_nt_good~1_combout ),
	.datae(!\dgrb_ctrl_ac_nt_good~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dgrb_ctrl_ac_nt_good~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dgrb_ctrl_ac_nt_good~6 .extended_lut = "off";
defparam \dgrb_ctrl_ac_nt_good~6 .lut_mask = 64'h0000000900000009;
defparam \dgrb_ctrl_ac_nt_good~6 .shared_arith = "off";

arriaii_lcell_comb \Selector32~0 (
	.dataa(!\sig_dimm_driving_dq~q ),
	.datab(!\sig_dgrb_last_state.s_adv_wd_lat~q ),
	.datac(!\sig_dgrb_state.s_adv_wd_lat~q ),
	.datad(!rdata_valid[0]),
	.datae(!seq_rdata_valid_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector32~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector32~0 .extended_lut = "off";
defparam \Selector32~0 .lut_mask = 64'h0002020200020202;
defparam \Selector32~0 .shared_arith = "off";

arriaii_lcell_comb \dgrb_ctrl_ac_nt_good~7 (
	.dataa(!q_b_15),
	.datab(!q_b_79),
	.datac(!dgrb_ctrl_ac_nt_good1),
	.datad(!\dgrb_ctrl_ac_nt_good~6_combout ),
	.datae(!\Selector32~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dgrb_ctrl_ac_nt_good~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dgrb_ctrl_ac_nt_good~7 .extended_lut = "off";
defparam \dgrb_ctrl_ac_nt_good~7 .lut_mask = 64'h0F0FFF660F0FFF66;
defparam \dgrb_ctrl_ac_nt_good~7 .shared_arith = "off";

arriaii_lcell_comb \pll_reconf_mux~0 (
	.dataa(!\sig_dgrb_state.s_seek_cdvw~q ),
	.datab(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datac(!\sig_dgrb_state.s_test_phases~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pll_reconf_mux~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pll_reconf_mux~0 .extended_lut = "off";
defparam \pll_reconf_mux~0 .lut_mask = 64'h8080808080808080;
defparam \pll_reconf_mux~0 .shared_arith = "off";

arriaii_lcell_comb \sig_rsc_pll_inc_dec_n~0 (
	.dataa(!\rsc_block:sig_rewind_direction~q ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_rewind_phase~q ),
	.datac(!\Equal13~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_rsc_pll_inc_dec_n~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_rsc_pll_inc_dec_n~0 .extended_lut = "off";
defparam \sig_rsc_pll_inc_dec_n~0 .lut_mask = 64'h0202020202020202;
defparam \sig_rsc_pll_inc_dec_n~0 .shared_arith = "off";

dffeas sig_rsc_pll_inc_dec_n(
	.clk(clk),
	.d(\sig_rsc_pll_inc_dec_n~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_rsc_pll_inc_dec_n~q ),
	.prn(vcc));
defparam sig_rsc_pll_inc_dec_n.is_wysiwyg = "true";
defparam sig_rsc_pll_inc_dec_n.power_up = "low";

arriaii_lcell_comb \sig_trk_pll_inc_dec_n~2 (
	.dataa(!\sig_trk_pll_inc_dec_n~q ),
	.datab(!\trk_block:sig_trk_last_state.s_trk_adjust_resync~q ),
	.datac(!\trk_block:sig_req_rsc_shift[7]~q ),
	.datad(!\LessThan11~1_combout ),
	.datae(!\sig_trk_pll_inc_dec_n~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_trk_pll_inc_dec_n~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_trk_pll_inc_dec_n~2 .extended_lut = "off";
defparam \sig_trk_pll_inc_dec_n~2 .lut_mask = 64'h0000111D0000111D;
defparam \sig_trk_pll_inc_dec_n~2 .shared_arith = "off";

dffeas sig_trk_pll_inc_dec_n(
	.clk(clk),
	.d(\sig_trk_pll_inc_dec_n~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_trk_pll_inc_dec_n~q ),
	.prn(vcc));
defparam sig_trk_pll_inc_dec_n.is_wysiwyg = "true";
defparam sig_trk_pll_inc_dec_n.power_up = "low";

arriaii_lcell_comb \seq_pll_inc_dec_n~0 (
	.dataa(!\pll_reconf_mux~0_combout ),
	.datab(!\sig_rsc_pll_inc_dec_n~q ),
	.datac(!\sig_trk_pll_inc_dec_n~q ),
	.datad(!\sig_dgrb_state.s_track~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_pll_inc_dec_n~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_pll_inc_dec_n~0 .extended_lut = "off";
defparam \seq_pll_inc_dec_n~0 .lut_mask = 64'h88D888D888D888D8;
defparam \seq_pll_inc_dec_n~0 .shared_arith = "off";

dffeas sig_phs_shft_busy_1t(
	.clk(clk),
	.d(\sig_phs_shft_busy~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_phs_shft_busy_1t~q ),
	.prn(vcc));
defparam sig_phs_shft_busy_1t.is_wysiwyg = "true";
defparam sig_phs_shft_busy_1t.power_up = "low";

arriaii_lcell_comb \Selector61~0 (
	.dataa(!\rsc_block:sig_rsc_state.s_rsc_rewind_phase~q ),
	.datab(!\Equal13~0_combout ),
	.datac(!\sig_phs_shft_busy~q ),
	.datad(!\sig_phs_shft_busy_1t~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector61~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector61~0 .extended_lut = "off";
defparam \Selector61~0 .lut_mask = 64'h1000100010001000;
defparam \Selector61~0 .shared_arith = "off";

arriaii_lcell_comb \Selector61~1 (
	.dataa(!\sig_phs_shft_start~q ),
	.datab(!\rsc_block:sig_rsc_state.s_rsc_next_phase~q ),
	.datac(!\Equal14~1_combout ),
	.datad(!\Selector71~0_combout ),
	.datae(!\Selector61~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector61~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector61~1 .extended_lut = "off";
defparam \Selector61~1 .lut_mask = 64'h22A2FFFF22A2FFFF;
defparam \Selector61~1 .shared_arith = "off";

dffeas sig_rsc_pll_start_reconfig(
	.clk(clk),
	.d(\Selector61~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_rsc_pll_start_reconfig~q ),
	.prn(vcc));
defparam sig_rsc_pll_start_reconfig.is_wysiwyg = "true";
defparam sig_rsc_pll_start_reconfig.power_up = "low";

arriaii_lcell_comb \sig_phs_shft_start~0 (
	.dataa(!\sig_phs_shft_busy~q ),
	.datab(!\phs_shft_busy_reg:phs_shft_busy_2r~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_phs_shft_start~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_phs_shft_start~0 .extended_lut = "off";
defparam \sig_phs_shft_start~0 .lut_mask = 64'h7777777777777777;
defparam \sig_phs_shft_start~0 .shared_arith = "off";

dffeas sig_phs_shft_start(
	.clk(clk),
	.d(\sig_phs_shft_start~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_phs_shft_start~q ),
	.prn(vcc));
defparam sig_phs_shft_start.is_wysiwyg = "true";
defparam sig_phs_shft_start.power_up = "low";

arriaii_lcell_comb \sig_trk_state~19 (
	.dataa(!\trk_block:sig_trk_state.s_trk_next_phase~q ),
	.datab(!\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.datac(!\shift_in_mmc_seq_value~0_combout ),
	.datad(!\Equal17~1_combout ),
	.datae(!\sig_trk_state~16_combout ),
	.dataf(!\sig_trk_state~18_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_trk_state~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_trk_state~19 .extended_lut = "off";
defparam \sig_trk_state~19 .lut_mask = 64'h0000000003005755;
defparam \sig_trk_state~19 .shared_arith = "off";

dffeas \trk_block:sig_trk_state.s_trk_next_phase (
	.clk(clk),
	.d(\sig_trk_state~19_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_trk_state.s_trk_next_phase~q ),
	.prn(vcc));
defparam \trk_block:sig_trk_state.s_trk_next_phase .is_wysiwyg = "true";
defparam \trk_block:sig_trk_state.s_trk_next_phase .power_up = "low";

arriaii_lcell_comb \Selector127~0 (
	.dataa(!\trk_block:sig_trk_last_state.s_trk_adjust_resync~q ),
	.datab(!\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.datac(!\sig_phs_shft_start~q ),
	.datad(!\trk_block:sig_trk_state.s_trk_next_phase~q ),
	.datae(!\sig_trk_state~11_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector127~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector127~0 .extended_lut = "off";
defparam \Selector127~0 .lut_mask = 64'h30F010F030F010F0;
defparam \Selector127~0 .shared_arith = "off";

dffeas sig_trk_pll_start_reconfig(
	.clk(clk),
	.d(\Selector127~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_track~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_trk_pll_start_reconfig~q ),
	.prn(vcc));
defparam sig_trk_pll_start_reconfig.is_wysiwyg = "true";
defparam sig_trk_pll_start_reconfig.power_up = "low";

arriaii_lcell_comb \seq_pll_start_reconfig~0 (
	.dataa(!\pll_reconf_mux~0_combout ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\sig_rsc_pll_start_reconfig~q ),
	.datad(!\sig_trk_pll_start_reconfig~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_pll_start_reconfig~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_pll_start_reconfig~0 .extended_lut = "off";
defparam \seq_pll_start_reconfig~0 .lut_mask = 64'h0A1B0A1B0A1B0A1B;
defparam \seq_pll_start_reconfig~0 .shared_arith = "off";

dffeas \sig_dgrb_last_state.s_release_admin (
	.clk(clk),
	.d(\sig_dgrb_state.s_release_admin~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgrb_last_state.s_release_admin~q ),
	.prn(vcc));
defparam \sig_dgrb_last_state.s_release_admin .is_wysiwyg = "true";
defparam \sig_dgrb_last_state.s_release_admin .power_up = "low";

arriaii_lcell_comb \ac_handshake_proc~2 (
	.dataa(!\sig_dgrb_last_state.s_release_admin~q ),
	.datab(!\sig_dgrb_state.s_idle~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_handshake_proc~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_handshake_proc~2 .extended_lut = "off";
defparam \ac_handshake_proc~2 .lut_mask = 64'h4444444444444444;
defparam \ac_handshake_proc~2 .shared_arith = "off";

arriaii_lcell_comb \sig_rsc_result[0]~0 (
	.dataa(!\sig_dgrb_state.s_read_mtp~q ),
	.datab(!\sig_cdvw_state.status.calculating~q ),
	.datac(!\rsc_block:sig_rsc_state.s_rsc_cdvw_wait~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_rsc_result[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_rsc_result[0]~0 .extended_lut = "off";
defparam \sig_rsc_result[0]~0 .lut_mask = 64'h0808080808080808;
defparam \sig_rsc_result[0]~0 .shared_arith = "off";

arriaii_lcell_comb \sig_rsc_err~0 (
	.dataa(!\sig_rsc_err~q ),
	.datab(!\sig_cdvw_state.status.valid_result~q ),
	.datac(!\sig_rsc_result[0]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_rsc_err~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_rsc_err~0 .extended_lut = "off";
defparam \sig_rsc_err~0 .lut_mask = 64'h5D5D5D5D5D5D5D5D;
defparam \sig_rsc_err~0 .shared_arith = "off";

dffeas sig_rsc_err(
	.clk(clk),
	.d(\sig_rsc_err~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_rsc_err~q ),
	.prn(vcc));
defparam sig_rsc_err.is_wysiwyg = "true";
defparam sig_rsc_err.power_up = "low";

arriaii_lcell_comb \Add20~1 (
	.dataa(!\trk_block:sig_rsc_drift[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(!\trk_block:sig_rsc_drift[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add20~1_sumout ),
	.cout(\Add20~2 ),
	.shareout());
defparam \Add20~1 .extended_lut = "off";
defparam \Add20~1 .lut_mask = 64'h0000AA550000AAAA;
defparam \Add20~1 .shared_arith = "off";

arriaii_lcell_comb \Add20~5 (
	.dataa(!\trk_block:sig_rsc_drift[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_rsc_drift[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add20~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add20~5_sumout ),
	.cout(\Add20~6 ),
	.shareout());
defparam \Add20~5 .extended_lut = "off";
defparam \Add20~5 .lut_mask = 64'h0000FFFF0000AA55;
defparam \Add20~5 .shared_arith = "off";

arriaii_lcell_comb \Add20~9 (
	.dataa(!\trk_block:sig_rsc_drift[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_rsc_drift[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add20~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add20~9_sumout ),
	.cout(\Add20~10 ),
	.shareout());
defparam \Add20~9 .extended_lut = "off";
defparam \Add20~9 .lut_mask = 64'h0000FFFF0000AA55;
defparam \Add20~9 .shared_arith = "off";

arriaii_lcell_comb \Add20~13 (
	.dataa(!\trk_block:sig_rsc_drift[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_rsc_drift[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add20~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add20~13_sumout ),
	.cout(\Add20~14 ),
	.shareout());
defparam \Add20~13 .extended_lut = "off";
defparam \Add20~13 .lut_mask = 64'h0000FFFF0000AA55;
defparam \Add20~13 .shared_arith = "off";

arriaii_lcell_comb \Add20~17 (
	.dataa(!\trk_block:sig_rsc_drift[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_rsc_drift[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add20~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add20~17_sumout ),
	.cout(\Add20~18 ),
	.shareout());
defparam \Add20~17 .extended_lut = "off";
defparam \Add20~17 .lut_mask = 64'h0000FFFF0000AA55;
defparam \Add20~17 .shared_arith = "off";

arriaii_lcell_comb \Selector129~0 (
	.dataa(!\trk_block:sig_trk_state.s_trk_adjust_resync~q ),
	.datab(!\Add20~1_sumout ),
	.datac(!\Add20~5_sumout ),
	.datad(!\Add20~9_sumout ),
	.datae(!\Add20~13_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector129~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector129~0 .extended_lut = "off";
defparam \Selector129~0 .lut_mask = 64'h0000000100000001;
defparam \Selector129~0 .shared_arith = "off";

arriaii_lcell_comb \Add20~21 (
	.dataa(!\trk_block:sig_rsc_drift[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_rsc_drift[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add20~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add20~21_sumout ),
	.cout(\Add20~22 ),
	.shareout());
defparam \Add20~21 .extended_lut = "off";
defparam \Add20~21 .lut_mask = 64'h0000FFFF0000AA55;
defparam \Add20~21 .shared_arith = "off";

arriaii_lcell_comb \Add20~25 (
	.dataa(!\trk_block:sig_rsc_drift[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\trk_block:sig_rsc_drift[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add20~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add20~25_sumout ),
	.cout(\Add20~26 ),
	.shareout());
defparam \Add20~25 .extended_lut = "off";
defparam \Add20~25 .lut_mask = 64'h0000FFFF0000AA55;
defparam \Add20~25 .shared_arith = "off";

arriaii_lcell_comb \Add20~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add20~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add20~29_sumout ),
	.cout(),
	.shareout());
defparam \Add20~29 .extended_lut = "off";
defparam \Add20~29 .lut_mask = 64'h0000FFFF00000000;
defparam \Add20~29 .shared_arith = "off";

arriaii_lcell_comb \Selector129~2 (
	.dataa(!\Selector128~1_combout ),
	.datab(!\Add20~17_sumout ),
	.datac(!\Selector129~0_combout ),
	.datad(!\Add20~21_sumout ),
	.datae(!\Add20~25_sumout ),
	.dataf(!\Add20~29_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector129~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector129~2 .extended_lut = "off";
defparam \Selector129~2 .lut_mask = 64'h5555555755555555;
defparam \Selector129~2 .shared_arith = "off";

dffeas sig_trk_err(
	.clk(clk),
	.d(\Selector129~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_track~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_trk_err~q ),
	.prn(vcc));
defparam sig_trk_err.is_wysiwyg = "true";
defparam sig_trk_err.power_up = "low";

arriaii_lcell_comb \sig_cmd_err~0 (
	.dataa(!q_b_1),
	.datab(!q_b_3),
	.datac(!q_b_17),
	.datad(!q_b_19),
	.datae(!q_b_33),
	.dataf(!q_b_35),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_cmd_err~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_cmd_err~0 .extended_lut = "off";
defparam \sig_cmd_err~0 .lut_mask = 64'h8000040000200001;
defparam \sig_cmd_err~0 .shared_arith = "off";

arriaii_lcell_comb \sig_cmd_err~1 (
	.dataa(!q_b_5),
	.datab(!q_b_7),
	.datac(!q_b_21),
	.datad(!q_b_23),
	.datae(!q_b_37),
	.dataf(!q_b_39),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_cmd_err~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_cmd_err~1 .extended_lut = "off";
defparam \sig_cmd_err~1 .lut_mask = 64'h8000040000200001;
defparam \sig_cmd_err~1 .shared_arith = "off";

arriaii_lcell_comb \sig_cmd_err~3 (
	.dataa(!q_b_0),
	.datab(!q_b_16),
	.datac(!q_b_32),
	.datad(!q_b_48),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_cmd_err~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_cmd_err~3 .extended_lut = "off";
defparam \sig_cmd_err~3 .lut_mask = 64'h8001800180018001;
defparam \sig_cmd_err~3 .shared_arith = "off";

arriaii_lcell_comb \sig_cmd_err~4 (
	.dataa(!q_b_2),
	.datab(!q_b_18),
	.datac(!q_b_34),
	.datad(!q_b_50),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_cmd_err~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_cmd_err~4 .extended_lut = "off";
defparam \sig_cmd_err~4 .lut_mask = 64'h8001800180018001;
defparam \sig_cmd_err~4 .shared_arith = "off";

arriaii_lcell_comb \sig_cmd_err~6 (
	.dataa(!q_b_1),
	.datab(!q_b_3),
	.datac(!q_b_49),
	.datad(!q_b_51),
	.datae(!q_b_7),
	.dataf(!q_b_55),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_cmd_err~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_cmd_err~6 .extended_lut = "off";
defparam \sig_cmd_err~6 .lut_mask = 64'h8421000000008421;
defparam \sig_cmd_err~6 .shared_arith = "off";

arriaii_lcell_comb \sig_cmd_err~7 (
	.dataa(!q_b_5),
	.datab(!q_b_53),
	.datac(!q_b_6),
	.datad(!q_b_22),
	.datae(!q_b_38),
	.dataf(!q_b_54),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_cmd_err~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_cmd_err~7 .extended_lut = "off";
defparam \sig_cmd_err~7 .lut_mask = 64'h9000000000000009;
defparam \sig_cmd_err~7 .shared_arith = "off";

arriaii_lcell_comb \sig_cmd_err~5 (
	.dataa(!\sig_cmd_err~2_combout ),
	.datab(!\sig_cmd_err~3_combout ),
	.datac(!\sig_cmd_err~4_combout ),
	.datad(!\sig_cmd_err~6_combout ),
	.datae(!\sig_cmd_err~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_cmd_err~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_cmd_err~5 .extended_lut = "off";
defparam \sig_cmd_err~5 .lut_mask = 64'h0000000100000001;
defparam \sig_cmd_err~5 .shared_arith = "off";

arriaii_lcell_comb \Selector32~2 (
	.dataa(!\Selector32~0_combout ),
	.datab(!sig_addr_cmd0cke0),
	.datac(!\sig_cmd_err~0_combout ),
	.datad(!\sig_cmd_err~1_combout ),
	.datae(!\sig_cmd_err~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector32~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector32~2 .extended_lut = "off";
defparam \Selector32~2 .lut_mask = 64'h1111111011111110;
defparam \Selector32~2 .shared_arith = "off";

arriaii_lcell_comb \Selector32~3 (
	.dataa(!\Selector32~1_combout ),
	.datab(!\Selector32~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector32~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector32~3 .extended_lut = "off";
defparam \Selector32~3 .lut_mask = 64'h7777777777777777;
defparam \Selector32~3 .shared_arith = "off";

dffeas sig_cmd_err(
	.clk(clk),
	.d(\Selector32~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_cmd_err~q ),
	.prn(vcc));
defparam sig_cmd_err.is_wysiwyg = "true";
defparam sig_cmd_err.power_up = "low";

arriaii_lcell_comb \dgrb_ctrl~0 (
	.dataa(!\sig_dgrb_state.s_seek_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\ctrl_dgrb_r.command.cmd_read_mtp~q ),
	.datad(!\sig_rsc_err~q ),
	.datae(!\sig_trk_err~q ),
	.dataf(!\sig_cmd_err~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dgrb_ctrl~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dgrb_ctrl~0 .extended_lut = "off";
defparam \dgrb_ctrl~0 .lut_mask = 64'h0050207080D0A0F0;
defparam \dgrb_ctrl~0 .shared_arith = "off";

arriaii_lcell_comb \seq_pll_select~0 (
	.dataa(!\sig_dgrb_state.s_track~q ),
	.datab(!sig_addr_cmd0cke0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_pll_select~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_pll_select~0 .extended_lut = "off";
defparam \seq_pll_select~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \seq_pll_select~0 .shared_arith = "off";

arriaii_lcell_comb \sig_trk_pll_select[1]~0 (
	.dataa(!\sig_trk_pll_inc_dec_n~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_trk_pll_select[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_trk_pll_select[1]~0 .extended_lut = "off";
defparam \sig_trk_pll_select[1]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \sig_trk_pll_select[1]~0 .shared_arith = "off";

dffeas \sig_trk_pll_select[1] (
	.clk(clk),
	.d(\sig_trk_pll_select[1]~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_trk_pll_select[1]~q ),
	.prn(vcc));
defparam \sig_trk_pll_select[1] .is_wysiwyg = "true";
defparam \sig_trk_pll_select[1] .power_up = "low";

arriaii_lcell_comb \seq_pll_select~1 (
	.dataa(!\sig_dgrb_state.s_seek_cdvw~q ),
	.datab(!\sig_dgrb_state.s_reset_cdvw~q ),
	.datac(!\sig_dgrb_state.s_test_phases~q ),
	.datad(!\sig_dgrb_state.s_track~q ),
	.datae(!\sig_trk_pll_select[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_pll_select~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_pll_select~1 .extended_lut = "off";
defparam \seq_pll_select~1 .lut_mask = 64'h8000808080008080;
defparam \seq_pll_select~1 .shared_arith = "off";

arriaii_lcell_comb \Selector179~0 (
	.dataa(!\ac_block:sig_burst_count[0]~q ),
	.datab(!\ac_block:sig_addr_cmd_state.s_ac_read_wd_lat~q ),
	.datac(!\ac_block:sig_addr_cmd_last_state.s_ac_read_wd_lat~q ),
	.datad(!\ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ),
	.datae(!\ac_block:sig_addr_cmd_last_state.s_ac_read_rdv~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector179~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector179~0 .extended_lut = "off";
defparam \Selector179~0 .lut_mask = 64'h020202AA020202AA;
defparam \Selector179~0 .shared_arith = "off";

arriaii_lcell_comb \Selector179~1 (
	.dataa(gnd),
	.datab(!\Equal21~1_combout ),
	.datac(!\Selector153~1_combout ),
	.datad(!\Selector183~0_combout ),
	.datae(!\Selector179~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector179~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector179~1 .extended_lut = "off";
defparam \Selector179~1 .lut_mask = 64'h0F3FFFFF0F3FFFFF;
defparam \Selector179~1 .shared_arith = "off";

arriaii_lcell_comb \btp_addr_array~0 (
	.dataa(!\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.datab(!\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\btp_addr_array~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \btp_addr_array~0 .extended_lut = "off";
defparam \btp_addr_array~0 .lut_mask = 64'h7777777777777777;
defparam \btp_addr_array~0 .shared_arith = "off";

dffeas \ac_block:btp_addr_array[0][4] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btp_addr_array~0_combout ),
	.q(\ac_block:btp_addr_array[0][4]~q ),
	.prn(vcc));
defparam \ac_block:btp_addr_array[0][4] .is_wysiwyg = "true";
defparam \ac_block:btp_addr_array[0][4] .power_up = "low";

dffeas \ctrl_dgrb_r.command_op.mtp_almt (
	.clk(clk),
	.d(\ctrl_dgrb.command_op.mtp_almt ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_dgrb_r.command_op.mtp_almt~q ),
	.prn(vcc));
defparam \ctrl_dgrb_r.command_op.mtp_almt .is_wysiwyg = "true";
defparam \ctrl_dgrb_r.command_op.mtp_almt .power_up = "low";

dffeas current_mtp_almt(
	.clk(clk),
	.d(\ctrl_dgrb_r.command_op.mtp_almt~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ac_muxctrl_broadcast_rcommand_req),
	.q(\current_mtp_almt~q ),
	.prn(vcc));
defparam current_mtp_almt.is_wysiwyg = "true";
defparam current_mtp_almt.power_up = "low";

dffeas \ac_block:btp_addr_array[0][3] (
	.clk(clk),
	.d(\current_mtp_almt~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btp_addr_array~0_combout ),
	.q(\ac_block:btp_addr_array[0][3]~q ),
	.prn(vcc));
defparam \ac_block:btp_addr_array[0][3] .is_wysiwyg = "true";
defparam \ac_block:btp_addr_array[0][3] .power_up = "low";

arriaii_lcell_comb \Selector153~2 (
	.dataa(!\ac_block:sig_count[0]~q ),
	.datab(!\Equal21~1_combout ),
	.datac(!\Selector183~0_combout ),
	.datad(!\ac_block:btp_addr_array[0][4]~q ),
	.datae(!\ac_block:btp_addr_array[0][3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector153~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector153~2 .extended_lut = "off";
defparam \Selector153~2 .lut_mask = 64'h0001020300010203;
defparam \Selector153~2 .shared_arith = "off";

arriaii_lcell_comb \Selector153~3 (
	.dataa(!\ac_block:sig_burst_count[0]~q ),
	.datab(!\ac_block:sig_addr_cmd_state.s_ac_read_wd_lat~q ),
	.datac(!\ac_block:sig_addr_cmd_last_state.s_ac_read_wd_lat~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector153~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector153~3 .extended_lut = "off";
defparam \Selector153~3 .lut_mask = 64'h3131313131313131;
defparam \Selector153~3 .shared_arith = "off";

arriaii_lcell_comb \sig_addr_cmd~0 (
	.dataa(!\ac_block:sig_burst_count[0]~q ),
	.datab(!\ac_block:sig_addr_cmd_last_state.s_ac_read_mtp~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_addr_cmd~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_addr_cmd~0 .extended_lut = "off";
defparam \sig_addr_cmd~0 .lut_mask = 64'h2222222222222222;
defparam \sig_addr_cmd~0 .shared_arith = "off";

arriaii_lcell_comb \Selector152~0 (
	.dataa(!\ac_block:sig_burst_count[0]~q ),
	.datab(!dgb_ac_access_gnt_r),
	.datac(!\ac_block:sig_addr_cmd_last_state.s_ac_read_poa_mtp~q ),
	.datad(!\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector152~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector152~0 .extended_lut = "off";
defparam \Selector152~0 .lut_mask = 64'h00FD00FD00FD00FD;
defparam \Selector152~0 .shared_arith = "off";

arriaii_lcell_comb \Selector152~1 (
	.dataa(!\ac_block:sig_burst_count[0]~q ),
	.datab(!\ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ),
	.datac(!\ac_block:sig_addr_cmd_state.s_ac_relax~q ),
	.datad(!\ac_block:sig_addr_cmd_last_state.s_ac_read_rdv~q ),
	.datae(!\Selector152~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector152~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector152~1 .extended_lut = "off";
defparam \Selector152~1 .lut_mask = 64'hC0E00000C0E00000;
defparam \Selector152~1 .shared_arith = "off";

arriaii_lcell_comb \Selector152~2 (
	.dataa(gnd),
	.datab(!\Equal21~1_combout ),
	.datac(!\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.datad(!\sig_addr_cmd~0_combout ),
	.datae(!\Selector152~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector152~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector152~2 .extended_lut = "off";
defparam \Selector152~2 .lut_mask = 64'h0000F0F30000F0F3;
defparam \Selector152~2 .shared_arith = "off";

arriaii_lcell_comb \Selector153~4 (
	.dataa(!\ac_block:sig_burst_count[0]~q ),
	.datab(!\Equal21~0_combout ),
	.datac(!\ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ),
	.datad(!\ac_block:sig_addr_cmd_last_state.s_ac_read_rdv~q ),
	.datae(!\Selector153~1_combout ),
	.dataf(!\current_mtp_almt~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector153~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector153~4 .extended_lut = "off";
defparam \Selector153~4 .lut_mask = 64'h0008333B00080008;
defparam \Selector153~4 .shared_arith = "off";

arriaii_lcell_comb \Selector153~5 (
	.dataa(!sig_addr_cmd0addr3),
	.datab(!\Selector153~2_combout ),
	.datac(!\Selector153~3_combout ),
	.datad(!\Selector152~2_combout ),
	.datae(!\Selector153~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector153~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector153~5 .extended_lut = "off";
defparam \Selector153~5 .lut_mask = 64'h7737FFFF7737FFFF;
defparam \Selector153~5 .shared_arith = "off";

arriaii_lcell_comb \Selector152~3 (
	.dataa(!\ac_block:sig_burst_count[0]~q ),
	.datab(!\ac_block:sig_addr_cmd_state.s_ac_read_wd_lat~q ),
	.datac(!\ac_block:sig_addr_cmd_last_state.s_ac_read_wd_lat~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector152~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector152~3 .extended_lut = "off";
defparam \Selector152~3 .lut_mask = 64'h0202020202020202;
defparam \Selector152~3 .shared_arith = "off";

arriaii_lcell_comb \Selector152~4 (
	.dataa(!\ac_block:sig_count[0]~q ),
	.datab(!\Equal21~1_combout ),
	.datac(!\Selector153~1_combout ),
	.datad(!\Selector183~0_combout ),
	.datae(!\ac_block:btp_addr_array[0][4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector152~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector152~4 .extended_lut = "off";
defparam \Selector152~4 .lut_mask = 64'h0202022202020222;
defparam \Selector152~4 .shared_arith = "off";

arriaii_lcell_comb \Selector152~5 (
	.dataa(!\ac_block:sig_addr_cmd_state.s_ac_read_wd_lat~q ),
	.datab(!sig_addr_cmd0addr4),
	.datac(!\Selector152~3_combout ),
	.datad(!\Selector152~2_combout ),
	.datae(!\Selector152~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector152~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector152~5 .extended_lut = "off";
defparam \Selector152~5 .lut_mask = 64'h3F1FFFFF3F1FFFFF;
defparam \Selector152~5 .shared_arith = "off";

arriaii_lcell_comb \Selector151~0 (
	.dataa(!\ac_block:sig_count[0]~q ),
	.datab(!\Equal21~1_combout ),
	.datac(!\Selector183~0_combout ),
	.datad(!\ac_block:btp_addr_array[0][4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector151~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector151~0 .extended_lut = "off";
defparam \Selector151~0 .lut_mask = 64'h0001000100010001;
defparam \Selector151~0 .shared_arith = "off";

arriaii_lcell_comb \Selector151~1 (
	.dataa(!\ac_block:sig_addr_cmd_state.s_ac_read_wd_lat~q ),
	.datab(!sig_addr_cmd0addr5),
	.datac(!\Selector152~3_combout ),
	.datad(!\Selector152~2_combout ),
	.datae(!\Selector151~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector151~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector151~1 .extended_lut = "off";
defparam \Selector151~1 .lut_mask = 64'h3F1FFFFF3F1FFFFF;
defparam \Selector151~1 .shared_arith = "off";

arriaii_lcell_comb \sig_addr_cmd[0].addr[12]~0 (
	.dataa(!\ac_block:sig_burst_count[0]~q ),
	.datab(!\ac_block:sig_count[0]~q ),
	.datac(!\Equal21~1_combout ),
	.datad(!\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.datae(!\Selector188~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_addr_cmd[0].addr[12]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_addr_cmd[0].addr[12]~0 .extended_lut = "off";
defparam \sig_addr_cmd[0].addr[12]~0 .lut_mask = 64'h55F300F055F300F0;
defparam \sig_addr_cmd[0].addr[12]~0 .shared_arith = "off";

arriaii_lcell_comb \sig_addr_cmd[0].addr[12]~1 (
	.dataa(!\ac_block:sig_addr_cmd_state.s_ac_read_wd_lat~q ),
	.datab(!\ac_block:sig_addr_cmd_last_state.s_ac_read_wd_lat~q ),
	.datac(!\ac_block:sig_addr_cmd_state.s_ac_read_rdv~q ),
	.datad(!\ac_block:sig_addr_cmd_state.s_ac_relax~q ),
	.datae(!\ac_block:sig_addr_cmd_last_state.s_ac_read_rdv~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_addr_cmd[0].addr[12]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_addr_cmd[0].addr[12]~1 .extended_lut = "off";
defparam \sig_addr_cmd[0].addr[12]~1 .lut_mask = 64'hB100BB00B100BB00;
defparam \sig_addr_cmd[0].addr[12]~1 .shared_arith = "off";

arriaii_lcell_comb \sig_addr_cmd[0].addr[12]~2 (
	.dataa(!dgb_ac_access_gnt_r),
	.datab(!\ac_block:sig_addr_cmd_last_state.s_ac_read_poa_mtp~q ),
	.datac(!\ac_block:sig_addr_cmd_state.s_ac_read_poa_mtp~q ),
	.datad(!\ac_block:sig_addr_cmd_state.s_ac_read_mtp~q ),
	.datae(!\sig_addr_cmd~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_addr_cmd[0].addr[12]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_addr_cmd[0].addr[12]~2 .extended_lut = "off";
defparam \sig_addr_cmd[0].addr[12]~2 .lut_mask = 64'hF100F1F1F100F1F1;
defparam \sig_addr_cmd[0].addr[12]~2 .shared_arith = "off";

arriaii_lcell_comb \sig_addr_cmd[0].addr[12]~3 (
	.dataa(!\ac_block:sig_addr_cmd_state.s_ac_idle~q ),
	.datab(!sig_addr_cmd0addr12),
	.datac(!\sig_addr_cmd[0].addr[12]~0_combout ),
	.datad(!\sig_addr_cmd[0].addr[12]~1_combout ),
	.datae(!\sig_addr_cmd[0].addr[12]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_addr_cmd[0].addr[12]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_addr_cmd[0].addr[12]~3 .extended_lut = "off";
defparam \sig_addr_cmd[0].addr[12]~3 .lut_mask = 64'h3333335333333353;
defparam \sig_addr_cmd[0].addr[12]~3 .shared_arith = "off";

dffeas \sig_dgrb_last_state.s_idle (
	.clk(clk),
	.d(\sig_dgrb_state.s_idle~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgrb_last_state.s_idle~q ),
	.prn(vcc));
defparam \sig_dgrb_last_state.s_idle .is_wysiwyg = "true";
defparam \sig_dgrb_last_state.s_idle .power_up = "low";

arriaii_lcell_comb \ac_handshake_proc~3 (
	.dataa(!\sig_dgrb_state.s_wait_admin~q ),
	.datab(!\sig_dgrb_last_state.s_idle~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_handshake_proc~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_handshake_proc~3 .extended_lut = "off";
defparam \ac_handshake_proc~3 .lut_mask = 64'h4444444444444444;
defparam \ac_handshake_proc~3 .shared_arith = "off";

arriaii_lcell_comb \seq_poa_lat_dec_1x~0 (
	.dataa(!\sig_dgrb_state.s_poa_cal~q ),
	.datab(!\poa_block:sig_poa_state~q ),
	.datac(!\sig_poa_match_en~q ),
	.datad(!\sig_poa_match~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_poa_lat_dec_1x~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_poa_lat_dec_1x~0 .extended_lut = "off";
defparam \seq_poa_lat_dec_1x~0 .lut_mask = 64'h0400040004000400;
defparam \seq_poa_lat_dec_1x~0 .shared_arith = "off";

arriaii_lcell_comb \dgrb_ctrl~1 (
	.dataa(!\ctrl_dgrb_r.command.cmd_read_mtp~q ),
	.datab(!\sig_cdvw_state.largest_window_size[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dgrb_ctrl~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dgrb_ctrl~1 .extended_lut = "off";
defparam \dgrb_ctrl~1 .lut_mask = 64'h1111111111111111;
defparam \dgrb_ctrl~1 .shared_arith = "off";

dffeas \sig_cmd_result[2] (
	.clk(clk),
	.d(\Selector32~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_cmd_result[2]~q ),
	.prn(vcc));
defparam \sig_cmd_result[2] .is_wysiwyg = "true";
defparam \sig_cmd_result[2] .power_up = "low";

dffeas \sig_cdvw_state.largest_window_size[2] (
	.clk(clk),
	.d(\sig_cdvw_state.current_window_size[2]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\v_cdvw_state~2_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.largest_window_centre[1]~0_combout ),
	.q(\sig_cdvw_state.largest_window_size[2]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.largest_window_size[2] .is_wysiwyg = "true";
defparam \sig_cdvw_state.largest_window_size[2] .power_up = "low";

dffeas \sig_trk_result[2] (
	.clk(clk),
	.d(\Selector128~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_track~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_trk_result[2]~q ),
	.prn(vcc));
defparam \sig_trk_result[2] .is_wysiwyg = "true";
defparam \sig_trk_result[2] .power_up = "low";

arriaii_lcell_comb \sig_rsc_result[2]~3 (
	.dataa(!\sig_cdvw_state.status.valid_result~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_rsc_result[2]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_rsc_result[2]~3 .extended_lut = "off";
defparam \sig_rsc_result[2]~3 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \sig_rsc_result[2]~3 .shared_arith = "off";

dffeas \sig_rsc_result[2] (
	.clk(clk),
	.d(\sig_rsc_result[2]~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_rsc_result[0]~0_combout ),
	.q(\sig_rsc_result[2]~q ),
	.prn(vcc));
defparam \sig_rsc_result[2] .is_wysiwyg = "true";
defparam \sig_rsc_result[2] .power_up = "low";

arriaii_lcell_comb \dgrb_ctrl.command_result[3]~0 (
	.dataa(!\sig_dgrb_state.s_seek_cdvw~q ),
	.datab(!\ctrl_dgrb_r.command.cmd_read_mtp~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dgrb_ctrl.command_result[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dgrb_ctrl.command_result[3]~0 .extended_lut = "off";
defparam \dgrb_ctrl.command_result[3]~0 .lut_mask = 64'h8888888888888888;
defparam \dgrb_ctrl.command_result[3]~0 .shared_arith = "off";

arriaii_lcell_comb \dgrb_ctrl.command_result[3]~1 (
	.dataa(!\sig_dgrb_state.s_seek_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\ctrl_dgrb_r.command.cmd_read_mtp~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dgrb_ctrl.command_result[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dgrb_ctrl.command_result[3]~1 .extended_lut = "off";
defparam \dgrb_ctrl.command_result[3]~1 .lut_mask = 64'h7070707070707070;
defparam \dgrb_ctrl.command_result[3]~1 .shared_arith = "off";

arriaii_lcell_comb \dgrb_ctrl~2 (
	.dataa(!\sig_cmd_result[2]~q ),
	.datab(!\sig_cdvw_state.largest_window_size[2]~q ),
	.datac(!\sig_trk_result[2]~q ),
	.datad(!\sig_rsc_result[2]~q ),
	.datae(!\dgrb_ctrl.command_result[3]~0_combout ),
	.dataf(!\dgrb_ctrl.command_result[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dgrb_ctrl~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dgrb_ctrl~2 .extended_lut = "off";
defparam \dgrb_ctrl~2 .lut_mask = 64'h3333555500FF0F0F;
defparam \dgrb_ctrl~2 .shared_arith = "off";

arriaii_lcell_comb \v_cdvw_state~29 (
	.dataa(!\sig_cdvw_state.valid_phase_seen~q ),
	.datab(!\find_centre_of_largest_data_valid_window~1_combout ),
	.datac(!\v_cdvw_state~1_combout ),
	.datad(!\cdvw_proc~1_combout ),
	.datae(!\cdvw_proc~2_combout ),
	.dataf(!\sig_cdvw_state.status.no_valid_phases~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~29 .extended_lut = "off";
defparam \v_cdvw_state~29 .lut_mask = 64'h0D00FF00FD00FF00;
defparam \v_cdvw_state~29 .shared_arith = "off";

dffeas \sig_cdvw_state.status.no_valid_phases (
	.clk(clk),
	.d(\v_cdvw_state~29_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_cdvw_state.status.no_valid_phases~q ),
	.prn(vcc));
defparam \sig_cdvw_state.status.no_valid_phases .is_wysiwyg = "true";
defparam \sig_cdvw_state.status.no_valid_phases .power_up = "low";

arriaii_lcell_comb \Selector131~1 (
	.dataa(!\Selector128~1_combout ),
	.datab(!\sig_cdvw_state.status.no_valid_phases~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector131~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector131~1 .extended_lut = "off";
defparam \Selector131~1 .lut_mask = 64'h1111111111111111;
defparam \Selector131~1 .shared_arith = "off";

arriaii_lcell_comb \Selector131~0 (
	.dataa(!\Add20~17_sumout ),
	.datab(!\Selector129~0_combout ),
	.datac(!\Add20~21_sumout ),
	.datad(!\Add20~25_sumout ),
	.datae(!\Add20~29_sumout ),
	.dataf(!\Selector131~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector131~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector131~0 .extended_lut = "off";
defparam \Selector131~0 .lut_mask = 64'h00010000FFFFFFFF;
defparam \Selector131~0 .shared_arith = "off";

dffeas \sig_trk_result[1] (
	.clk(clk),
	.d(\Selector131~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_track~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_trk_result[1]~q ),
	.prn(vcc));
defparam \sig_trk_result[1] .is_wysiwyg = "true";
defparam \sig_trk_result[1] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~30 (
	.dataa(!\sig_cdvw_state.valid_phase_seen~q ),
	.datab(!\find_centre_of_largest_data_valid_window~1_combout ),
	.datac(!\v_cdvw_state~1_combout ),
	.datad(!\v_cdvw_state~2_combout ),
	.datae(!\sig_cdvw_state.status.no_invalid_phases~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~30 .extended_lut = "off";
defparam \v_cdvw_state~30 .lut_mask = 64'h0100F1000100F100;
defparam \v_cdvw_state~30 .shared_arith = "off";

dffeas \sig_cdvw_state.status.no_invalid_phases (
	.clk(clk),
	.d(\v_cdvw_state~30_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_cdvw_state.status.no_invalid_phases~q ),
	.prn(vcc));
defparam \sig_cdvw_state.status.no_invalid_phases .is_wysiwyg = "true";
defparam \sig_cdvw_state.status.no_invalid_phases .power_up = "low";

arriaii_lcell_comb \sig_rsc_result~1 (
	.dataa(!\sig_cdvw_state.status.no_valid_phases~q ),
	.datab(!\sig_cdvw_state.status.no_invalid_phases~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_rsc_result~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_rsc_result~1 .extended_lut = "off";
defparam \sig_rsc_result~1 .lut_mask = 64'h4444444444444444;
defparam \sig_rsc_result~1 .shared_arith = "off";

dffeas \sig_rsc_result[1] (
	.clk(clk),
	.d(\sig_rsc_result~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_cdvw_state.status.valid_result~q ),
	.sload(gnd),
	.ena(\sig_rsc_result[0]~0_combout ),
	.q(\sig_rsc_result[1]~q ),
	.prn(vcc));
defparam \sig_rsc_result[1] .is_wysiwyg = "true";
defparam \sig_rsc_result[1] .power_up = "low";

arriaii_lcell_comb \dgrb_ctrl~3 (
	.dataa(!\sig_cmd_result[2]~q ),
	.datab(!\sig_cdvw_state.largest_window_size[1]~q ),
	.datac(!\sig_trk_result[1]~q ),
	.datad(!\sig_rsc_result[1]~q ),
	.datae(!\dgrb_ctrl.command_result[3]~0_combout ),
	.dataf(!\dgrb_ctrl.command_result[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dgrb_ctrl~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dgrb_ctrl~3 .extended_lut = "off";
defparam \dgrb_ctrl~3 .lut_mask = 64'h3333555500FF0F0F;
defparam \dgrb_ctrl~3 .shared_arith = "off";

arriaii_lcell_comb \Add0~1 (
	.dataa(!rdata_valid[0]),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dgrb_main_block:sig_count[0]~q ),
	.datae(gnd),
	.dataf(!seq_rdata_valid_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000055FF000000FF;
defparam \Add0~1 .shared_arith = "off";

arriaii_lcell_comb \dgrb_main_block:sig_count[0]~0 (
	.dataa(!\sig_dimm_driving_dq~q ),
	.datab(!\sig_dgrb_state.s_idle~q ),
	.datac(!\sig_dgrb_state.s_adv_rd_lat_setup~q ),
	.datad(!\sig_dgrb_state.s_adv_rd_lat~q ),
	.datae(!\sig_dgrb_last_state.s_adv_rd_lat_setup~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dgrb_main_block:sig_count[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dgrb_main_block:sig_count[0]~0 .extended_lut = "off";
defparam \dgrb_main_block:sig_count[0]~0 .lut_mask = 64'hCFAAC0A0CFAAC0A0;
defparam \dgrb_main_block:sig_count[0]~0 .shared_arith = "off";

dffeas \dgrb_main_block:sig_count[0] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_adv_rd_lat~q ),
	.sload(gnd),
	.ena(\dgrb_main_block:sig_count[0]~0_combout ),
	.q(\dgrb_main_block:sig_count[0]~q ),
	.prn(vcc));
defparam \dgrb_main_block:sig_count[0] .is_wysiwyg = "true";
defparam \dgrb_main_block:sig_count[0] .power_up = "low";

arriaii_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dgrb_main_block:sig_count[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \dgrb_main_block:sig_count[1] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_adv_rd_lat~q ),
	.sload(gnd),
	.ena(\dgrb_main_block:sig_count[0]~0_combout ),
	.q(\dgrb_main_block:sig_count[1]~q ),
	.prn(vcc));
defparam \dgrb_main_block:sig_count[1] .is_wysiwyg = "true";
defparam \dgrb_main_block:sig_count[1] .power_up = "low";

arriaii_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dgrb_main_block:sig_count[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \dgrb_main_block:sig_count[2] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_adv_rd_lat~q ),
	.sload(gnd),
	.ena(\dgrb_main_block:sig_count[0]~0_combout ),
	.q(\dgrb_main_block:sig_count[2]~q ),
	.prn(vcc));
defparam \dgrb_main_block:sig_count[2] .is_wysiwyg = "true";
defparam \dgrb_main_block:sig_count[2] .power_up = "low";

arriaii_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dgrb_main_block:sig_count[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \dgrb_main_block:sig_count[3] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_adv_rd_lat~q ),
	.sload(gnd),
	.ena(\dgrb_main_block:sig_count[0]~0_combout ),
	.q(\dgrb_main_block:sig_count[3]~q ),
	.prn(vcc));
defparam \dgrb_main_block:sig_count[3] .is_wysiwyg = "true";
defparam \dgrb_main_block:sig_count[3] .power_up = "low";

arriaii_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dgrb_main_block:sig_count[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \dgrb_main_block:sig_count[4] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_adv_rd_lat~q ),
	.sload(gnd),
	.ena(\dgrb_main_block:sig_count[0]~0_combout ),
	.q(\dgrb_main_block:sig_count[4]~q ),
	.prn(vcc));
defparam \dgrb_main_block:sig_count[4] .is_wysiwyg = "true";
defparam \dgrb_main_block:sig_count[4] .power_up = "low";

arriaii_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dgrb_main_block:sig_count[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \dgrb_main_block:sig_count[5] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_adv_rd_lat~q ),
	.sload(gnd),
	.ena(\dgrb_main_block:sig_count[0]~0_combout ),
	.q(\dgrb_main_block:sig_count[5]~q ),
	.prn(vcc));
defparam \dgrb_main_block:sig_count[5] .is_wysiwyg = "true";
defparam \dgrb_main_block:sig_count[5] .power_up = "low";

arriaii_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dgrb_main_block:sig_count[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~25 .shared_arith = "off";

dffeas \dgrb_main_block:sig_count[6] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_adv_rd_lat~q ),
	.sload(gnd),
	.ena(\dgrb_main_block:sig_count[0]~0_combout ),
	.q(\dgrb_main_block:sig_count[6]~q ),
	.prn(vcc));
defparam \dgrb_main_block:sig_count[6] .is_wysiwyg = "true";
defparam \dgrb_main_block:sig_count[6] .power_up = "low";

arriaii_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dgrb_main_block:sig_count[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add0~29 .shared_arith = "off";

dffeas \dgrb_main_block:sig_count[7] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_adv_rd_lat~q ),
	.sload(gnd),
	.ena(\dgrb_main_block:sig_count[0]~0_combout ),
	.q(\dgrb_main_block:sig_count[7]~q ),
	.prn(vcc));
defparam \dgrb_main_block:sig_count[7] .is_wysiwyg = "true";
defparam \dgrb_main_block:sig_count[7] .power_up = "low";

arriaii_lcell_comb \Selector32~1 (
	.dataa(!\sig_dimm_driving_dq~q ),
	.datab(!\sig_dgrb_state.s_adv_rd_lat~q ),
	.datac(!\dgrb_main_block:sig_count[7]~q ),
	.datad(!\dgrb_main_block:sig_count[6]~q ),
	.datae(!\dgrb_main_block:sig_count[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector32~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector32~1 .extended_lut = "off";
defparam \Selector32~1 .lut_mask = 64'h0222222202222222;
defparam \Selector32~1 .shared_arith = "off";

dffeas \sig_cmd_result[3] (
	.clk(clk),
	.d(\Selector32~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_cmd_result[3]~q ),
	.prn(vcc));
defparam \sig_cmd_result[3] .is_wysiwyg = "true";
defparam \sig_cmd_result[3] .power_up = "low";

dffeas \sig_cdvw_state.largest_window_size[0] (
	.clk(clk),
	.d(\sig_cdvw_state.current_window_size[0]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\v_cdvw_state~2_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.largest_window_centre[1]~0_combout ),
	.q(\sig_cdvw_state.largest_window_size[0]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.largest_window_size[0] .is_wysiwyg = "true";
defparam \sig_cdvw_state.largest_window_size[0] .power_up = "low";

arriaii_lcell_comb \v_cdvw_state~31 (
	.dataa(!\find_centre_of_largest_data_valid_window~1_combout ),
	.datab(!\v_cdvw_state~1_combout ),
	.datac(!\sig_cdvw_state.multiple_eq_windows~q ),
	.datad(!\v_cdvw_state~2_combout ),
	.datae(!\sig_cdvw_state.status.multiple_equal_windows~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\v_cdvw_state~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \v_cdvw_state~31 .extended_lut = "off";
defparam \v_cdvw_state~31 .lut_mask = 64'h0200CE000200CE00;
defparam \v_cdvw_state~31 .shared_arith = "off";

dffeas \sig_cdvw_state.status.multiple_equal_windows (
	.clk(clk),
	.d(\v_cdvw_state~31_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_cdvw_state.status.multiple_equal_windows~q ),
	.prn(vcc));
defparam \sig_cdvw_state.status.multiple_equal_windows .is_wysiwyg = "true";
defparam \sig_cdvw_state.status.multiple_equal_windows .power_up = "low";

arriaii_lcell_comb \sig_trk_result~0 (
	.dataa(!\sig_cdvw_state.status.valid_result~q ),
	.datab(!\sig_cdvw_state.status.calculating~q ),
	.datac(!\sig_cdvw_state.status.multiple_equal_windows~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_trk_result~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_trk_result~0 .extended_lut = "off";
defparam \sig_trk_result~0 .lut_mask = 64'h8080808080808080;
defparam \sig_trk_result~0 .shared_arith = "off";

dffeas \sig_trk_result[0] (
	.clk(clk),
	.d(\sig_trk_result~0_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_track~q ),
	.sload(!\trk_block:sig_trk_state.s_trk_cdvw_wait~q ),
	.ena(vcc),
	.q(\sig_trk_result[0]~q ),
	.prn(vcc));
defparam \sig_trk_result[0] .is_wysiwyg = "true";
defparam \sig_trk_result[0] .power_up = "low";

arriaii_lcell_comb \sig_rsc_result~2 (
	.dataa(!\sig_cdvw_state.status.valid_result~q ),
	.datab(!\sig_cdvw_state.status.multiple_equal_windows~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_rsc_result~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_rsc_result~2 .extended_lut = "off";
defparam \sig_rsc_result~2 .lut_mask = 64'h8888888888888888;
defparam \sig_rsc_result~2 .shared_arith = "off";

dffeas \sig_rsc_result[0] (
	.clk(clk),
	.d(\sig_rsc_result~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sig_rsc_result[0]~0_combout ),
	.q(\sig_rsc_result[0]~q ),
	.prn(vcc));
defparam \sig_rsc_result[0] .is_wysiwyg = "true";
defparam \sig_rsc_result[0] .power_up = "low";

arriaii_lcell_comb \dgrb_ctrl~4 (
	.dataa(!\sig_cmd_result[3]~q ),
	.datab(!\sig_cdvw_state.largest_window_size[0]~q ),
	.datac(!\sig_trk_result[0]~q ),
	.datad(!\sig_rsc_result[0]~q ),
	.datae(!\dgrb_ctrl.command_result[3]~0_combout ),
	.dataf(!\dgrb_ctrl.command_result[3]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dgrb_ctrl~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dgrb_ctrl~4 .extended_lut = "off";
defparam \dgrb_ctrl~4 .lut_mask = 64'h3333555500FF0F0F;
defparam \dgrb_ctrl~4 .shared_arith = "off";

arriaii_lcell_comb \Selector129~1 (
	.dataa(!\Add20~17_sumout ),
	.datab(!\Selector129~0_combout ),
	.datac(!\Add20~21_sumout ),
	.datad(!\Add20~25_sumout ),
	.datae(!\Add20~29_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector129~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector129~1 .extended_lut = "off";
defparam \Selector129~1 .lut_mask = 64'h0001000000010000;
defparam \Selector129~1 .shared_arith = "off";

dffeas \sig_trk_result[4] (
	.clk(clk),
	.d(\Selector129~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_track~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_trk_result[4]~q ),
	.prn(vcc));
defparam \sig_trk_result[4] .is_wysiwyg = "true";
defparam \sig_trk_result[4] .power_up = "low";

arriaii_lcell_comb \dgrb_ctrl~5 (
	.dataa(!\sig_cdvw_state.largest_window_size[3]~q ),
	.datab(!\dgrb_ctrl.command_result[3]~0_combout ),
	.datac(!\dgrb_ctrl.command_result[3]~1_combout ),
	.datad(!\sig_cmd_result[3]~q ),
	.datae(!\sig_trk_result[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dgrb_ctrl~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dgrb_ctrl~5 .extended_lut = "off";
defparam \dgrb_ctrl~5 .lut_mask = 64'h4070437340704373;
defparam \dgrb_ctrl~5 .shared_arith = "off";

dffeas \sig_cdvw_state.largest_window_size[4] (
	.clk(clk),
	.d(\sig_cdvw_state.current_window_size[4]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\v_cdvw_state~2_combout ),
	.sload(gnd),
	.ena(\sig_cdvw_state.largest_window_centre[1]~0_combout ),
	.q(\sig_cdvw_state.largest_window_size[4]~q ),
	.prn(vcc));
defparam \sig_cdvw_state.largest_window_size[4] .is_wysiwyg = "true";
defparam \sig_cdvw_state.largest_window_size[4] .power_up = "low";

arriaii_lcell_comb \dgrb_ctrl~6 (
	.dataa(!\sig_dgrb_state.s_seek_cdvw~q ),
	.datab(!\sig_dgrb_state.s_track~q ),
	.datac(!\ctrl_dgrb_r.command.cmd_read_mtp~q ),
	.datad(!\sig_cmd_err~q ),
	.datae(!\sig_cdvw_state.largest_window_size[4]~q ),
	.dataf(!\sig_trk_result[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dgrb_ctrl~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dgrb_ctrl~6 .extended_lut = "off";
defparam \dgrb_ctrl~6 .lut_mask = 64'h00800F8F30B03FBF;
defparam \dgrb_ctrl~6 .shared_arith = "off";

arriaii_lcell_comb \sig_trk_last_state~2 (
	.dataa(!\sig_dgrb_state.s_track~q ),
	.datab(!\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_trk_last_state~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_trk_last_state~2 .extended_lut = "off";
defparam \sig_trk_last_state~2 .lut_mask = 64'h1111111111111111;
defparam \sig_trk_last_state~2 .shared_arith = "off";

dffeas \trk_block:sig_trk_last_state.s_trk_mimic_sample (
	.clk(clk),
	.d(\sig_trk_last_state~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:sig_trk_last_state.s_trk_mimic_sample~q ),
	.prn(vcc));
defparam \trk_block:sig_trk_last_state.s_trk_mimic_sample .is_wysiwyg = "true";
defparam \trk_block:sig_trk_last_state.s_trk_mimic_sample .power_up = "low";

arriaii_lcell_comb \sig_mmc_start~1 (
	.dataa(!\Equal17~1_combout ),
	.datab(!\trk_block:sig_trk_last_state.s_trk_mimic_sample~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_mmc_start~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_mmc_start~1 .extended_lut = "off";
defparam \sig_mmc_start~1 .lut_mask = 64'h8888888888888888;
defparam \sig_mmc_start~1 .shared_arith = "off";

dffeas \trk_block:sig_mmc_start (
	.clk(clk),
	.d(\sig_mmc_start~1_combout ),
	.asdata(GND_port),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\sig_dgrb_state.s_track~q ),
	.sload(!\trk_block:sig_trk_state.s_trk_mimic_sample~q ),
	.ena(vcc),
	.q(\trk_block:sig_mmc_start~q ),
	.prn(vcc));
defparam \trk_block:sig_mmc_start .is_wysiwyg = "true";
defparam \trk_block:sig_mmc_start .power_up = "low";

dffeas \trk_block:mimic_sample_req:seq_mmc_start_r[0] (
	.clk(clk),
	.d(\trk_block:sig_mmc_start~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:mimic_sample_req:seq_mmc_start_r[0]~q ),
	.prn(vcc));
defparam \trk_block:mimic_sample_req:seq_mmc_start_r[0] .is_wysiwyg = "true";
defparam \trk_block:mimic_sample_req:seq_mmc_start_r[0] .power_up = "low";

dffeas \trk_block:mimic_sample_req:seq_mmc_start_r[1] (
	.clk(clk),
	.d(\trk_block:mimic_sample_req:seq_mmc_start_r[0]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:mimic_sample_req:seq_mmc_start_r[1]~q ),
	.prn(vcc));
defparam \trk_block:mimic_sample_req:seq_mmc_start_r[1] .is_wysiwyg = "true";
defparam \trk_block:mimic_sample_req:seq_mmc_start_r[1] .power_up = "low";

dffeas \trk_block:mimic_sample_req:seq_mmc_start_r[2] (
	.clk(clk),
	.d(\trk_block:mimic_sample_req:seq_mmc_start_r[1]~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\trk_block:mimic_sample_req:seq_mmc_start_r[2]~q ),
	.prn(vcc));
defparam \trk_block:mimic_sample_req:seq_mmc_start_r[2] .is_wysiwyg = "true";
defparam \trk_block:mimic_sample_req:seq_mmc_start_r[2] .power_up = "low";

arriaii_lcell_comb \seq_mmc_start~0 (
	.dataa(!\trk_block:sig_mmc_start~q ),
	.datab(!\trk_block:mimic_sample_req:seq_mmc_start_r[0]~q ),
	.datac(!\trk_block:mimic_sample_req:seq_mmc_start_r[2]~q ),
	.datad(!\trk_block:mimic_sample_req:seq_mmc_start_r[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\seq_mmc_start~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \seq_mmc_start~0 .extended_lut = "off";
defparam \seq_mmc_start~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \seq_mmc_start~0 .shared_arith = "off";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_dgwb (
	clk,
	sig_addr_cmd0addr2,
	sig_addr_cmd0addr3,
	sig_addr_cmd0addr4,
	sig_addr_cmd0addr5,
	sig_addr_cmd0cas_n,
	rst_n,
	dgb_ac_access_gnt_r,
	curr_cmdcmd_was,
	curr_cmdcmd_write_btp,
	curr_cmdcmd_write_mtp,
	curr_ctrlcommand_ack,
	dgwb_ctrlcommand_done,
	dgwb_wdp_ovride1,
	ac_muxctrl_broadcast_rcommand_req,
	sig_addr_cmd0cke0,
	dgwb_ac_access_req1,
	sig_addr_cmd1cs_n0,
	sig_addr_cmd0addr12,
	sig_addr_cmd0rst_n,
	dgwb_wdata_120,
	dgwb_wdata_56,
	dgwb_wdata_88,
	dgwb_wdata_24,
	dgwb_wdata_121,
	dgwb_wdata_57,
	dgwb_wdata_89,
	dgwb_wdata_25,
	dgwb_wdata_122,
	dgwb_wdata_58,
	dgwb_wdata_90,
	dgwb_wdata_26,
	dgwb_wdata_123,
	dgwb_wdata_59,
	dgwb_wdata_91,
	dgwb_wdata_27,
	dgwb_wdata_124,
	dgwb_wdata_60,
	dgwb_wdata_92,
	dgwb_wdata_28,
	dgwb_wdata_125,
	dgwb_wdata_61,
	dgwb_wdata_93,
	dgwb_wdata_29,
	dgwb_wdata_126,
	dgwb_wdata_62,
	dgwb_wdata_94,
	dgwb_wdata_30,
	dgwb_wdata_127,
	dgwb_wdata_63,
	dgwb_wdata_95,
	dgwb_wdata_31,
	dgwb_ctrlcommand_ack,
	dgwb_wdp_ovride2)/* synthesis synthesis_greybox=0 */;
input 	clk;
output 	sig_addr_cmd0addr2;
output 	sig_addr_cmd0addr3;
output 	sig_addr_cmd0addr4;
output 	sig_addr_cmd0addr5;
output 	sig_addr_cmd0cas_n;
input 	rst_n;
input 	dgb_ac_access_gnt_r;
input 	curr_cmdcmd_was;
input 	curr_cmdcmd_write_btp;
input 	curr_cmdcmd_write_mtp;
input 	curr_ctrlcommand_ack;
output 	dgwb_ctrlcommand_done;
output 	dgwb_wdp_ovride1;
input 	ac_muxctrl_broadcast_rcommand_req;
output 	sig_addr_cmd0cke0;
output 	dgwb_ac_access_req1;
output 	sig_addr_cmd1cs_n0;
output 	sig_addr_cmd0addr12;
output 	sig_addr_cmd0rst_n;
output 	dgwb_wdata_120;
output 	dgwb_wdata_56;
output 	dgwb_wdata_88;
output 	dgwb_wdata_24;
output 	dgwb_wdata_121;
output 	dgwb_wdata_57;
output 	dgwb_wdata_89;
output 	dgwb_wdata_25;
output 	dgwb_wdata_122;
output 	dgwb_wdata_58;
output 	dgwb_wdata_90;
output 	dgwb_wdata_26;
output 	dgwb_wdata_123;
output 	dgwb_wdata_59;
output 	dgwb_wdata_91;
output 	dgwb_wdata_27;
output 	dgwb_wdata_124;
output 	dgwb_wdata_60;
output 	dgwb_wdata_92;
output 	dgwb_wdata_28;
output 	dgwb_wdata_125;
output 	dgwb_wdata_61;
output 	dgwb_wdata_93;
output 	dgwb_wdata_29;
output 	dgwb_wdata_126;
output 	dgwb_wdata_62;
output 	dgwb_wdata_94;
output 	dgwb_wdata_30;
output 	dgwb_wdata_127;
output 	dgwb_wdata_63;
output 	dgwb_wdata_95;
output 	dgwb_wdata_31;
output 	dgwb_ctrlcommand_ack;
output 	dgwb_wdp_ovride2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add1~1_sumout ;
wire \sig_dgwb_last_state.s_write_01_pairs~q ;
wire \Selector9~4_combout ;
wire \sig_dgwb_state.s_write_01_pairs~q ;
wire \Selector11~5_combout ;
wire \sig_dgwb_last_state.s_write_1100_step~q ;
wire \Selector10~0_combout ;
wire \sig_dgwb_state.s_write_1100_step~q ;
wire \Selector11~6_combout ;
wire \Selector6~0_combout ;
wire \Selector6~1_combout ;
wire \Selector6~2_combout ;
wire \sig_dgwb_state.s_write_ones~q ;
wire \sig_dgwb_last_state.s_write_ones~q ;
wire \Selector5~2_combout ;
wire \sig_dgwb_state.s_write_btp~q ;
wire \sig_dgwb_last_state.s_write_0011_step~q ;
wire \Selector5~3_combout ;
wire \Selector5~4_combout ;
wire \sig_dgwb_last_state.s_write_zeros~q ;
wire \Selector5~5_combout ;
wire \Selector5~6_combout ;
wire \Selector5~7_combout ;
wire \Selector12~0_combout ;
wire \sig_dgwb_state.s_write_wlat~q ;
wire \sig_dgwb_last_state.s_write_wlat~q ;
wire \Selector11~11_combout ;
wire \Selector11~7_combout ;
wire \Selector11~8_combout ;
wire \Selector11~9_combout ;
wire \sig_dgwb_state.s_release_admin~q ;
wire \Selector11~4_combout ;
wire \sig_dgwb_state.s_idle~q ;
wire \Selector4~0_combout ;
wire \sig_dgwb_state.s_wait_admin~q ;
wire \Selector8~0_combout ;
wire \sig_dgwb_state.s_write_mtp~q ;
wire \Selector7~0_combout ;
wire \sig_dgwb_state.s_write_zeros~q ;
wire \sig_addr_cmd[0].addr[4]~3_combout ;
wire \generate_wdata~q ;
wire \ac_write_block:sig_count[3]~2_combout ;
wire \ac_write_block:sig_count[3]~3_combout ;
wire \ac_write_block:sig_count[3]~1_combout ;
wire \ac_write_block:sig_count[0]~q ;
wire \Add1~2 ;
wire \Add1~5_sumout ;
wire \ac_write_block:sig_count[1]~q ;
wire \Add1~6 ;
wire \Add1~9_sumout ;
wire \ac_write_block:sig_count[2]~q ;
wire \Add1~10 ;
wire \Add1~13_sumout ;
wire \ac_write_block:sig_count[3]~q ;
wire \Add1~14 ;
wire \Add1~17_sumout ;
wire \ac_write_block:sig_count[4]~q ;
wire \ac_write_block:sig_count[3]~0_combout ;
wire \Add1~18 ;
wire \Add1~21_sumout ;
wire \ac_write_block:sig_count[5]~q ;
wire \Add1~22 ;
wire \Add1~25_sumout ;
wire \ac_write_block:sig_count[6]~q ;
wire \Add1~26 ;
wire \Add1~29_sumout ;
wire \ac_write_block:sig_count[7]~q ;
wire \Selector91~0_combout ;
wire \Selector32~0_combout ;
wire \Selector91~1_combout ;
wire \access_complete~q ;
wire \Selector11~10_combout ;
wire \sig_dgwb_state.s_write_0011_step~q ;
wire \Equal1~0_combout ;
wire \Selector26~0_combout ;
wire \Selector26~1_combout ;
wire \sig_addr_cmd[0].addr[4]~0_combout ;
wire \sig_addr_cmd[0].addr[4]~1_combout ;
wire \sig_addr_cmd[0].addr[4]~4_combout ;
wire \sig_addr_cmd[0].addr[4]~5_combout ;
wire \sig_addr_cmd[0].addr[4]~2_combout ;
wire \sig_addr_cmd~0_combout ;
wire \Selector25~0_combout ;
wire \Selector24~0_combout ;
wire \Selector23~0_combout ;
wire \sig_dgwb_last_state.s_release_admin~q ;
wire \ac_handshake_proc~2_combout ;
wire \dgwb_dqs_burst~0_combout ;
wire \ac_handshake_proc~3_combout ;
wire \Selector50~0_combout ;
wire \Selector50~1_combout ;
wire \Selector50~2_combout ;
wire \sig_addr_cmd[0].addr[12]~0_combout ;
wire \Selector58~0_combout ;
wire \Selector74~0_combout ;
wire \WideOr4~0_combout ;
wire \Selector66~0_combout ;
wire \WideOr7~0_combout ;
wire \Selector82~0_combout ;
wire \Selector57~0_combout ;
wire \Selector73~0_combout ;
wire \Selector65~0_combout ;
wire \Selector81~0_combout ;
wire \Selector56~0_combout ;
wire \Selector72~0_combout ;
wire \Selector64~0_combout ;
wire \Selector80~0_combout ;
wire \Selector55~0_combout ;
wire \Selector71~0_combout ;
wire \Selector63~0_combout ;
wire \Selector79~0_combout ;
wire \Selector54~0_combout ;
wire \Selector70~0_combout ;
wire \Selector62~0_combout ;
wire \Selector78~0_combout ;
wire \Selector53~0_combout ;
wire \Selector69~0_combout ;
wire \Selector61~0_combout ;
wire \Selector77~0_combout ;
wire \Selector52~0_combout ;
wire \Selector68~0_combout ;
wire \Selector60~0_combout ;
wire \Selector76~0_combout ;
wire \Selector51~0_combout ;
wire \Selector67~0_combout ;
wire \Selector59~0_combout ;
wire \Selector75~0_combout ;
wire \sig_dgwb_last_state.s_idle~q ;
wire \ac_handshake_proc~4_combout ;


dffeas \sig_addr_cmd[0].addr[2] (
	.clk(clk),
	.d(\Selector26~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_dgwb_state.s_write_wlat~q ),
	.sload(\sig_dgwb_state.s_write_1100_step~q ),
	.ena(\sig_addr_cmd[0].addr[4]~2_combout ),
	.q(sig_addr_cmd0addr2),
	.prn(vcc));
defparam \sig_addr_cmd[0].addr[2] .is_wysiwyg = "true";
defparam \sig_addr_cmd[0].addr[2] .power_up = "low";

dffeas \sig_addr_cmd[0].addr[3] (
	.clk(clk),
	.d(\Selector25~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\sig_dgwb_state.s_write_wlat~q ),
	.sload(\sig_dgwb_state.s_write_1100_step~q ),
	.ena(\sig_addr_cmd[0].addr[4]~2_combout ),
	.q(sig_addr_cmd0addr3),
	.prn(vcc));
defparam \sig_addr_cmd[0].addr[3] .is_wysiwyg = "true";
defparam \sig_addr_cmd[0].addr[3] .power_up = "low";

dffeas \sig_addr_cmd[0].addr[4] (
	.clk(clk),
	.d(\Selector24~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sig_dgwb_state.s_write_wlat~q ),
	.ena(\sig_addr_cmd[0].addr[4]~2_combout ),
	.q(sig_addr_cmd0addr4),
	.prn(vcc));
defparam \sig_addr_cmd[0].addr[4] .is_wysiwyg = "true";
defparam \sig_addr_cmd[0].addr[4] .power_up = "low";

dffeas \sig_addr_cmd[0].addr[5] (
	.clk(clk),
	.d(\Selector23~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sig_dgwb_state.s_write_wlat~q ),
	.ena(\sig_addr_cmd[0].addr[4]~2_combout ),
	.q(sig_addr_cmd0addr5),
	.prn(vcc));
defparam \sig_addr_cmd[0].addr[5] .is_wysiwyg = "true";
defparam \sig_addr_cmd[0].addr[5] .power_up = "low";

dffeas \sig_addr_cmd[0].cas_n (
	.clk(clk),
	.d(\Selector32~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sig_dgwb_state.s_write_wlat~q ),
	.ena(\sig_addr_cmd[0].addr[4]~2_combout ),
	.q(sig_addr_cmd0cas_n),
	.prn(vcc));
defparam \sig_addr_cmd[0].cas_n .is_wysiwyg = "true";
defparam \sig_addr_cmd[0].cas_n .power_up = "low";

dffeas \dgwb_ctrl.command_done (
	.clk(clk),
	.d(\ac_handshake_proc~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_ctrlcommand_done),
	.prn(vcc));
defparam \dgwb_ctrl.command_done .is_wysiwyg = "true";
defparam \dgwb_ctrl.command_done .power_up = "low";

dffeas dgwb_wdp_ovride(
	.clk(clk),
	.d(\dgwb_dqs_burst~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdp_ovride1),
	.prn(vcc));
defparam dgwb_wdp_ovride.is_wysiwyg = "true";
defparam dgwb_wdp_ovride.power_up = "low";

dffeas \sig_addr_cmd[0].cke[0] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sig_addr_cmd0cke0),
	.prn(vcc));
defparam \sig_addr_cmd[0].cke[0] .is_wysiwyg = "true";
defparam \sig_addr_cmd[0].cke[0] .power_up = "low";

dffeas dgwb_ac_access_req(
	.clk(clk),
	.d(\ac_handshake_proc~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_ac_access_req1),
	.prn(vcc));
defparam dgwb_ac_access_req.is_wysiwyg = "true";
defparam dgwb_ac_access_req.power_up = "low";

dffeas \sig_addr_cmd[1].cs_n[0] (
	.clk(clk),
	.d(\Selector50~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sig_addr_cmd1cs_n0),
	.prn(vcc));
defparam \sig_addr_cmd[1].cs_n[0] .is_wysiwyg = "true";
defparam \sig_addr_cmd[1].cs_n[0] .power_up = "low";

dffeas \sig_addr_cmd[0].addr[12] (
	.clk(clk),
	.d(\sig_addr_cmd[0].addr[12]~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sig_addr_cmd0addr12),
	.prn(vcc));
defparam \sig_addr_cmd[0].addr[12] .is_wysiwyg = "true";
defparam \sig_addr_cmd[0].addr[12] .power_up = "low";

dffeas \sig_addr_cmd[0].rst_n (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sig_addr_cmd0rst_n),
	.prn(vcc));
defparam \sig_addr_cmd[0].rst_n .is_wysiwyg = "true";
defparam \sig_addr_cmd[0].rst_n .power_up = "low";

dffeas \dgwb_wdata[120] (
	.clk(clk),
	.d(\Selector58~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_120),
	.prn(vcc));
defparam \dgwb_wdata[120] .is_wysiwyg = "true";
defparam \dgwb_wdata[120] .power_up = "low";

dffeas \dgwb_wdata[56] (
	.clk(clk),
	.d(\Selector74~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_56),
	.prn(vcc));
defparam \dgwb_wdata[56] .is_wysiwyg = "true";
defparam \dgwb_wdata[56] .power_up = "low";

dffeas \dgwb_wdata[88] (
	.clk(clk),
	.d(\Selector66~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_88),
	.prn(vcc));
defparam \dgwb_wdata[88] .is_wysiwyg = "true";
defparam \dgwb_wdata[88] .power_up = "low";

dffeas \dgwb_wdata[24] (
	.clk(clk),
	.d(\Selector82~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_24),
	.prn(vcc));
defparam \dgwb_wdata[24] .is_wysiwyg = "true";
defparam \dgwb_wdata[24] .power_up = "low";

dffeas \dgwb_wdata[121] (
	.clk(clk),
	.d(\Selector57~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_121),
	.prn(vcc));
defparam \dgwb_wdata[121] .is_wysiwyg = "true";
defparam \dgwb_wdata[121] .power_up = "low";

dffeas \dgwb_wdata[57] (
	.clk(clk),
	.d(\Selector73~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_57),
	.prn(vcc));
defparam \dgwb_wdata[57] .is_wysiwyg = "true";
defparam \dgwb_wdata[57] .power_up = "low";

dffeas \dgwb_wdata[89] (
	.clk(clk),
	.d(\Selector65~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_89),
	.prn(vcc));
defparam \dgwb_wdata[89] .is_wysiwyg = "true";
defparam \dgwb_wdata[89] .power_up = "low";

dffeas \dgwb_wdata[25] (
	.clk(clk),
	.d(\Selector81~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_25),
	.prn(vcc));
defparam \dgwb_wdata[25] .is_wysiwyg = "true";
defparam \dgwb_wdata[25] .power_up = "low";

dffeas \dgwb_wdata[122] (
	.clk(clk),
	.d(\Selector56~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_122),
	.prn(vcc));
defparam \dgwb_wdata[122] .is_wysiwyg = "true";
defparam \dgwb_wdata[122] .power_up = "low";

dffeas \dgwb_wdata[58] (
	.clk(clk),
	.d(\Selector72~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_58),
	.prn(vcc));
defparam \dgwb_wdata[58] .is_wysiwyg = "true";
defparam \dgwb_wdata[58] .power_up = "low";

dffeas \dgwb_wdata[90] (
	.clk(clk),
	.d(\Selector64~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_90),
	.prn(vcc));
defparam \dgwb_wdata[90] .is_wysiwyg = "true";
defparam \dgwb_wdata[90] .power_up = "low";

dffeas \dgwb_wdata[26] (
	.clk(clk),
	.d(\Selector80~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_26),
	.prn(vcc));
defparam \dgwb_wdata[26] .is_wysiwyg = "true";
defparam \dgwb_wdata[26] .power_up = "low";

dffeas \dgwb_wdata[123] (
	.clk(clk),
	.d(\Selector55~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_123),
	.prn(vcc));
defparam \dgwb_wdata[123] .is_wysiwyg = "true";
defparam \dgwb_wdata[123] .power_up = "low";

dffeas \dgwb_wdata[59] (
	.clk(clk),
	.d(\Selector71~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_59),
	.prn(vcc));
defparam \dgwb_wdata[59] .is_wysiwyg = "true";
defparam \dgwb_wdata[59] .power_up = "low";

dffeas \dgwb_wdata[91] (
	.clk(clk),
	.d(\Selector63~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_91),
	.prn(vcc));
defparam \dgwb_wdata[91] .is_wysiwyg = "true";
defparam \dgwb_wdata[91] .power_up = "low";

dffeas \dgwb_wdata[27] (
	.clk(clk),
	.d(\Selector79~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_27),
	.prn(vcc));
defparam \dgwb_wdata[27] .is_wysiwyg = "true";
defparam \dgwb_wdata[27] .power_up = "low";

dffeas \dgwb_wdata[124] (
	.clk(clk),
	.d(\Selector54~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_124),
	.prn(vcc));
defparam \dgwb_wdata[124] .is_wysiwyg = "true";
defparam \dgwb_wdata[124] .power_up = "low";

dffeas \dgwb_wdata[60] (
	.clk(clk),
	.d(\Selector70~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_60),
	.prn(vcc));
defparam \dgwb_wdata[60] .is_wysiwyg = "true";
defparam \dgwb_wdata[60] .power_up = "low";

dffeas \dgwb_wdata[92] (
	.clk(clk),
	.d(\Selector62~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_92),
	.prn(vcc));
defparam \dgwb_wdata[92] .is_wysiwyg = "true";
defparam \dgwb_wdata[92] .power_up = "low";

dffeas \dgwb_wdata[28] (
	.clk(clk),
	.d(\Selector78~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_28),
	.prn(vcc));
defparam \dgwb_wdata[28] .is_wysiwyg = "true";
defparam \dgwb_wdata[28] .power_up = "low";

dffeas \dgwb_wdata[125] (
	.clk(clk),
	.d(\Selector53~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_125),
	.prn(vcc));
defparam \dgwb_wdata[125] .is_wysiwyg = "true";
defparam \dgwb_wdata[125] .power_up = "low";

dffeas \dgwb_wdata[61] (
	.clk(clk),
	.d(\Selector69~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_61),
	.prn(vcc));
defparam \dgwb_wdata[61] .is_wysiwyg = "true";
defparam \dgwb_wdata[61] .power_up = "low";

dffeas \dgwb_wdata[93] (
	.clk(clk),
	.d(\Selector61~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_93),
	.prn(vcc));
defparam \dgwb_wdata[93] .is_wysiwyg = "true";
defparam \dgwb_wdata[93] .power_up = "low";

dffeas \dgwb_wdata[29] (
	.clk(clk),
	.d(\Selector77~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_29),
	.prn(vcc));
defparam \dgwb_wdata[29] .is_wysiwyg = "true";
defparam \dgwb_wdata[29] .power_up = "low";

dffeas \dgwb_wdata[126] (
	.clk(clk),
	.d(\Selector52~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_126),
	.prn(vcc));
defparam \dgwb_wdata[126] .is_wysiwyg = "true";
defparam \dgwb_wdata[126] .power_up = "low";

dffeas \dgwb_wdata[62] (
	.clk(clk),
	.d(\Selector68~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_62),
	.prn(vcc));
defparam \dgwb_wdata[62] .is_wysiwyg = "true";
defparam \dgwb_wdata[62] .power_up = "low";

dffeas \dgwb_wdata[94] (
	.clk(clk),
	.d(\Selector60~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_94),
	.prn(vcc));
defparam \dgwb_wdata[94] .is_wysiwyg = "true";
defparam \dgwb_wdata[94] .power_up = "low";

dffeas \dgwb_wdata[30] (
	.clk(clk),
	.d(\Selector76~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_30),
	.prn(vcc));
defparam \dgwb_wdata[30] .is_wysiwyg = "true";
defparam \dgwb_wdata[30] .power_up = "low";

dffeas \dgwb_wdata[127] (
	.clk(clk),
	.d(\Selector51~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_127),
	.prn(vcc));
defparam \dgwb_wdata[127] .is_wysiwyg = "true";
defparam \dgwb_wdata[127] .power_up = "low";

dffeas \dgwb_wdata[63] (
	.clk(clk),
	.d(\Selector67~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_63),
	.prn(vcc));
defparam \dgwb_wdata[63] .is_wysiwyg = "true";
defparam \dgwb_wdata[63] .power_up = "low";

dffeas \dgwb_wdata[95] (
	.clk(clk),
	.d(\Selector59~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_95),
	.prn(vcc));
defparam \dgwb_wdata[95] .is_wysiwyg = "true";
defparam \dgwb_wdata[95] .power_up = "low";

dffeas \dgwb_wdata[31] (
	.clk(clk),
	.d(\Selector75~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_wdata_31),
	.prn(vcc));
defparam \dgwb_wdata[31] .is_wysiwyg = "true";
defparam \dgwb_wdata[31] .power_up = "low";

dffeas \dgwb_ctrl.command_ack (
	.clk(clk),
	.d(\ac_handshake_proc~4_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dgwb_ctrlcommand_ack),
	.prn(vcc));
defparam \dgwb_ctrl.command_ack .is_wysiwyg = "true";
defparam \dgwb_ctrl.command_ack .power_up = "low";

arriaii_lcell_comb \dgwb_wdp_ovride~_wirecell (
	.dataa(!dgwb_wdp_ovride1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(dgwb_wdp_ovride2),
	.sumout(),
	.cout(),
	.shareout());
defparam \dgwb_wdp_ovride~_wirecell .extended_lut = "off";
defparam \dgwb_wdp_ovride~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dgwb_wdp_ovride~_wirecell .shared_arith = "off";

arriaii_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\ac_write_block:sig_count[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(\Add1~2 ),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h00000000000000FF;
defparam \Add1~1 .shared_arith = "off";

dffeas \sig_dgwb_last_state.s_write_01_pairs (
	.clk(clk),
	.d(\sig_dgwb_state.s_write_01_pairs~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_last_state.s_write_01_pairs~q ),
	.prn(vcc));
defparam \sig_dgwb_last_state.s_write_01_pairs .is_wysiwyg = "true";
defparam \sig_dgwb_last_state.s_write_01_pairs .power_up = "low";

arriaii_lcell_comb \Selector9~4 (
	.dataa(!\sig_dgwb_state.s_write_mtp~q ),
	.datab(!\access_complete~q ),
	.datac(!\sig_dgwb_last_state.s_write_01_pairs~q ),
	.datad(!\sig_dgwb_state.s_write_01_pairs~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector9~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector9~4 .extended_lut = "off";
defparam \Selector9~4 .lut_mask = 64'h55FD55FD55FD55FD;
defparam \Selector9~4 .shared_arith = "off";

dffeas \sig_dgwb_state.s_write_01_pairs (
	.clk(clk),
	.d(\Selector9~4_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_state.s_write_01_pairs~q ),
	.prn(vcc));
defparam \sig_dgwb_state.s_write_01_pairs .is_wysiwyg = "true";
defparam \sig_dgwb_state.s_write_01_pairs .power_up = "low";

arriaii_lcell_comb \Selector11~5 (
	.dataa(!\sig_dgwb_last_state.s_write_01_pairs~q ),
	.datab(!\sig_dgwb_state.s_write_01_pairs~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector11~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector11~5 .extended_lut = "off";
defparam \Selector11~5 .lut_mask = 64'h1111111111111111;
defparam \Selector11~5 .shared_arith = "off";

dffeas \sig_dgwb_last_state.s_write_1100_step (
	.clk(clk),
	.d(\sig_dgwb_state.s_write_1100_step~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_last_state.s_write_1100_step~q ),
	.prn(vcc));
defparam \sig_dgwb_last_state.s_write_1100_step .is_wysiwyg = "true";
defparam \sig_dgwb_last_state.s_write_1100_step .power_up = "low";

arriaii_lcell_comb \Selector10~0 (
	.dataa(!\Selector11~4_combout ),
	.datab(!\access_complete~q ),
	.datac(!\Selector11~5_combout ),
	.datad(!\sig_dgwb_state.s_write_1100_step~q ),
	.datae(!\sig_dgwb_last_state.s_write_1100_step~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector10~0 .extended_lut = "off";
defparam \Selector10~0 .lut_mask = 64'h0155014401550144;
defparam \Selector10~0 .shared_arith = "off";

dffeas \sig_dgwb_state.s_write_1100_step (
	.clk(clk),
	.d(\Selector10~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_state.s_write_1100_step~q ),
	.prn(vcc));
defparam \sig_dgwb_state.s_write_1100_step .is_wysiwyg = "true";
defparam \sig_dgwb_state.s_write_1100_step .power_up = "low";

arriaii_lcell_comb \Selector11~6 (
	.dataa(!\access_complete~q ),
	.datab(!\sig_dgwb_state.s_write_1100_step~q ),
	.datac(!\sig_dgwb_last_state.s_write_1100_step~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector11~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector11~6 .extended_lut = "off";
defparam \Selector11~6 .lut_mask = 64'h0101010101010101;
defparam \Selector11~6 .shared_arith = "off";

arriaii_lcell_comb \Selector6~0 (
	.dataa(!\Selector11~4_combout ),
	.datab(!\access_complete~q ),
	.datac(!\Selector11~5_combout ),
	.datad(!\Selector11~6_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~0 .extended_lut = "off";
defparam \Selector6~0 .lut_mask = 64'h5400540054005400;
defparam \Selector6~0 .shared_arith = "off";

arriaii_lcell_comb \Selector6~1 (
	.dataa(!\sig_dgwb_last_state.s_write_zeros~q ),
	.datab(!\sig_dgwb_state.s_write_zeros~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector6~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~1 .extended_lut = "off";
defparam \Selector6~1 .lut_mask = 64'h1111111111111111;
defparam \Selector6~1 .shared_arith = "off";

arriaii_lcell_comb \Selector6~2 (
	.dataa(!\access_complete~q ),
	.datab(!\sig_dgwb_state.s_write_ones~q ),
	.datac(!\sig_dgwb_last_state.s_write_ones~q ),
	.datad(!\Selector6~0_combout ),
	.datae(!\Selector6~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector6~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~2 .extended_lut = "off";
defparam \Selector6~2 .lut_mask = 64'h0032007700320077;
defparam \Selector6~2 .shared_arith = "off";

dffeas \sig_dgwb_state.s_write_ones (
	.clk(clk),
	.d(\Selector6~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_state.s_write_ones~q ),
	.prn(vcc));
defparam \sig_dgwb_state.s_write_ones .is_wysiwyg = "true";
defparam \sig_dgwb_state.s_write_ones .power_up = "low";

dffeas \sig_dgwb_last_state.s_write_ones (
	.clk(clk),
	.d(\sig_dgwb_state.s_write_ones~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_last_state.s_write_ones~q ),
	.prn(vcc));
defparam \sig_dgwb_last_state.s_write_ones .is_wysiwyg = "true";
defparam \sig_dgwb_last_state.s_write_ones .power_up = "low";

arriaii_lcell_comb \Selector5~2 (
	.dataa(!dgb_ac_access_gnt_r),
	.datab(!curr_cmdcmd_write_btp),
	.datac(!\sig_dgwb_state.s_wait_admin~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~2 .extended_lut = "off";
defparam \Selector5~2 .lut_mask = 64'h0101010101010101;
defparam \Selector5~2 .shared_arith = "off";

dffeas \sig_dgwb_state.s_write_btp (
	.clk(clk),
	.d(\Selector5~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_state.s_write_btp~q ),
	.prn(vcc));
defparam \sig_dgwb_state.s_write_btp .is_wysiwyg = "true";
defparam \sig_dgwb_state.s_write_btp .power_up = "low";

dffeas \sig_dgwb_last_state.s_write_0011_step (
	.clk(clk),
	.d(\sig_dgwb_state.s_write_0011_step~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_last_state.s_write_0011_step~q ),
	.prn(vcc));
defparam \sig_dgwb_last_state.s_write_0011_step .is_wysiwyg = "true";
defparam \sig_dgwb_last_state.s_write_0011_step .power_up = "low";

arriaii_lcell_comb \Selector5~3 (
	.dataa(!dgb_ac_access_gnt_r),
	.datab(!\sig_dgwb_state.s_release_admin~q ),
	.datac(!\access_complete~q ),
	.datad(!\sig_dgwb_last_state.s_write_0011_step~q ),
	.datae(!\sig_dgwb_state.s_write_0011_step~q ),
	.dataf(!\sig_dgwb_last_state.s_write_wlat~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~3 .extended_lut = "off";
defparam \Selector5~3 .lut_mask = 64'h2222000F2E2E000F;
defparam \Selector5~3 .shared_arith = "off";

arriaii_lcell_comb \Selector5~4 (
	.dataa(!\access_complete~q ),
	.datab(!\sig_dgwb_last_state.s_write_01_pairs~q ),
	.datac(!\sig_dgwb_state.s_write_01_pairs~q ),
	.datad(!\sig_dgwb_state.s_write_1100_step~q ),
	.datae(!\sig_dgwb_last_state.s_write_1100_step~q ),
	.dataf(!\Selector5~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~4 .extended_lut = "off";
defparam \Selector5~4 .lut_mask = 64'h01010151F101F151;
defparam \Selector5~4 .shared_arith = "off";

dffeas \sig_dgwb_last_state.s_write_zeros (
	.clk(clk),
	.d(\sig_dgwb_state.s_write_zeros~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_last_state.s_write_zeros~q ),
	.prn(vcc));
defparam \sig_dgwb_last_state.s_write_zeros .is_wysiwyg = "true";
defparam \sig_dgwb_last_state.s_write_zeros .power_up = "low";

arriaii_lcell_comb \Selector5~5 (
	.dataa(!\sig_dgwb_state.s_write_ones~q ),
	.datab(!\sig_dgwb_last_state.s_write_ones~q ),
	.datac(!\sig_dgwb_last_state.s_write_zeros~q ),
	.datad(!\sig_dgwb_state.s_write_zeros~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~5 .extended_lut = "off";
defparam \Selector5~5 .lut_mask = 64'h110F110F110F110F;
defparam \Selector5~5 .shared_arith = "off";

arriaii_lcell_comb \Selector5~6 (
	.dataa(!curr_ctrlcommand_ack),
	.datab(!\sig_dgwb_state.s_idle~q ),
	.datac(!ac_muxctrl_broadcast_rcommand_req),
	.datad(!\access_complete~q ),
	.datae(!\Selector5~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~6 .extended_lut = "off";
defparam \Selector5~6 .lut_mask = 64'h0808083B0808083B;
defparam \Selector5~6 .shared_arith = "off";

arriaii_lcell_comb \Selector5~7 (
	.dataa(!\sig_dgwb_state.s_idle~q ),
	.datab(!\sig_dgwb_state.s_write_ones~q ),
	.datac(!\sig_dgwb_state.s_write_zeros~q ),
	.datad(!\Selector5~4_combout ),
	.datae(!\Selector5~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~7 .extended_lut = "off";
defparam \Selector5~7 .lut_mask = 64'h0040FFFF0040FFFF;
defparam \Selector5~7 .shared_arith = "off";

arriaii_lcell_comb \Selector12~0 (
	.dataa(!\sig_dgwb_state.s_write_wlat~q ),
	.datab(!curr_cmdcmd_was),
	.datac(!dgb_ac_access_gnt_r),
	.datad(!\sig_dgwb_state.s_write_mtp~q ),
	.datae(!\sig_dgwb_state.s_wait_admin~q ),
	.dataf(!\sig_dgwb_state.s_write_btp~q ),
	.datag(!\Selector5~7_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector12~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector12~0 .extended_lut = "on";
defparam \Selector12~0 .lut_mask = 64'h5000030000000000;
defparam \Selector12~0 .shared_arith = "off";

dffeas \sig_dgwb_state.s_write_wlat (
	.clk(clk),
	.d(\Selector12~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_state.s_write_wlat~q ),
	.prn(vcc));
defparam \sig_dgwb_state.s_write_wlat .is_wysiwyg = "true";
defparam \sig_dgwb_state.s_write_wlat .power_up = "low";

dffeas \sig_dgwb_last_state.s_write_wlat (
	.clk(clk),
	.d(\sig_dgwb_state.s_write_wlat~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_last_state.s_write_wlat~q ),
	.prn(vcc));
defparam \sig_dgwb_last_state.s_write_wlat .is_wysiwyg = "true";
defparam \sig_dgwb_last_state.s_write_wlat .power_up = "low";

arriaii_lcell_comb \Selector11~11 (
	.dataa(!\sig_dgwb_state.s_write_0011_step~q ),
	.datab(!\sig_dgwb_last_state.s_write_ones~q ),
	.datac(!\sig_dgwb_last_state.s_write_wlat~q ),
	.datad(!\sig_dgwb_state.s_write_ones~q ),
	.datae(!\sig_dgwb_state.s_write_wlat~q ),
	.dataf(!\access_complete~q ),
	.datag(!\sig_dgwb_last_state.s_write_0011_step~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector11~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector11~11 .extended_lut = "on";
defparam \Selector11~11 .lut_mask = 64'h0000000005330F33;
defparam \Selector11~11 .shared_arith = "off";

arriaii_lcell_comb \Selector11~7 (
	.dataa(!\sig_dgwb_state.s_write_btp~q ),
	.datab(!\sig_dgwb_state.s_write_mtp~q ),
	.datac(!\access_complete~q ),
	.datad(!\sig_dgwb_last_state.s_write_zeros~q ),
	.datae(!\sig_dgwb_state.s_write_zeros~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector11~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector11~7 .extended_lut = "off";
defparam \Selector11~7 .lut_mask = 64'h8888888088888880;
defparam \Selector11~7 .shared_arith = "off";

arriaii_lcell_comb \Selector11~8 (
	.dataa(!dgb_ac_access_gnt_r),
	.datab(!curr_ctrlcommand_ack),
	.datac(!\sig_dgwb_state.s_idle~q ),
	.datad(!ac_muxctrl_broadcast_rcommand_req),
	.datae(!\sig_dgwb_state.s_wait_admin~q ),
	.dataf(!\Selector11~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector11~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector11~8 .extended_lut = "off";
defparam \Selector11~8 .lut_mask = 64'h00000000FF3F1111;
defparam \Selector11~8 .shared_arith = "off";

arriaii_lcell_comb \Selector11~9 (
	.dataa(!\Selector11~11_combout ),
	.datab(!\Selector6~0_combout ),
	.datac(!\Selector11~8_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector11~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector11~9 .extended_lut = "off";
defparam \Selector11~9 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \Selector11~9 .shared_arith = "off";

dffeas \sig_dgwb_state.s_release_admin (
	.clk(clk),
	.d(\Selector11~11_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector11~9_combout ),
	.q(\sig_dgwb_state.s_release_admin~q ),
	.prn(vcc));
defparam \sig_dgwb_state.s_release_admin .is_wysiwyg = "true";
defparam \sig_dgwb_state.s_release_admin .power_up = "low";

arriaii_lcell_comb \Selector11~4 (
	.dataa(!dgb_ac_access_gnt_r),
	.datab(!\sig_dgwb_state.s_release_admin~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector11~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector11~4 .extended_lut = "off";
defparam \Selector11~4 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \Selector11~4 .shared_arith = "off";

dffeas \sig_dgwb_state.s_idle (
	.clk(clk),
	.d(\Selector11~4_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Selector11~9_combout ),
	.q(\sig_dgwb_state.s_idle~q ),
	.prn(vcc));
defparam \sig_dgwb_state.s_idle .is_wysiwyg = "true";
defparam \sig_dgwb_state.s_idle .power_up = "low";

arriaii_lcell_comb \Selector4~0 (
	.dataa(!dgb_ac_access_gnt_r),
	.datab(!curr_ctrlcommand_ack),
	.datac(!\sig_dgwb_state.s_idle~q ),
	.datad(!ac_muxctrl_broadcast_rcommand_req),
	.datae(!\sig_dgwb_state.s_wait_admin~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~0 .extended_lut = "off";
defparam \Selector4~0 .lut_mask = 64'h00C0BBFB00C0BBFB;
defparam \Selector4~0 .shared_arith = "off";

dffeas \sig_dgwb_state.s_wait_admin (
	.clk(clk),
	.d(\Selector4~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_state.s_wait_admin~q ),
	.prn(vcc));
defparam \sig_dgwb_state.s_wait_admin .is_wysiwyg = "true";
defparam \sig_dgwb_state.s_wait_admin .power_up = "low";

arriaii_lcell_comb \Selector8~0 (
	.dataa(!dgb_ac_access_gnt_r),
	.datab(!curr_cmdcmd_write_mtp),
	.datac(!\sig_dgwb_state.s_wait_admin~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector8~0 .extended_lut = "off";
defparam \Selector8~0 .lut_mask = 64'h0101010101010101;
defparam \Selector8~0 .shared_arith = "off";

dffeas \sig_dgwb_state.s_write_mtp (
	.clk(clk),
	.d(\Selector8~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_state.s_write_mtp~q ),
	.prn(vcc));
defparam \sig_dgwb_state.s_write_mtp .is_wysiwyg = "true";
defparam \sig_dgwb_state.s_write_mtp .power_up = "low";

arriaii_lcell_comb \Selector7~0 (
	.dataa(!\sig_dgwb_state.s_write_btp~q ),
	.datab(!\sig_dgwb_state.s_write_mtp~q ),
	.datac(!\access_complete~q ),
	.datad(!\sig_dgwb_last_state.s_write_zeros~q ),
	.datae(!\sig_dgwb_state.s_write_zeros~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector7~0 .extended_lut = "off";
defparam \Selector7~0 .lut_mask = 64'h4444CCC44444CCC4;
defparam \Selector7~0 .shared_arith = "off";

dffeas \sig_dgwb_state.s_write_zeros (
	.clk(clk),
	.d(\Selector7~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_state.s_write_zeros~q ),
	.prn(vcc));
defparam \sig_dgwb_state.s_write_zeros .is_wysiwyg = "true";
defparam \sig_dgwb_state.s_write_zeros .power_up = "low";

arriaii_lcell_comb \sig_addr_cmd[0].addr[4]~3 (
	.dataa(!\sig_dgwb_state.s_write_wlat~q ),
	.datab(!\sig_dgwb_last_state.s_write_wlat~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_addr_cmd[0].addr[4]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_addr_cmd[0].addr[4]~3 .extended_lut = "off";
defparam \sig_addr_cmd[0].addr[4]~3 .lut_mask = 64'h1111111111111111;
defparam \sig_addr_cmd[0].addr[4]~3 .shared_arith = "off";

dffeas generate_wdata(
	.clk(clk),
	.d(\sig_addr_cmd[0].addr[4]~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\generate_wdata~q ),
	.prn(vcc));
defparam generate_wdata.is_wysiwyg = "true";
defparam generate_wdata.power_up = "low";

arriaii_lcell_comb \ac_write_block:sig_count[3]~2 (
	.dataa(!\sig_dgwb_last_state.s_write_zeros~q ),
	.datab(!\sig_dgwb_state.s_write_zeros~q ),
	.datac(!\sig_dgwb_last_state.s_write_0011_step~q ),
	.datad(!\sig_dgwb_state.s_write_01_pairs~q ),
	.datae(!\sig_dgwb_state.s_write_1100_step~q ),
	.dataf(!\sig_dgwb_last_state.s_write_1100_step~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_write_block:sig_count[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_write_block:sig_count[3]~2 .extended_lut = "off";
defparam \ac_write_block:sig_count[3]~2 .lut_mask = 64'h1D1111111D11DD11;
defparam \ac_write_block:sig_count[3]~2 .shared_arith = "off";

arriaii_lcell_comb \ac_write_block:sig_count[3]~3 (
	.dataa(!\sig_dgwb_last_state.s_write_ones~q ),
	.datab(!\sig_dgwb_state.s_write_zeros~q ),
	.datac(!\generate_wdata~q ),
	.datad(!\ac_write_block:sig_count[3]~2_combout ),
	.datae(!\sig_dgwb_state.s_write_wlat~q ),
	.dataf(!\Selector11~5_combout ),
	.datag(!\sig_dgwb_state.s_write_ones~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_write_block:sig_count[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_write_block:sig_count[3]~3 .extended_lut = "on";
defparam \ac_write_block:sig_count[3]~3 .lut_mask = 64'h05F50F0FC5F50F0F;
defparam \ac_write_block:sig_count[3]~3 .shared_arith = "off";

arriaii_lcell_comb \ac_write_block:sig_count[3]~1 (
	.dataa(!\dgwb_dqs_burst~0_combout ),
	.datab(!\sig_addr_cmd[0].addr[4]~3_combout ),
	.datac(!\generate_wdata~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_write_block:sig_count[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_write_block:sig_count[3]~1 .extended_lut = "off";
defparam \ac_write_block:sig_count[3]~1 .lut_mask = 64'h4545454545454545;
defparam \ac_write_block:sig_count[3]~1 .shared_arith = "off";

dffeas \ac_write_block:sig_count[0] (
	.clk(clk),
	.d(\Add1~1_sumout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\ac_write_block:sig_count[3]~3_combout ),
	.sload(gnd),
	.ena(\ac_write_block:sig_count[3]~1_combout ),
	.q(\ac_write_block:sig_count[0]~q ),
	.prn(vcc));
defparam \ac_write_block:sig_count[0] .is_wysiwyg = "true";
defparam \ac_write_block:sig_count[0] .power_up = "low";

arriaii_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\ac_write_block:sig_count[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~5 .shared_arith = "off";

dffeas \ac_write_block:sig_count[1] (
	.clk(clk),
	.d(\Add1~5_sumout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\ac_write_block:sig_count[3]~3_combout ),
	.sload(gnd),
	.ena(\ac_write_block:sig_count[3]~1_combout ),
	.q(\ac_write_block:sig_count[1]~q ),
	.prn(vcc));
defparam \ac_write_block:sig_count[1] .is_wysiwyg = "true";
defparam \ac_write_block:sig_count[1] .power_up = "low";

arriaii_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\ac_write_block:sig_count[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~9 .shared_arith = "off";

dffeas \ac_write_block:sig_count[2] (
	.clk(clk),
	.d(\Add1~9_sumout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\ac_write_block:sig_count[3]~3_combout ),
	.sload(gnd),
	.ena(\ac_write_block:sig_count[3]~1_combout ),
	.q(\ac_write_block:sig_count[2]~q ),
	.prn(vcc));
defparam \ac_write_block:sig_count[2] .is_wysiwyg = "true";
defparam \ac_write_block:sig_count[2] .power_up = "low";

arriaii_lcell_comb \Add1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\ac_write_block:sig_count[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~13 .shared_arith = "off";

dffeas \ac_write_block:sig_count[3] (
	.clk(clk),
	.d(\Add1~13_sumout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\ac_write_block:sig_count[3]~3_combout ),
	.sload(gnd),
	.ena(\ac_write_block:sig_count[3]~1_combout ),
	.q(\ac_write_block:sig_count[3]~q ),
	.prn(vcc));
defparam \ac_write_block:sig_count[3] .is_wysiwyg = "true";
defparam \ac_write_block:sig_count[3] .power_up = "low";

arriaii_lcell_comb \Add1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\ac_write_block:sig_count[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~17 .shared_arith = "off";

dffeas \ac_write_block:sig_count[4] (
	.clk(clk),
	.d(\Add1~17_sumout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\ac_write_block:sig_count[3]~3_combout ),
	.sload(gnd),
	.ena(\ac_write_block:sig_count[3]~1_combout ),
	.q(\ac_write_block:sig_count[4]~q ),
	.prn(vcc));
defparam \ac_write_block:sig_count[4] .is_wysiwyg = "true";
defparam \ac_write_block:sig_count[4] .power_up = "low";

arriaii_lcell_comb \ac_write_block:sig_count[3]~0 (
	.dataa(!\sig_dgwb_state.s_write_wlat~q ),
	.datab(!\generate_wdata~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_write_block:sig_count[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_write_block:sig_count[3]~0 .extended_lut = "off";
defparam \ac_write_block:sig_count[3]~0 .lut_mask = 64'h1111111111111111;
defparam \ac_write_block:sig_count[3]~0 .shared_arith = "off";

arriaii_lcell_comb \Add1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\ac_write_block:sig_count[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~21_sumout ),
	.cout(\Add1~22 ),
	.shareout());
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~21 .shared_arith = "off";

dffeas \ac_write_block:sig_count[5] (
	.clk(clk),
	.d(\Add1~21_sumout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\ac_write_block:sig_count[3]~3_combout ),
	.sload(gnd),
	.ena(\ac_write_block:sig_count[3]~1_combout ),
	.q(\ac_write_block:sig_count[5]~q ),
	.prn(vcc));
defparam \ac_write_block:sig_count[5] .is_wysiwyg = "true";
defparam \ac_write_block:sig_count[5] .power_up = "low";

arriaii_lcell_comb \Add1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\ac_write_block:sig_count[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~25_sumout ),
	.cout(\Add1~26 ),
	.shareout());
defparam \Add1~25 .extended_lut = "off";
defparam \Add1~25 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~25 .shared_arith = "off";

dffeas \ac_write_block:sig_count[6] (
	.clk(clk),
	.d(\Add1~25_sumout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\ac_write_block:sig_count[3]~3_combout ),
	.sload(gnd),
	.ena(\ac_write_block:sig_count[3]~1_combout ),
	.q(\ac_write_block:sig_count[6]~q ),
	.prn(vcc));
defparam \ac_write_block:sig_count[6] .is_wysiwyg = "true";
defparam \ac_write_block:sig_count[6] .power_up = "low";

arriaii_lcell_comb \Add1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\ac_write_block:sig_count[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~29_sumout ),
	.cout(),
	.shareout());
defparam \Add1~29 .extended_lut = "off";
defparam \Add1~29 .lut_mask = 64'h0000FFFF000000FF;
defparam \Add1~29 .shared_arith = "off";

dffeas \ac_write_block:sig_count[7] (
	.clk(clk),
	.d(\Add1~29_sumout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(!\ac_write_block:sig_count[3]~3_combout ),
	.sload(gnd),
	.ena(\ac_write_block:sig_count[3]~1_combout ),
	.q(\ac_write_block:sig_count[7]~q ),
	.prn(vcc));
defparam \ac_write_block:sig_count[7] .is_wysiwyg = "true";
defparam \ac_write_block:sig_count[7] .power_up = "low";

arriaii_lcell_comb \Selector91~0 (
	.dataa(!\ac_write_block:sig_count[2]~q ),
	.datab(!\ac_write_block:sig_count[3]~q ),
	.datac(!\ac_write_block:sig_count[6]~q ),
	.datad(!\ac_write_block:sig_count[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector91~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector91~0 .extended_lut = "off";
defparam \Selector91~0 .lut_mask = 64'h0001000100010001;
defparam \Selector91~0 .shared_arith = "off";

arriaii_lcell_comb \Selector32~0 (
	.dataa(!\sig_dgwb_state.s_write_ones~q ),
	.datab(!\sig_dgwb_state.s_write_0011_step~q ),
	.datac(!\sig_dgwb_state.s_write_01_pairs~q ),
	.datad(!\sig_dgwb_state.s_write_1100_step~q ),
	.datae(!\sig_dgwb_state.s_write_zeros~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector32~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector32~0 .extended_lut = "off";
defparam \Selector32~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \Selector32~0 .shared_arith = "off";

arriaii_lcell_comb \Selector91~1 (
	.dataa(!\ac_write_block:sig_count[5]~q ),
	.datab(!\ac_write_block:sig_count[4]~q ),
	.datac(!\ac_write_block:sig_count[3]~0_combout ),
	.datad(!\ac_write_block:sig_count[7]~q ),
	.datae(!\ac_write_block:sig_count[0]~q ),
	.dataf(!\Selector91~0_combout ),
	.datag(!\Selector32~0_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector91~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector91~1 .extended_lut = "on";
defparam \Selector91~1 .lut_mask = 64'h0000000008000800;
defparam \Selector91~1 .shared_arith = "off";

dffeas access_complete(
	.clk(clk),
	.d(\Selector91~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\access_complete~q ),
	.prn(vcc));
defparam access_complete.is_wysiwyg = "true";
defparam access_complete.power_up = "low";

arriaii_lcell_comb \Selector11~10 (
	.dataa(!\Selector11~4_combout ),
	.datab(!\access_complete~q ),
	.datac(!\sig_dgwb_last_state.s_write_0011_step~q ),
	.datad(!\sig_dgwb_state.s_write_0011_step~q ),
	.datae(!\Selector11~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector11~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector11~10 .extended_lut = "off";
defparam \Selector11~10 .lut_mask = 64'h0054555500545555;
defparam \Selector11~10 .shared_arith = "off";

dffeas \sig_dgwb_state.s_write_0011_step (
	.clk(clk),
	.d(\Selector11~10_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_state.s_write_0011_step~q ),
	.prn(vcc));
defparam \sig_dgwb_state.s_write_0011_step .is_wysiwyg = "true";
defparam \sig_dgwb_state.s_write_0011_step .power_up = "low";

arriaii_lcell_comb \Equal1~0 (
	.dataa(!\ac_write_block:sig_count[6]~q ),
	.datab(!\ac_write_block:sig_count[0]~q ),
	.datac(!\ac_write_block:sig_count[1]~q ),
	.datad(!\ac_write_block:sig_count[7]~q ),
	.datae(!\ac_write_block:sig_count[4]~q ),
	.dataf(!\ac_write_block:sig_count[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'h8000000000000000;
defparam \Equal1~0 .shared_arith = "off";

arriaii_lcell_comb \Selector26~0 (
	.dataa(!\sig_dgwb_state.s_write_ones~q ),
	.datab(!\sig_dgwb_state.s_write_zeros~q ),
	.datac(!\ac_write_block:sig_count[2]~q ),
	.datad(!\ac_write_block:sig_count[3]~q ),
	.datae(!\Equal1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector26~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector26~0 .extended_lut = "off";
defparam \Selector26~0 .lut_mask = 64'h4444074444440744;
defparam \Selector26~0 .shared_arith = "off";

arriaii_lcell_comb \Selector26~1 (
	.dataa(!\sig_dgwb_state.s_write_0011_step~q ),
	.datab(!\sig_dgwb_state.s_write_01_pairs~q ),
	.datac(!\Selector26~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector26~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector26~1 .extended_lut = "off";
defparam \Selector26~1 .lut_mask = 64'h5D5D5D5D5D5D5D5D;
defparam \Selector26~1 .shared_arith = "off";

arriaii_lcell_comb \sig_addr_cmd[0].addr[4]~0 (
	.dataa(!\sig_dgwb_state.s_write_ones~q ),
	.datab(!\sig_dgwb_last_state.s_write_ones~q ),
	.datac(!\sig_dgwb_state.s_write_1100_step~q ),
	.datad(!\sig_dgwb_last_state.s_write_1100_step~q ),
	.datae(!\sig_dgwb_last_state.s_write_zeros~q ),
	.dataf(!\sig_dgwb_state.s_write_zeros~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_addr_cmd[0].addr[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_addr_cmd[0].addr[4]~0 .extended_lut = "off";
defparam \sig_addr_cmd[0].addr[4]~0 .lut_mask = 64'hBBB0BBB00000BBB0;
defparam \sig_addr_cmd[0].addr[4]~0 .shared_arith = "off";

arriaii_lcell_comb \sig_addr_cmd[0].addr[4]~1 (
	.dataa(!\sig_dgwb_state.s_write_wlat~q ),
	.datab(!\sig_dgwb_last_state.s_write_0011_step~q ),
	.datac(!\sig_dgwb_state.s_write_0011_step~q ),
	.datad(!\sig_dgwb_last_state.s_write_wlat~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_addr_cmd[0].addr[4]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_addr_cmd[0].addr[4]~1 .extended_lut = "off";
defparam \sig_addr_cmd[0].addr[4]~1 .lut_mask = 64'h0357035703570357;
defparam \sig_addr_cmd[0].addr[4]~1 .shared_arith = "off";

arriaii_lcell_comb \sig_addr_cmd[0].addr[4]~4 (
	.dataa(!\sig_dgwb_last_state.s_write_01_pairs~q ),
	.datab(!\sig_dgwb_state.s_write_01_pairs~q ),
	.datac(!\ac_write_block:sig_count[2]~q ),
	.datad(!\ac_write_block:sig_count[3]~q ),
	.datae(!\sig_dgwb_state.s_write_ones~q ),
	.dataf(!\sig_dgwb_state.s_release_admin~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_addr_cmd[0].addr[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_addr_cmd[0].addr[4]~4 .extended_lut = "off";
defparam \sig_addr_cmd[0].addr[4]~4 .lut_mask = 64'hDCCCDCC000000000;
defparam \sig_addr_cmd[0].addr[4]~4 .shared_arith = "off";

arriaii_lcell_comb \sig_addr_cmd[0].addr[4]~5 (
	.dataa(!\sig_dgwb_state.s_write_01_pairs~q ),
	.datab(!\Equal1~0_combout ),
	.datac(!\sig_dgwb_state.s_write_ones~q ),
	.datad(!\sig_dgwb_state.s_write_zeros~q ),
	.datae(!\sig_dgwb_state.s_wait_admin~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_addr_cmd[0].addr[4]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_addr_cmd[0].addr[4]~5 .extended_lut = "off";
defparam \sig_addr_cmd[0].addr[4]~5 .lut_mask = 64'hB3330000B3330000;
defparam \sig_addr_cmd[0].addr[4]~5 .shared_arith = "off";

arriaii_lcell_comb \sig_addr_cmd[0].addr[4]~2 (
	.dataa(!\sig_addr_cmd[0].addr[4]~0_combout ),
	.datab(!\sig_addr_cmd[0].addr[4]~1_combout ),
	.datac(!\sig_dgwb_state.s_write_btp~q ),
	.datad(!\sig_dgwb_state.s_write_mtp~q ),
	.datae(!\sig_addr_cmd[0].addr[4]~4_combout ),
	.dataf(!\sig_addr_cmd[0].addr[4]~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_addr_cmd[0].addr[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_addr_cmd[0].addr[4]~2 .extended_lut = "off";
defparam \sig_addr_cmd[0].addr[4]~2 .lut_mask = 64'h0000000000004000;
defparam \sig_addr_cmd[0].addr[4]~2 .shared_arith = "off";

arriaii_lcell_comb \sig_addr_cmd~0 (
	.dataa(!\ac_write_block:sig_count[2]~q ),
	.datab(!\ac_write_block:sig_count[3]~q ),
	.datac(!\Equal1~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_addr_cmd~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_addr_cmd~0 .extended_lut = "off";
defparam \sig_addr_cmd~0 .lut_mask = 64'h0E0E0E0E0E0E0E0E;
defparam \sig_addr_cmd~0 .shared_arith = "off";

arriaii_lcell_comb \Selector25~0 (
	.dataa(!\sig_dgwb_state.s_write_ones~q ),
	.datab(!\sig_dgwb_state.s_write_01_pairs~q ),
	.datac(!\sig_dgwb_state.s_write_zeros~q ),
	.datad(!\sig_addr_cmd~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector25~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector25~0 .extended_lut = "off";
defparam \Selector25~0 .lut_mask = 64'h7F737F737F737F73;
defparam \Selector25~0 .shared_arith = "off";

arriaii_lcell_comb \Selector24~0 (
	.dataa(!\sig_dgwb_state.s_write_0011_step~q ),
	.datab(!\sig_dgwb_state.s_write_1100_step~q ),
	.datac(!\sig_dgwb_state.s_write_zeros~q ),
	.datad(gnd),
	.datae(!\ac_write_block:sig_count[3]~q ),
	.dataf(!\Equal1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector24~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector24~0 .extended_lut = "off";
defparam \Selector24~0 .lut_mask = 64'h7F7F7F7F77777F7F;
defparam \Selector24~0 .shared_arith = "off";

arriaii_lcell_comb \Selector23~0 (
	.dataa(!\sig_dgwb_state.s_write_ones~q ),
	.datab(!\sig_dgwb_state.s_write_01_pairs~q ),
	.datac(gnd),
	.datad(!\ac_write_block:sig_count[3]~q ),
	.datae(!\Equal1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector23~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector23~0 .extended_lut = "off";
defparam \Selector23~0 .lut_mask = 64'h7777337777773377;
defparam \Selector23~0 .shared_arith = "off";

dffeas \sig_dgwb_last_state.s_release_admin (
	.clk(clk),
	.d(\sig_dgwb_state.s_release_admin~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_last_state.s_release_admin~q ),
	.prn(vcc));
defparam \sig_dgwb_last_state.s_release_admin .is_wysiwyg = "true";
defparam \sig_dgwb_last_state.s_release_admin .power_up = "low";

arriaii_lcell_comb \ac_handshake_proc~2 (
	.dataa(!\sig_dgwb_last_state.s_release_admin~q ),
	.datab(!\sig_dgwb_state.s_idle~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_handshake_proc~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_handshake_proc~2 .extended_lut = "off";
defparam \ac_handshake_proc~2 .lut_mask = 64'h4444444444444444;
defparam \ac_handshake_proc~2 .shared_arith = "off";

arriaii_lcell_comb \dgwb_dqs_burst~0 (
	.dataa(!\sig_dgwb_state.s_idle~q ),
	.datab(!\sig_dgwb_state.s_write_btp~q ),
	.datac(!\sig_dgwb_state.s_write_mtp~q ),
	.datad(!\sig_dgwb_state.s_wait_admin~q ),
	.datae(!\sig_dgwb_state.s_release_admin~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dgwb_dqs_burst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dgwb_dqs_burst~0 .extended_lut = "off";
defparam \dgwb_dqs_burst~0 .lut_mask = 64'h4000000040000000;
defparam \dgwb_dqs_burst~0 .shared_arith = "off";

arriaii_lcell_comb \ac_handshake_proc~3 (
	.dataa(!\sig_dgwb_state.s_idle~q ),
	.datab(!\sig_dgwb_state.s_release_admin~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_handshake_proc~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_handshake_proc~3 .extended_lut = "off";
defparam \ac_handshake_proc~3 .lut_mask = 64'h4444444444444444;
defparam \ac_handshake_proc~3 .shared_arith = "off";

arriaii_lcell_comb \Selector50~0 (
	.dataa(!\sig_dgwb_last_state.s_write_0011_step~q ),
	.datab(!\sig_dgwb_state.s_write_0011_step~q ),
	.datac(!\sig_dgwb_state.s_write_1100_step~q ),
	.datad(!\sig_dgwb_last_state.s_write_1100_step~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector50~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector50~0 .extended_lut = "off";
defparam \Selector50~0 .lut_mask = 64'h2F222F222F222F22;
defparam \Selector50~0 .shared_arith = "off";

arriaii_lcell_comb \Selector50~1 (
	.dataa(!\sig_dgwb_state.s_write_ones~q ),
	.datab(!\sig_dgwb_state.s_write_wlat~q ),
	.datac(!\sig_dgwb_last_state.s_write_wlat~q ),
	.datad(!\sig_dgwb_last_state.s_write_ones~q ),
	.datae(!\sig_addr_cmd~0_combout ),
	.dataf(!\Selector50~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector50~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector50~1 .extended_lut = "off";
defparam \Selector50~1 .lut_mask = 64'hCFCFCF8A00000000;
defparam \Selector50~1 .shared_arith = "off";

arriaii_lcell_comb \Selector50~2 (
	.dataa(!\Selector11~5_combout ),
	.datab(!\Selector6~1_combout ),
	.datac(!\ac_write_block:sig_count[2]~q ),
	.datad(!\ac_write_block:sig_count[3]~q ),
	.datae(!\Equal1~0_combout ),
	.dataf(!\Selector50~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector50~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector50~2 .extended_lut = "off";
defparam \Selector50~2 .lut_mask = 64'hFFFFFFFF00007333;
defparam \Selector50~2 .shared_arith = "off";

arriaii_lcell_comb \sig_addr_cmd[0].addr[12]~0 (
	.dataa(!sig_addr_cmd0addr12),
	.datab(!\sig_dgwb_state.s_write_wlat~q ),
	.datac(!\sig_addr_cmd[0].addr[4]~2_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sig_addr_cmd[0].addr[12]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sig_addr_cmd[0].addr[12]~0 .extended_lut = "off";
defparam \sig_addr_cmd[0].addr[12]~0 .lut_mask = 64'h5353535353535353;
defparam \sig_addr_cmd[0].addr[12]~0 .shared_arith = "off";

arriaii_lcell_comb \Selector58~0 (
	.dataa(!\sig_dgwb_state.s_write_ones~q ),
	.datab(!\sig_dgwb_state.s_write_0011_step~q ),
	.datac(!\ac_write_block:sig_count[0]~q ),
	.datad(!\ac_write_block:sig_count[3]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector58~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector58~0 .extended_lut = "off";
defparam \Selector58~0 .lut_mask = 64'h777F777F777F777F;
defparam \Selector58~0 .shared_arith = "off";

arriaii_lcell_comb \Selector74~0 (
	.dataa(!\sig_dgwb_state.s_write_ones~q ),
	.datab(!\sig_dgwb_state.s_write_1100_step~q ),
	.datac(!\ac_write_block:sig_count[0]~q ),
	.datad(!\ac_write_block:sig_count[3]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector74~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector74~0 .extended_lut = "off";
defparam \Selector74~0 .lut_mask = 64'h777F777F777F777F;
defparam \Selector74~0 .shared_arith = "off";

arriaii_lcell_comb \WideOr4~0 (
	.dataa(!\sig_dgwb_state.s_write_ones~q ),
	.datab(!\sig_dgwb_state.s_write_0011_step~q ),
	.datac(!\sig_dgwb_state.s_write_01_pairs~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr4~0 .extended_lut = "off";
defparam \WideOr4~0 .lut_mask = 64'h8080808080808080;
defparam \WideOr4~0 .shared_arith = "off";

arriaii_lcell_comb \Selector66~0 (
	.dataa(!\ac_write_block:sig_count[0]~q ),
	.datab(!\ac_write_block:sig_count[3]~0_combout ),
	.datac(!\WideOr4~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector66~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector66~0 .extended_lut = "off";
defparam \Selector66~0 .lut_mask = 64'hF1F1F1F1F1F1F1F1;
defparam \Selector66~0 .shared_arith = "off";

arriaii_lcell_comb \WideOr7~0 (
	.dataa(!\sig_dgwb_state.s_write_ones~q ),
	.datab(!\sig_dgwb_state.s_write_01_pairs~q ),
	.datac(!\sig_dgwb_state.s_write_1100_step~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr7~0 .extended_lut = "off";
defparam \WideOr7~0 .lut_mask = 64'h8080808080808080;
defparam \WideOr7~0 .shared_arith = "off";

arriaii_lcell_comb \Selector82~0 (
	.dataa(!\ac_write_block:sig_count[0]~q ),
	.datab(!\WideOr7~0_combout ),
	.datac(!\ac_write_block:sig_count[3]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector82~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector82~0 .extended_lut = "off";
defparam \Selector82~0 .lut_mask = 64'hCDCDCDCDCDCDCDCD;
defparam \Selector82~0 .shared_arith = "off";

arriaii_lcell_comb \Selector57~0 (
	.dataa(!\sig_dgwb_state.s_write_ones~q ),
	.datab(!\sig_dgwb_state.s_write_0011_step~q ),
	.datac(!\ac_write_block:sig_count[1]~q ),
	.datad(!\ac_write_block:sig_count[3]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector57~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector57~0 .extended_lut = "off";
defparam \Selector57~0 .lut_mask = 64'h777F777F777F777F;
defparam \Selector57~0 .shared_arith = "off";

arriaii_lcell_comb \Selector73~0 (
	.dataa(!\sig_dgwb_state.s_write_ones~q ),
	.datab(!\sig_dgwb_state.s_write_1100_step~q ),
	.datac(!\ac_write_block:sig_count[1]~q ),
	.datad(!\ac_write_block:sig_count[3]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector73~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector73~0 .extended_lut = "off";
defparam \Selector73~0 .lut_mask = 64'h777F777F777F777F;
defparam \Selector73~0 .shared_arith = "off";

arriaii_lcell_comb \Selector65~0 (
	.dataa(!\ac_write_block:sig_count[1]~q ),
	.datab(!\ac_write_block:sig_count[3]~0_combout ),
	.datac(!\WideOr4~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector65~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector65~0 .extended_lut = "off";
defparam \Selector65~0 .lut_mask = 64'hF1F1F1F1F1F1F1F1;
defparam \Selector65~0 .shared_arith = "off";

arriaii_lcell_comb \Selector81~0 (
	.dataa(!\ac_write_block:sig_count[1]~q ),
	.datab(!\WideOr7~0_combout ),
	.datac(!\ac_write_block:sig_count[3]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector81~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector81~0 .extended_lut = "off";
defparam \Selector81~0 .lut_mask = 64'hCDCDCDCDCDCDCDCD;
defparam \Selector81~0 .shared_arith = "off";

arriaii_lcell_comb \Selector56~0 (
	.dataa(!\sig_dgwb_state.s_write_ones~q ),
	.datab(!\sig_dgwb_state.s_write_0011_step~q ),
	.datac(!\ac_write_block:sig_count[2]~q ),
	.datad(!\ac_write_block:sig_count[3]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector56~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector56~0 .extended_lut = "off";
defparam \Selector56~0 .lut_mask = 64'h777F777F777F777F;
defparam \Selector56~0 .shared_arith = "off";

arriaii_lcell_comb \Selector72~0 (
	.dataa(!\sig_dgwb_state.s_write_ones~q ),
	.datab(!\sig_dgwb_state.s_write_1100_step~q ),
	.datac(!\ac_write_block:sig_count[2]~q ),
	.datad(!\ac_write_block:sig_count[3]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector72~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector72~0 .extended_lut = "off";
defparam \Selector72~0 .lut_mask = 64'h777F777F777F777F;
defparam \Selector72~0 .shared_arith = "off";

arriaii_lcell_comb \Selector64~0 (
	.dataa(!\ac_write_block:sig_count[2]~q ),
	.datab(!\ac_write_block:sig_count[3]~0_combout ),
	.datac(!\WideOr4~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector64~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector64~0 .extended_lut = "off";
defparam \Selector64~0 .lut_mask = 64'hF1F1F1F1F1F1F1F1;
defparam \Selector64~0 .shared_arith = "off";

arriaii_lcell_comb \Selector80~0 (
	.dataa(!\ac_write_block:sig_count[2]~q ),
	.datab(!\WideOr7~0_combout ),
	.datac(!\ac_write_block:sig_count[3]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector80~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector80~0 .extended_lut = "off";
defparam \Selector80~0 .lut_mask = 64'hCDCDCDCDCDCDCDCD;
defparam \Selector80~0 .shared_arith = "off";

arriaii_lcell_comb \Selector55~0 (
	.dataa(!\sig_dgwb_state.s_write_ones~q ),
	.datab(!\sig_dgwb_state.s_write_0011_step~q ),
	.datac(!\ac_write_block:sig_count[3]~q ),
	.datad(!\ac_write_block:sig_count[3]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector55~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector55~0 .extended_lut = "off";
defparam \Selector55~0 .lut_mask = 64'h777F777F777F777F;
defparam \Selector55~0 .shared_arith = "off";

arriaii_lcell_comb \Selector71~0 (
	.dataa(!\sig_dgwb_state.s_write_ones~q ),
	.datab(!\sig_dgwb_state.s_write_1100_step~q ),
	.datac(!\ac_write_block:sig_count[3]~q ),
	.datad(!\ac_write_block:sig_count[3]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector71~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector71~0 .extended_lut = "off";
defparam \Selector71~0 .lut_mask = 64'h777F777F777F777F;
defparam \Selector71~0 .shared_arith = "off";

arriaii_lcell_comb \Selector63~0 (
	.dataa(!\ac_write_block:sig_count[3]~q ),
	.datab(!\ac_write_block:sig_count[3]~0_combout ),
	.datac(!\WideOr4~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector63~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector63~0 .extended_lut = "off";
defparam \Selector63~0 .lut_mask = 64'hF1F1F1F1F1F1F1F1;
defparam \Selector63~0 .shared_arith = "off";

arriaii_lcell_comb \Selector79~0 (
	.dataa(!\ac_write_block:sig_count[3]~q ),
	.datab(!\WideOr7~0_combout ),
	.datac(!\ac_write_block:sig_count[3]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector79~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector79~0 .extended_lut = "off";
defparam \Selector79~0 .lut_mask = 64'hCDCDCDCDCDCDCDCD;
defparam \Selector79~0 .shared_arith = "off";

arriaii_lcell_comb \Selector54~0 (
	.dataa(!\sig_dgwb_state.s_write_ones~q ),
	.datab(!\sig_dgwb_state.s_write_0011_step~q ),
	.datac(!\ac_write_block:sig_count[4]~q ),
	.datad(!\ac_write_block:sig_count[3]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector54~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector54~0 .extended_lut = "off";
defparam \Selector54~0 .lut_mask = 64'h777F777F777F777F;
defparam \Selector54~0 .shared_arith = "off";

arriaii_lcell_comb \Selector70~0 (
	.dataa(!\sig_dgwb_state.s_write_ones~q ),
	.datab(!\sig_dgwb_state.s_write_1100_step~q ),
	.datac(!\ac_write_block:sig_count[4]~q ),
	.datad(!\ac_write_block:sig_count[3]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector70~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector70~0 .extended_lut = "off";
defparam \Selector70~0 .lut_mask = 64'h777F777F777F777F;
defparam \Selector70~0 .shared_arith = "off";

arriaii_lcell_comb \Selector62~0 (
	.dataa(!\ac_write_block:sig_count[4]~q ),
	.datab(!\ac_write_block:sig_count[3]~0_combout ),
	.datac(!\WideOr4~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector62~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector62~0 .extended_lut = "off";
defparam \Selector62~0 .lut_mask = 64'hF1F1F1F1F1F1F1F1;
defparam \Selector62~0 .shared_arith = "off";

arriaii_lcell_comb \Selector78~0 (
	.dataa(!\ac_write_block:sig_count[4]~q ),
	.datab(!\WideOr7~0_combout ),
	.datac(!\ac_write_block:sig_count[3]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector78~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector78~0 .extended_lut = "off";
defparam \Selector78~0 .lut_mask = 64'hCDCDCDCDCDCDCDCD;
defparam \Selector78~0 .shared_arith = "off";

arriaii_lcell_comb \Selector53~0 (
	.dataa(!\sig_dgwb_state.s_write_ones~q ),
	.datab(!\sig_dgwb_state.s_write_0011_step~q ),
	.datac(!\ac_write_block:sig_count[5]~q ),
	.datad(!\ac_write_block:sig_count[3]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector53~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector53~0 .extended_lut = "off";
defparam \Selector53~0 .lut_mask = 64'h777F777F777F777F;
defparam \Selector53~0 .shared_arith = "off";

arriaii_lcell_comb \Selector69~0 (
	.dataa(!\sig_dgwb_state.s_write_ones~q ),
	.datab(!\sig_dgwb_state.s_write_1100_step~q ),
	.datac(!\ac_write_block:sig_count[5]~q ),
	.datad(!\ac_write_block:sig_count[3]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector69~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector69~0 .extended_lut = "off";
defparam \Selector69~0 .lut_mask = 64'h777F777F777F777F;
defparam \Selector69~0 .shared_arith = "off";

arriaii_lcell_comb \Selector61~0 (
	.dataa(!\ac_write_block:sig_count[5]~q ),
	.datab(!\ac_write_block:sig_count[3]~0_combout ),
	.datac(!\WideOr4~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector61~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector61~0 .extended_lut = "off";
defparam \Selector61~0 .lut_mask = 64'hF1F1F1F1F1F1F1F1;
defparam \Selector61~0 .shared_arith = "off";

arriaii_lcell_comb \Selector77~0 (
	.dataa(!\ac_write_block:sig_count[5]~q ),
	.datab(!\WideOr7~0_combout ),
	.datac(!\ac_write_block:sig_count[3]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector77~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector77~0 .extended_lut = "off";
defparam \Selector77~0 .lut_mask = 64'hCDCDCDCDCDCDCDCD;
defparam \Selector77~0 .shared_arith = "off";

arriaii_lcell_comb \Selector52~0 (
	.dataa(!\sig_dgwb_state.s_write_ones~q ),
	.datab(!\sig_dgwb_state.s_write_0011_step~q ),
	.datac(!\ac_write_block:sig_count[6]~q ),
	.datad(!\ac_write_block:sig_count[3]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector52~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector52~0 .extended_lut = "off";
defparam \Selector52~0 .lut_mask = 64'h777F777F777F777F;
defparam \Selector52~0 .shared_arith = "off";

arriaii_lcell_comb \Selector68~0 (
	.dataa(!\sig_dgwb_state.s_write_ones~q ),
	.datab(!\sig_dgwb_state.s_write_1100_step~q ),
	.datac(!\ac_write_block:sig_count[6]~q ),
	.datad(!\ac_write_block:sig_count[3]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector68~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector68~0 .extended_lut = "off";
defparam \Selector68~0 .lut_mask = 64'h777F777F777F777F;
defparam \Selector68~0 .shared_arith = "off";

arriaii_lcell_comb \Selector60~0 (
	.dataa(!\ac_write_block:sig_count[6]~q ),
	.datab(!\ac_write_block:sig_count[3]~0_combout ),
	.datac(!\WideOr4~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector60~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector60~0 .extended_lut = "off";
defparam \Selector60~0 .lut_mask = 64'hF1F1F1F1F1F1F1F1;
defparam \Selector60~0 .shared_arith = "off";

arriaii_lcell_comb \Selector76~0 (
	.dataa(!\ac_write_block:sig_count[6]~q ),
	.datab(!\WideOr7~0_combout ),
	.datac(!\ac_write_block:sig_count[3]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector76~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector76~0 .extended_lut = "off";
defparam \Selector76~0 .lut_mask = 64'hCDCDCDCDCDCDCDCD;
defparam \Selector76~0 .shared_arith = "off";

arriaii_lcell_comb \Selector51~0 (
	.dataa(!\sig_dgwb_state.s_write_ones~q ),
	.datab(!\sig_dgwb_state.s_write_0011_step~q ),
	.datac(!\ac_write_block:sig_count[7]~q ),
	.datad(!\ac_write_block:sig_count[3]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector51~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector51~0 .extended_lut = "off";
defparam \Selector51~0 .lut_mask = 64'h777F777F777F777F;
defparam \Selector51~0 .shared_arith = "off";

arriaii_lcell_comb \Selector67~0 (
	.dataa(!\sig_dgwb_state.s_write_ones~q ),
	.datab(!\sig_dgwb_state.s_write_1100_step~q ),
	.datac(!\ac_write_block:sig_count[7]~q ),
	.datad(!\ac_write_block:sig_count[3]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector67~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector67~0 .extended_lut = "off";
defparam \Selector67~0 .lut_mask = 64'h777F777F777F777F;
defparam \Selector67~0 .shared_arith = "off";

arriaii_lcell_comb \Selector59~0 (
	.dataa(!\ac_write_block:sig_count[7]~q ),
	.datab(!\ac_write_block:sig_count[3]~0_combout ),
	.datac(!\WideOr4~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector59~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector59~0 .extended_lut = "off";
defparam \Selector59~0 .lut_mask = 64'hF1F1F1F1F1F1F1F1;
defparam \Selector59~0 .shared_arith = "off";

arriaii_lcell_comb \Selector75~0 (
	.dataa(!\ac_write_block:sig_count[7]~q ),
	.datab(!\WideOr7~0_combout ),
	.datac(!\ac_write_block:sig_count[3]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector75~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector75~0 .extended_lut = "off";
defparam \Selector75~0 .lut_mask = 64'hCDCDCDCDCDCDCDCD;
defparam \Selector75~0 .shared_arith = "off";

dffeas \sig_dgwb_last_state.s_idle (
	.clk(clk),
	.d(\sig_dgwb_state.s_idle~q ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sig_dgwb_last_state.s_idle~q ),
	.prn(vcc));
defparam \sig_dgwb_last_state.s_idle .is_wysiwyg = "true";
defparam \sig_dgwb_last_state.s_idle .power_up = "low";

arriaii_lcell_comb \ac_handshake_proc~4 (
	.dataa(!\sig_dgwb_state.s_wait_admin~q ),
	.datab(!\sig_dgwb_last_state.s_idle~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac_handshake_proc~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac_handshake_proc~4 .extended_lut = "off";
defparam \ac_handshake_proc~4 .lut_mask = 64'h4444444444444444;
defparam \ac_handshake_proc~4 .shared_arith = "off";

endmodule

module ddr3_int_ddr3_int_phy_alt_mem_phy_write_dp (
	phy_clk_1x,
	mem_clk_2x,
	write_clk_2x,
	wdp_dm_l_2x_0,
	wdp_dm_h_2x_0,
	wdp_dm_l_2x_1,
	wdp_dm_h_2x_1,
	wdp_dm_l_2x_2,
	wdp_dm_h_2x_2,
	wdp_dm_l_2x_3,
	wdp_dm_h_2x_3,
	wdp_wdata_l_2x_0,
	wdp_wdata_h_2x_0,
	dq_oe_2x_0,
	wdp_wdata_l_2x_1,
	wdp_wdata_h_2x_1,
	wdp_wdata_l_2x_2,
	wdp_wdata_h_2x_2,
	wdp_wdata_l_2x_3,
	wdp_wdata_h_2x_3,
	wdp_wdata_l_2x_4,
	wdp_wdata_h_2x_4,
	dq_oe_2x_1,
	wdp_wdata_l_2x_5,
	wdp_wdata_h_2x_5,
	wdp_wdata_l_2x_6,
	wdp_wdata_h_2x_6,
	wdp_wdata_l_2x_7,
	wdp_wdata_h_2x_7,
	wdp_wdata_l_2x_8,
	wdp_wdata_h_2x_8,
	dq_oe_2x_2,
	wdp_wdata_l_2x_9,
	wdp_wdata_h_2x_9,
	wdp_wdata_l_2x_10,
	wdp_wdata_h_2x_10,
	wdp_wdata_l_2x_11,
	wdp_wdata_h_2x_11,
	wdp_wdata_l_2x_12,
	wdp_wdata_h_2x_12,
	dq_oe_2x_3,
	wdp_wdata_l_2x_13,
	wdp_wdata_h_2x_13,
	wdp_wdata_l_2x_14,
	wdp_wdata_h_2x_14,
	wdp_wdata_l_2x_15,
	wdp_wdata_h_2x_15,
	wdp_wdata_l_2x_16,
	wdp_wdata_h_2x_16,
	dq_oe_2x_4,
	wdp_wdata_l_2x_17,
	wdp_wdata_h_2x_17,
	wdp_wdata_l_2x_18,
	wdp_wdata_h_2x_18,
	wdp_wdata_l_2x_19,
	wdp_wdata_h_2x_19,
	wdp_wdata_l_2x_20,
	wdp_wdata_h_2x_20,
	dq_oe_2x_5,
	wdp_wdata_l_2x_21,
	wdp_wdata_h_2x_21,
	wdp_wdata_l_2x_22,
	wdp_wdata_h_2x_22,
	wdp_wdata_l_2x_23,
	wdp_wdata_h_2x_23,
	wdp_wdata_l_2x_24,
	wdp_wdata_h_2x_24,
	dq_oe_2x_6,
	wdp_wdata_l_2x_25,
	wdp_wdata_h_2x_25,
	wdp_wdata_l_2x_26,
	wdp_wdata_h_2x_26,
	wdp_wdata_l_2x_27,
	wdp_wdata_h_2x_27,
	wdp_wdata_l_2x_28,
	wdp_wdata_h_2x_28,
	dq_oe_2x_7,
	wdp_wdata_l_2x_29,
	wdp_wdata_h_2x_29,
	wdp_wdata_l_2x_30,
	wdp_wdata_h_2x_30,
	wdp_wdata_l_2x_31,
	wdp_wdata_h_2x_31,
	q_b_96,
	q_b_32,
	q_b_64,
	q_b_0,
	q_b_97,
	q_b_33,
	q_b_65,
	q_b_1,
	q_b_98,
	q_b_34,
	q_b_66,
	q_b_2,
	q_b_99,
	q_b_35,
	q_b_67,
	q_b_3,
	q_b_100,
	q_b_36,
	q_b_68,
	q_b_4,
	q_b_101,
	q_b_37,
	q_b_69,
	q_b_5,
	q_b_102,
	q_b_38,
	q_b_70,
	q_b_6,
	q_b_103,
	q_b_39,
	q_b_71,
	q_b_7,
	q_b_104,
	q_b_40,
	q_b_72,
	q_b_8,
	q_b_105,
	q_b_41,
	q_b_73,
	q_b_9,
	q_b_106,
	q_b_42,
	q_b_74,
	q_b_10,
	q_b_107,
	q_b_43,
	q_b_75,
	q_b_11,
	q_b_108,
	q_b_44,
	q_b_76,
	q_b_12,
	q_b_109,
	q_b_45,
	q_b_77,
	q_b_13,
	q_b_110,
	q_b_46,
	q_b_78,
	q_b_14,
	q_b_111,
	q_b_47,
	q_b_79,
	q_b_15,
	q_b_112,
	q_b_48,
	q_b_80,
	q_b_16,
	q_b_113,
	q_b_49,
	q_b_81,
	q_b_17,
	q_b_114,
	q_b_50,
	q_b_82,
	q_b_18,
	q_b_115,
	q_b_51,
	q_b_83,
	q_b_19,
	q_b_116,
	q_b_52,
	q_b_84,
	q_b_20,
	q_b_117,
	q_b_53,
	q_b_85,
	q_b_21,
	q_b_118,
	q_b_54,
	q_b_86,
	q_b_22,
	q_b_119,
	q_b_55,
	q_b_87,
	q_b_23,
	q_b_120,
	q_b_56,
	q_b_88,
	q_b_24,
	q_b_121,
	q_b_57,
	q_b_89,
	q_b_25,
	q_b_122,
	q_b_58,
	q_b_90,
	q_b_26,
	q_b_123,
	q_b_59,
	q_b_91,
	q_b_27,
	q_b_124,
	q_b_60,
	q_b_92,
	q_b_28,
	q_b_125,
	q_b_61,
	q_b_93,
	q_b_29,
	q_b_126,
	q_b_62,
	q_b_94,
	q_b_30,
	q_b_127,
	q_b_63,
	q_b_95,
	q_b_31,
	reset_phy_clk_1x_n,
	ctl_init_fail,
	ctl_init_success,
	reset_write_clk_2x_n,
	dqs_burst_2x_r3_0,
	dqs_burst_2x_r3_1,
	dqs_burst_2x_r3_2,
	dqs_burst_2x_r3_3,
	reset_mem_clk_2x_n,
	afi_dm_4,
	dgwb_wdp_ovride,
	seq_wdp_ovride,
	afi_dm_12,
	afi_dm_0,
	afi_dm_8,
	afi_dm_5,
	afi_dm_13,
	afi_dm_1,
	afi_dm_9,
	afi_dm_6,
	afi_dm_14,
	afi_dm_2,
	afi_dm_10,
	afi_dm_7,
	afi_dm_15,
	afi_dm_3,
	afi_dm_11,
	int_wdata_valid,
	dgwb_wdata_120,
	dgwb_wdata_56,
	dgwb_wdata_88,
	dgwb_wdata_24,
	dgwb_wdata_121,
	dgwb_wdata_57,
	dgwb_wdata_89,
	dgwb_wdata_25,
	dgwb_wdata_122,
	dgwb_wdata_58,
	dgwb_wdata_90,
	dgwb_wdata_26,
	dgwb_wdata_123,
	dgwb_wdata_59,
	dgwb_wdata_91,
	dgwb_wdata_27,
	dgwb_wdata_124,
	dgwb_wdata_60,
	dgwb_wdata_92,
	dgwb_wdata_28,
	dgwb_wdata_125,
	dgwb_wdata_61,
	dgwb_wdata_93,
	dgwb_wdata_29,
	dgwb_wdata_126,
	dgwb_wdata_62,
	dgwb_wdata_94,
	dgwb_wdata_30,
	dgwb_wdata_127,
	dgwb_wdata_63,
	dgwb_wdata_95,
	dgwb_wdata_31,
	int_dqs_burst,
	int_dqs_burst_hr,
	dgwb_wdp_ovride1)/* synthesis synthesis_greybox=0 */;
input 	phy_clk_1x;
input 	mem_clk_2x;
input 	write_clk_2x;
output 	wdp_dm_l_2x_0;
output 	wdp_dm_h_2x_0;
output 	wdp_dm_l_2x_1;
output 	wdp_dm_h_2x_1;
output 	wdp_dm_l_2x_2;
output 	wdp_dm_h_2x_2;
output 	wdp_dm_l_2x_3;
output 	wdp_dm_h_2x_3;
output 	wdp_wdata_l_2x_0;
output 	wdp_wdata_h_2x_0;
output 	dq_oe_2x_0;
output 	wdp_wdata_l_2x_1;
output 	wdp_wdata_h_2x_1;
output 	wdp_wdata_l_2x_2;
output 	wdp_wdata_h_2x_2;
output 	wdp_wdata_l_2x_3;
output 	wdp_wdata_h_2x_3;
output 	wdp_wdata_l_2x_4;
output 	wdp_wdata_h_2x_4;
output 	dq_oe_2x_1;
output 	wdp_wdata_l_2x_5;
output 	wdp_wdata_h_2x_5;
output 	wdp_wdata_l_2x_6;
output 	wdp_wdata_h_2x_6;
output 	wdp_wdata_l_2x_7;
output 	wdp_wdata_h_2x_7;
output 	wdp_wdata_l_2x_8;
output 	wdp_wdata_h_2x_8;
output 	dq_oe_2x_2;
output 	wdp_wdata_l_2x_9;
output 	wdp_wdata_h_2x_9;
output 	wdp_wdata_l_2x_10;
output 	wdp_wdata_h_2x_10;
output 	wdp_wdata_l_2x_11;
output 	wdp_wdata_h_2x_11;
output 	wdp_wdata_l_2x_12;
output 	wdp_wdata_h_2x_12;
output 	dq_oe_2x_3;
output 	wdp_wdata_l_2x_13;
output 	wdp_wdata_h_2x_13;
output 	wdp_wdata_l_2x_14;
output 	wdp_wdata_h_2x_14;
output 	wdp_wdata_l_2x_15;
output 	wdp_wdata_h_2x_15;
output 	wdp_wdata_l_2x_16;
output 	wdp_wdata_h_2x_16;
output 	dq_oe_2x_4;
output 	wdp_wdata_l_2x_17;
output 	wdp_wdata_h_2x_17;
output 	wdp_wdata_l_2x_18;
output 	wdp_wdata_h_2x_18;
output 	wdp_wdata_l_2x_19;
output 	wdp_wdata_h_2x_19;
output 	wdp_wdata_l_2x_20;
output 	wdp_wdata_h_2x_20;
output 	dq_oe_2x_5;
output 	wdp_wdata_l_2x_21;
output 	wdp_wdata_h_2x_21;
output 	wdp_wdata_l_2x_22;
output 	wdp_wdata_h_2x_22;
output 	wdp_wdata_l_2x_23;
output 	wdp_wdata_h_2x_23;
output 	wdp_wdata_l_2x_24;
output 	wdp_wdata_h_2x_24;
output 	dq_oe_2x_6;
output 	wdp_wdata_l_2x_25;
output 	wdp_wdata_h_2x_25;
output 	wdp_wdata_l_2x_26;
output 	wdp_wdata_h_2x_26;
output 	wdp_wdata_l_2x_27;
output 	wdp_wdata_h_2x_27;
output 	wdp_wdata_l_2x_28;
output 	wdp_wdata_h_2x_28;
output 	dq_oe_2x_7;
output 	wdp_wdata_l_2x_29;
output 	wdp_wdata_h_2x_29;
output 	wdp_wdata_l_2x_30;
output 	wdp_wdata_h_2x_30;
output 	wdp_wdata_l_2x_31;
output 	wdp_wdata_h_2x_31;
input 	q_b_96;
input 	q_b_32;
input 	q_b_64;
input 	q_b_0;
input 	q_b_97;
input 	q_b_33;
input 	q_b_65;
input 	q_b_1;
input 	q_b_98;
input 	q_b_34;
input 	q_b_66;
input 	q_b_2;
input 	q_b_99;
input 	q_b_35;
input 	q_b_67;
input 	q_b_3;
input 	q_b_100;
input 	q_b_36;
input 	q_b_68;
input 	q_b_4;
input 	q_b_101;
input 	q_b_37;
input 	q_b_69;
input 	q_b_5;
input 	q_b_102;
input 	q_b_38;
input 	q_b_70;
input 	q_b_6;
input 	q_b_103;
input 	q_b_39;
input 	q_b_71;
input 	q_b_7;
input 	q_b_104;
input 	q_b_40;
input 	q_b_72;
input 	q_b_8;
input 	q_b_105;
input 	q_b_41;
input 	q_b_73;
input 	q_b_9;
input 	q_b_106;
input 	q_b_42;
input 	q_b_74;
input 	q_b_10;
input 	q_b_107;
input 	q_b_43;
input 	q_b_75;
input 	q_b_11;
input 	q_b_108;
input 	q_b_44;
input 	q_b_76;
input 	q_b_12;
input 	q_b_109;
input 	q_b_45;
input 	q_b_77;
input 	q_b_13;
input 	q_b_110;
input 	q_b_46;
input 	q_b_78;
input 	q_b_14;
input 	q_b_111;
input 	q_b_47;
input 	q_b_79;
input 	q_b_15;
input 	q_b_112;
input 	q_b_48;
input 	q_b_80;
input 	q_b_16;
input 	q_b_113;
input 	q_b_49;
input 	q_b_81;
input 	q_b_17;
input 	q_b_114;
input 	q_b_50;
input 	q_b_82;
input 	q_b_18;
input 	q_b_115;
input 	q_b_51;
input 	q_b_83;
input 	q_b_19;
input 	q_b_116;
input 	q_b_52;
input 	q_b_84;
input 	q_b_20;
input 	q_b_117;
input 	q_b_53;
input 	q_b_85;
input 	q_b_21;
input 	q_b_118;
input 	q_b_54;
input 	q_b_86;
input 	q_b_22;
input 	q_b_119;
input 	q_b_55;
input 	q_b_87;
input 	q_b_23;
input 	q_b_120;
input 	q_b_56;
input 	q_b_88;
input 	q_b_24;
input 	q_b_121;
input 	q_b_57;
input 	q_b_89;
input 	q_b_25;
input 	q_b_122;
input 	q_b_58;
input 	q_b_90;
input 	q_b_26;
input 	q_b_123;
input 	q_b_59;
input 	q_b_91;
input 	q_b_27;
input 	q_b_124;
input 	q_b_60;
input 	q_b_92;
input 	q_b_28;
input 	q_b_125;
input 	q_b_61;
input 	q_b_93;
input 	q_b_29;
input 	q_b_126;
input 	q_b_62;
input 	q_b_94;
input 	q_b_30;
input 	q_b_127;
input 	q_b_63;
input 	q_b_95;
input 	q_b_31;
input 	reset_phy_clk_1x_n;
input 	ctl_init_fail;
input 	ctl_init_success;
input 	reset_write_clk_2x_n;
output 	dqs_burst_2x_r3_0;
output 	dqs_burst_2x_r3_1;
output 	dqs_burst_2x_r3_2;
output 	dqs_burst_2x_r3_3;
input 	reset_mem_clk_2x_n;
input 	afi_dm_4;
input 	dgwb_wdp_ovride;
input 	seq_wdp_ovride;
input 	afi_dm_12;
input 	afi_dm_0;
input 	afi_dm_8;
input 	afi_dm_5;
input 	afi_dm_13;
input 	afi_dm_1;
input 	afi_dm_9;
input 	afi_dm_6;
input 	afi_dm_14;
input 	afi_dm_2;
input 	afi_dm_10;
input 	afi_dm_7;
input 	afi_dm_15;
input 	afi_dm_3;
input 	afi_dm_11;
input 	int_wdata_valid;
input 	dgwb_wdata_120;
input 	dgwb_wdata_56;
input 	dgwb_wdata_88;
input 	dgwb_wdata_24;
input 	dgwb_wdata_121;
input 	dgwb_wdata_57;
input 	dgwb_wdata_89;
input 	dgwb_wdata_25;
input 	dgwb_wdata_122;
input 	dgwb_wdata_58;
input 	dgwb_wdata_90;
input 	dgwb_wdata_26;
input 	dgwb_wdata_123;
input 	dgwb_wdata_59;
input 	dgwb_wdata_91;
input 	dgwb_wdata_27;
input 	dgwb_wdata_124;
input 	dgwb_wdata_60;
input 	dgwb_wdata_92;
input 	dgwb_wdata_28;
input 	dgwb_wdata_125;
input 	dgwb_wdata_61;
input 	dgwb_wdata_93;
input 	dgwb_wdata_29;
input 	dgwb_wdata_126;
input 	dgwb_wdata_62;
input 	dgwb_wdata_94;
input 	dgwb_wdata_30;
input 	dgwb_wdata_127;
input 	dgwb_wdata_63;
input 	dgwb_wdata_95;
input 	dgwb_wdata_31;
input 	int_dqs_burst;
input 	int_dqs_burst_hr;
input 	dgwb_wdp_ovride1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \dqs_burst_sel[0]~q ;
wire \dqs_burst_sel[1]~q ;
wire \dqs_burst_sel[2]~q ;
wire \dqs_burst_sel[3]~q ;
wire \dqs_burst2_2x_r2[0]~q ;
wire \dqs_burst2_2x_r3[0]~q ;
wire \dqs_burst_sel~0_combout ;
wire \dqs_burst2_2x_r2[1]~q ;
wire \dqs_burst2_2x_r3[1]~q ;
wire \dqs_burst_sel~1_combout ;
wire \dqs_burst2_2x_r2[2]~q ;
wire \dqs_burst2_2x_r3[2]~q ;
wire \dqs_burst_sel~2_combout ;
wire \dqs_burst2_2x_r2[3]~q ;
wire \dqs_burst2_2x_r3[3]~q ;
wire \dqs_burst_sel~3_combout ;
wire \dqs_burst2_2x_r1[0]~q ;
wire \dqs_burst2_2x_r1[1]~q ;
wire \dqs_burst2_2x_r1[2]~q ;
wire \dqs_burst2_2x_r1[3]~q ;
wire \dqs_burst2_1x_r[0]~q ;
wire \dqs_burst2_1x_r[1]~q ;
wire \dqs_burst2_1x_r[2]~q ;
wire \dqs_burst2_1x_r[3]~q ;
wire \mem_dm_r1[4]~q ;
wire \mem_dm_r2[4]~q ;
wire \mem_dm_r1[12]~q ;
wire \mem_dm_r2[12]~q ;
wire \mem_wdata_valid[0]~0_combout ;
wire \wdata_dm_1x_r~q ;
wire \wdata_dm_2x_r1~q ;
wire \wdata_dm_2x_r2~q ;
wire \dm_sel~0_combout ;
wire \dm_sel~q ;
wire \mem_dm_r1[0]~q ;
wire \mem_dm_r2[0]~q ;
wire \mem_dm_r1[8]~q ;
wire \mem_dm_r2[8]~q ;
wire \mem_dm_r1[5]~q ;
wire \mem_dm_r2[5]~q ;
wire \mem_dm_r1[13]~q ;
wire \mem_dm_r2[13]~q ;
wire \mem_dm_r1[1]~q ;
wire \mem_dm_r2[1]~q ;
wire \mem_dm_r1[9]~q ;
wire \mem_dm_r2[9]~q ;
wire \mem_dm_r1[6]~q ;
wire \mem_dm_r2[6]~q ;
wire \mem_dm_r1[14]~q ;
wire \mem_dm_r2[14]~q ;
wire \mem_dm_r1[2]~q ;
wire \mem_dm_r2[2]~q ;
wire \mem_dm_r1[10]~q ;
wire \mem_dm_r2[10]~q ;
wire \mem_dm_r1[7]~q ;
wire \mem_dm_r2[7]~q ;
wire \mem_dm_r1[15]~q ;
wire \mem_dm_r2[15]~q ;
wire \mem_dm_r1[3]~q ;
wire \mem_dm_r2[3]~q ;
wire \mem_dm_r1[11]~q ;
wire \mem_dm_r2[11]~q ;
wire \mem_wdata[96]~0_combout ;
wire \mem_wdata_r1[96]~q ;
wire \mem_wdata_r2[96]~q ;
wire \mem_wdata[32]~1_combout ;
wire \mem_wdata_r1[32]~q ;
wire \mem_wdata_r2[32]~q ;
wire \wdata_valid_1x_r[0]~q ;
wire \wdata_valid_2x_r1[0]~q ;
wire \wdata_valid_2x_r2[0]~q ;
wire \wdata_sel~0_combout ;
wire \wdata_sel[0]~q ;
wire \mem_wdata[64]~2_combout ;
wire \mem_wdata_r1[64]~q ;
wire \mem_wdata_r2[64]~q ;
wire \mem_wdata[0]~3_combout ;
wire \mem_wdata_r1[0]~q ;
wire \mem_wdata_r2[0]~q ;
wire \wdata_valid_1x_r1[8]~q ;
wire \wdata_valid_1x_r2[8]~q ;
wire \wdata_valid_1x_r1[0]~q ;
wire \wdata_valid_1x_r2[0]~q ;
wire \mem_wdata[97]~4_combout ;
wire \mem_wdata_r1[97]~q ;
wire \mem_wdata_r2[97]~q ;
wire \mem_wdata[33]~5_combout ;
wire \mem_wdata_r1[33]~q ;
wire \mem_wdata_r2[33]~q ;
wire \mem_wdata[65]~6_combout ;
wire \mem_wdata_r1[65]~q ;
wire \mem_wdata_r2[65]~q ;
wire \mem_wdata[1]~7_combout ;
wire \mem_wdata_r1[1]~q ;
wire \mem_wdata_r2[1]~q ;
wire \mem_wdata[98]~8_combout ;
wire \mem_wdata_r1[98]~q ;
wire \mem_wdata_r2[98]~q ;
wire \mem_wdata[34]~9_combout ;
wire \mem_wdata_r1[34]~q ;
wire \mem_wdata_r2[34]~q ;
wire \mem_wdata[66]~10_combout ;
wire \mem_wdata_r1[66]~q ;
wire \mem_wdata_r2[66]~q ;
wire \mem_wdata[2]~11_combout ;
wire \mem_wdata_r1[2]~q ;
wire \mem_wdata_r2[2]~q ;
wire \mem_wdata[99]~12_combout ;
wire \mem_wdata_r1[99]~q ;
wire \mem_wdata_r2[99]~q ;
wire \mem_wdata[35]~13_combout ;
wire \mem_wdata_r1[35]~q ;
wire \mem_wdata_r2[35]~q ;
wire \mem_wdata[67]~14_combout ;
wire \mem_wdata_r1[67]~q ;
wire \mem_wdata_r2[67]~q ;
wire \mem_wdata[3]~15_combout ;
wire \mem_wdata_r1[3]~q ;
wire \mem_wdata_r2[3]~q ;
wire \mem_wdata[100]~16_combout ;
wire \mem_wdata_r1[100]~q ;
wire \mem_wdata_r2[100]~q ;
wire \mem_wdata[36]~17_combout ;
wire \mem_wdata_r1[36]~q ;
wire \mem_wdata_r2[36]~q ;
wire \wdata_valid_1x_r[1]~q ;
wire \wdata_valid_2x_r1[1]~q ;
wire \wdata_valid_2x_r2[1]~q ;
wire \wdata_sel~1_combout ;
wire \wdata_sel[1]~q ;
wire \mem_wdata[68]~18_combout ;
wire \mem_wdata_r1[68]~q ;
wire \mem_wdata_r2[68]~q ;
wire \mem_wdata[4]~19_combout ;
wire \mem_wdata_r1[4]~q ;
wire \mem_wdata_r2[4]~q ;
wire \wdata_valid_1x_r1[9]~q ;
wire \wdata_valid_1x_r2[9]~q ;
wire \wdata_valid_1x_r1[1]~q ;
wire \wdata_valid_1x_r2[1]~q ;
wire \mem_wdata[101]~20_combout ;
wire \mem_wdata_r1[101]~q ;
wire \mem_wdata_r2[101]~q ;
wire \mem_wdata[37]~21_combout ;
wire \mem_wdata_r1[37]~q ;
wire \mem_wdata_r2[37]~q ;
wire \mem_wdata[69]~22_combout ;
wire \mem_wdata_r1[69]~q ;
wire \mem_wdata_r2[69]~q ;
wire \mem_wdata[5]~23_combout ;
wire \mem_wdata_r1[5]~q ;
wire \mem_wdata_r2[5]~q ;
wire \mem_wdata[102]~24_combout ;
wire \mem_wdata_r1[102]~q ;
wire \mem_wdata_r2[102]~q ;
wire \mem_wdata[38]~25_combout ;
wire \mem_wdata_r1[38]~q ;
wire \mem_wdata_r2[38]~q ;
wire \mem_wdata[70]~26_combout ;
wire \mem_wdata_r1[70]~q ;
wire \mem_wdata_r2[70]~q ;
wire \mem_wdata[6]~27_combout ;
wire \mem_wdata_r1[6]~q ;
wire \mem_wdata_r2[6]~q ;
wire \mem_wdata[103]~28_combout ;
wire \mem_wdata_r1[103]~q ;
wire \mem_wdata_r2[103]~q ;
wire \mem_wdata[39]~29_combout ;
wire \mem_wdata_r1[39]~q ;
wire \mem_wdata_r2[39]~q ;
wire \mem_wdata[71]~30_combout ;
wire \mem_wdata_r1[71]~q ;
wire \mem_wdata_r2[71]~q ;
wire \mem_wdata[7]~31_combout ;
wire \mem_wdata_r1[7]~q ;
wire \mem_wdata_r2[7]~q ;
wire \mem_wdata[104]~32_combout ;
wire \mem_wdata_r1[104]~q ;
wire \mem_wdata_r2[104]~q ;
wire \mem_wdata[40]~33_combout ;
wire \mem_wdata_r1[40]~q ;
wire \mem_wdata_r2[40]~q ;
wire \wdata_valid_1x_r[2]~q ;
wire \wdata_valid_2x_r1[2]~q ;
wire \wdata_valid_2x_r2[2]~q ;
wire \wdata_sel~2_combout ;
wire \wdata_sel[2]~q ;
wire \mem_wdata[72]~34_combout ;
wire \mem_wdata_r1[72]~q ;
wire \mem_wdata_r2[72]~q ;
wire \mem_wdata[8]~35_combout ;
wire \mem_wdata_r1[8]~q ;
wire \mem_wdata_r2[8]~q ;
wire \wdata_valid_1x_r1[10]~q ;
wire \wdata_valid_1x_r2[10]~q ;
wire \wdata_valid_1x_r1[2]~q ;
wire \wdata_valid_1x_r2[2]~q ;
wire \mem_wdata[105]~36_combout ;
wire \mem_wdata_r1[105]~q ;
wire \mem_wdata_r2[105]~q ;
wire \mem_wdata[41]~37_combout ;
wire \mem_wdata_r1[41]~q ;
wire \mem_wdata_r2[41]~q ;
wire \mem_wdata[73]~38_combout ;
wire \mem_wdata_r1[73]~q ;
wire \mem_wdata_r2[73]~q ;
wire \mem_wdata[9]~39_combout ;
wire \mem_wdata_r1[9]~q ;
wire \mem_wdata_r2[9]~q ;
wire \mem_wdata[106]~40_combout ;
wire \mem_wdata_r1[106]~q ;
wire \mem_wdata_r2[106]~q ;
wire \mem_wdata[42]~41_combout ;
wire \mem_wdata_r1[42]~q ;
wire \mem_wdata_r2[42]~q ;
wire \mem_wdata[74]~42_combout ;
wire \mem_wdata_r1[74]~q ;
wire \mem_wdata_r2[74]~q ;
wire \mem_wdata[10]~43_combout ;
wire \mem_wdata_r1[10]~q ;
wire \mem_wdata_r2[10]~q ;
wire \mem_wdata[107]~44_combout ;
wire \mem_wdata_r1[107]~q ;
wire \mem_wdata_r2[107]~q ;
wire \mem_wdata[43]~45_combout ;
wire \mem_wdata_r1[43]~q ;
wire \mem_wdata_r2[43]~q ;
wire \mem_wdata[75]~46_combout ;
wire \mem_wdata_r1[75]~q ;
wire \mem_wdata_r2[75]~q ;
wire \mem_wdata[11]~47_combout ;
wire \mem_wdata_r1[11]~q ;
wire \mem_wdata_r2[11]~q ;
wire \mem_wdata[108]~48_combout ;
wire \mem_wdata_r1[108]~q ;
wire \mem_wdata_r2[108]~q ;
wire \mem_wdata[44]~49_combout ;
wire \mem_wdata_r1[44]~q ;
wire \mem_wdata_r2[44]~q ;
wire \wdata_valid_1x_r[3]~q ;
wire \wdata_valid_2x_r1[3]~q ;
wire \wdata_valid_2x_r2[3]~q ;
wire \wdata_sel~3_combout ;
wire \wdata_sel[3]~q ;
wire \mem_wdata[76]~50_combout ;
wire \mem_wdata_r1[76]~q ;
wire \mem_wdata_r2[76]~q ;
wire \mem_wdata[12]~51_combout ;
wire \mem_wdata_r1[12]~q ;
wire \mem_wdata_r2[12]~q ;
wire \wdata_valid_1x_r1[11]~q ;
wire \wdata_valid_1x_r2[11]~q ;
wire \wdata_valid_1x_r1[3]~q ;
wire \wdata_valid_1x_r2[3]~q ;
wire \mem_wdata[109]~52_combout ;
wire \mem_wdata_r1[109]~q ;
wire \mem_wdata_r2[109]~q ;
wire \mem_wdata[45]~53_combout ;
wire \mem_wdata_r1[45]~q ;
wire \mem_wdata_r2[45]~q ;
wire \mem_wdata[77]~54_combout ;
wire \mem_wdata_r1[77]~q ;
wire \mem_wdata_r2[77]~q ;
wire \mem_wdata[13]~55_combout ;
wire \mem_wdata_r1[13]~q ;
wire \mem_wdata_r2[13]~q ;
wire \mem_wdata[110]~56_combout ;
wire \mem_wdata_r1[110]~q ;
wire \mem_wdata_r2[110]~q ;
wire \mem_wdata[46]~57_combout ;
wire \mem_wdata_r1[46]~q ;
wire \mem_wdata_r2[46]~q ;
wire \mem_wdata[78]~58_combout ;
wire \mem_wdata_r1[78]~q ;
wire \mem_wdata_r2[78]~q ;
wire \mem_wdata[14]~59_combout ;
wire \mem_wdata_r1[14]~q ;
wire \mem_wdata_r2[14]~q ;
wire \mem_wdata[111]~60_combout ;
wire \mem_wdata_r1[111]~q ;
wire \mem_wdata_r2[111]~q ;
wire \mem_wdata[47]~61_combout ;
wire \mem_wdata_r1[47]~q ;
wire \mem_wdata_r2[47]~q ;
wire \mem_wdata[79]~62_combout ;
wire \mem_wdata_r1[79]~q ;
wire \mem_wdata_r2[79]~q ;
wire \mem_wdata[15]~63_combout ;
wire \mem_wdata_r1[15]~q ;
wire \mem_wdata_r2[15]~q ;
wire \mem_wdata[112]~64_combout ;
wire \mem_wdata_r1[112]~q ;
wire \mem_wdata_r2[112]~q ;
wire \mem_wdata[48]~65_combout ;
wire \mem_wdata_r1[48]~q ;
wire \mem_wdata_r2[48]~q ;
wire \wdata_valid_1x_r[4]~q ;
wire \wdata_valid_2x_r1[4]~q ;
wire \wdata_valid_2x_r2[4]~q ;
wire \wdata_sel~4_combout ;
wire \wdata_sel[4]~q ;
wire \mem_wdata[80]~66_combout ;
wire \mem_wdata_r1[80]~q ;
wire \mem_wdata_r2[80]~q ;
wire \mem_wdata[16]~67_combout ;
wire \mem_wdata_r1[16]~q ;
wire \mem_wdata_r2[16]~q ;
wire \wdata_valid_1x_r1[12]~q ;
wire \wdata_valid_1x_r2[12]~q ;
wire \wdata_valid_1x_r1[4]~q ;
wire \wdata_valid_1x_r2[4]~q ;
wire \mem_wdata[113]~68_combout ;
wire \mem_wdata_r1[113]~q ;
wire \mem_wdata_r2[113]~q ;
wire \mem_wdata[49]~69_combout ;
wire \mem_wdata_r1[49]~q ;
wire \mem_wdata_r2[49]~q ;
wire \mem_wdata[81]~70_combout ;
wire \mem_wdata_r1[81]~q ;
wire \mem_wdata_r2[81]~q ;
wire \mem_wdata[17]~71_combout ;
wire \mem_wdata_r1[17]~q ;
wire \mem_wdata_r2[17]~q ;
wire \mem_wdata[114]~72_combout ;
wire \mem_wdata_r1[114]~q ;
wire \mem_wdata_r2[114]~q ;
wire \mem_wdata[50]~73_combout ;
wire \mem_wdata_r1[50]~q ;
wire \mem_wdata_r2[50]~q ;
wire \mem_wdata[82]~74_combout ;
wire \mem_wdata_r1[82]~q ;
wire \mem_wdata_r2[82]~q ;
wire \mem_wdata[18]~75_combout ;
wire \mem_wdata_r1[18]~q ;
wire \mem_wdata_r2[18]~q ;
wire \mem_wdata[115]~76_combout ;
wire \mem_wdata_r1[115]~q ;
wire \mem_wdata_r2[115]~q ;
wire \mem_wdata[51]~77_combout ;
wire \mem_wdata_r1[51]~q ;
wire \mem_wdata_r2[51]~q ;
wire \mem_wdata[83]~78_combout ;
wire \mem_wdata_r1[83]~q ;
wire \mem_wdata_r2[83]~q ;
wire \mem_wdata[19]~79_combout ;
wire \mem_wdata_r1[19]~q ;
wire \mem_wdata_r2[19]~q ;
wire \mem_wdata[116]~80_combout ;
wire \mem_wdata_r1[116]~q ;
wire \mem_wdata_r2[116]~q ;
wire \mem_wdata[52]~81_combout ;
wire \mem_wdata_r1[52]~q ;
wire \mem_wdata_r2[52]~q ;
wire \wdata_valid_1x_r[5]~q ;
wire \wdata_valid_2x_r1[5]~q ;
wire \wdata_valid_2x_r2[5]~q ;
wire \wdata_sel~5_combout ;
wire \wdata_sel[5]~q ;
wire \mem_wdata[84]~82_combout ;
wire \mem_wdata_r1[84]~q ;
wire \mem_wdata_r2[84]~q ;
wire \mem_wdata[20]~83_combout ;
wire \mem_wdata_r1[20]~q ;
wire \mem_wdata_r2[20]~q ;
wire \wdata_valid_1x_r1[13]~q ;
wire \wdata_valid_1x_r2[13]~q ;
wire \wdata_valid_1x_r1[5]~q ;
wire \wdata_valid_1x_r2[5]~q ;
wire \mem_wdata[117]~84_combout ;
wire \mem_wdata_r1[117]~q ;
wire \mem_wdata_r2[117]~q ;
wire \mem_wdata[53]~85_combout ;
wire \mem_wdata_r1[53]~q ;
wire \mem_wdata_r2[53]~q ;
wire \mem_wdata[85]~86_combout ;
wire \mem_wdata_r1[85]~q ;
wire \mem_wdata_r2[85]~q ;
wire \mem_wdata[21]~87_combout ;
wire \mem_wdata_r1[21]~q ;
wire \mem_wdata_r2[21]~q ;
wire \mem_wdata[118]~88_combout ;
wire \mem_wdata_r1[118]~q ;
wire \mem_wdata_r2[118]~q ;
wire \mem_wdata[54]~89_combout ;
wire \mem_wdata_r1[54]~q ;
wire \mem_wdata_r2[54]~q ;
wire \mem_wdata[86]~90_combout ;
wire \mem_wdata_r1[86]~q ;
wire \mem_wdata_r2[86]~q ;
wire \mem_wdata[22]~91_combout ;
wire \mem_wdata_r1[22]~q ;
wire \mem_wdata_r2[22]~q ;
wire \mem_wdata[119]~92_combout ;
wire \mem_wdata_r1[119]~q ;
wire \mem_wdata_r2[119]~q ;
wire \mem_wdata[55]~93_combout ;
wire \mem_wdata_r1[55]~q ;
wire \mem_wdata_r2[55]~q ;
wire \mem_wdata[87]~94_combout ;
wire \mem_wdata_r1[87]~q ;
wire \mem_wdata_r2[87]~q ;
wire \mem_wdata[23]~95_combout ;
wire \mem_wdata_r1[23]~q ;
wire \mem_wdata_r2[23]~q ;
wire \mem_wdata[120]~96_combout ;
wire \mem_wdata_r1[120]~q ;
wire \mem_wdata_r2[120]~q ;
wire \mem_wdata[56]~97_combout ;
wire \mem_wdata_r1[56]~q ;
wire \mem_wdata_r2[56]~q ;
wire \wdata_valid_1x_r[6]~q ;
wire \wdata_valid_2x_r1[6]~q ;
wire \wdata_valid_2x_r2[6]~q ;
wire \wdata_sel~6_combout ;
wire \wdata_sel[6]~q ;
wire \mem_wdata[88]~98_combout ;
wire \mem_wdata_r1[88]~q ;
wire \mem_wdata_r2[88]~q ;
wire \mem_wdata[24]~99_combout ;
wire \mem_wdata_r1[24]~q ;
wire \mem_wdata_r2[24]~q ;
wire \wdata_valid_1x_r1[14]~q ;
wire \wdata_valid_1x_r2[14]~q ;
wire \wdata_valid_1x_r1[6]~q ;
wire \wdata_valid_1x_r2[6]~q ;
wire \mem_wdata[121]~100_combout ;
wire \mem_wdata_r1[121]~q ;
wire \mem_wdata_r2[121]~q ;
wire \mem_wdata[57]~101_combout ;
wire \mem_wdata_r1[57]~q ;
wire \mem_wdata_r2[57]~q ;
wire \mem_wdata[89]~102_combout ;
wire \mem_wdata_r1[89]~q ;
wire \mem_wdata_r2[89]~q ;
wire \mem_wdata[25]~103_combout ;
wire \mem_wdata_r1[25]~q ;
wire \mem_wdata_r2[25]~q ;
wire \mem_wdata[122]~104_combout ;
wire \mem_wdata_r1[122]~q ;
wire \mem_wdata_r2[122]~q ;
wire \mem_wdata[58]~105_combout ;
wire \mem_wdata_r1[58]~q ;
wire \mem_wdata_r2[58]~q ;
wire \mem_wdata[90]~106_combout ;
wire \mem_wdata_r1[90]~q ;
wire \mem_wdata_r2[90]~q ;
wire \mem_wdata[26]~107_combout ;
wire \mem_wdata_r1[26]~q ;
wire \mem_wdata_r2[26]~q ;
wire \mem_wdata[123]~108_combout ;
wire \mem_wdata_r1[123]~q ;
wire \mem_wdata_r2[123]~q ;
wire \mem_wdata[59]~109_combout ;
wire \mem_wdata_r1[59]~q ;
wire \mem_wdata_r2[59]~q ;
wire \mem_wdata[91]~110_combout ;
wire \mem_wdata_r1[91]~q ;
wire \mem_wdata_r2[91]~q ;
wire \mem_wdata[27]~111_combout ;
wire \mem_wdata_r1[27]~q ;
wire \mem_wdata_r2[27]~q ;
wire \mem_wdata[124]~112_combout ;
wire \mem_wdata_r1[124]~q ;
wire \mem_wdata_r2[124]~q ;
wire \mem_wdata[60]~113_combout ;
wire \mem_wdata_r1[60]~q ;
wire \mem_wdata_r2[60]~q ;
wire \wdata_valid_1x_r[7]~q ;
wire \wdata_valid_2x_r1[7]~q ;
wire \wdata_valid_2x_r2[7]~q ;
wire \wdata_sel~7_combout ;
wire \wdata_sel[7]~q ;
wire \mem_wdata[92]~114_combout ;
wire \mem_wdata_r1[92]~q ;
wire \mem_wdata_r2[92]~q ;
wire \mem_wdata[28]~115_combout ;
wire \mem_wdata_r1[28]~q ;
wire \mem_wdata_r2[28]~q ;
wire \wdata_valid_1x_r1[15]~q ;
wire \wdata_valid_1x_r2[15]~q ;
wire \wdata_valid_1x_r1[7]~q ;
wire \wdata_valid_1x_r2[7]~q ;
wire \mem_wdata[125]~116_combout ;
wire \mem_wdata_r1[125]~q ;
wire \mem_wdata_r2[125]~q ;
wire \mem_wdata[61]~117_combout ;
wire \mem_wdata_r1[61]~q ;
wire \mem_wdata_r2[61]~q ;
wire \mem_wdata[93]~118_combout ;
wire \mem_wdata_r1[93]~q ;
wire \mem_wdata_r2[93]~q ;
wire \mem_wdata[29]~119_combout ;
wire \mem_wdata_r1[29]~q ;
wire \mem_wdata_r2[29]~q ;
wire \mem_wdata[126]~120_combout ;
wire \mem_wdata_r1[126]~q ;
wire \mem_wdata_r2[126]~q ;
wire \mem_wdata[62]~121_combout ;
wire \mem_wdata_r1[62]~q ;
wire \mem_wdata_r2[62]~q ;
wire \mem_wdata[94]~122_combout ;
wire \mem_wdata_r1[94]~q ;
wire \mem_wdata_r2[94]~q ;
wire \mem_wdata[30]~123_combout ;
wire \mem_wdata_r1[30]~q ;
wire \mem_wdata_r2[30]~q ;
wire \mem_wdata[127]~124_combout ;
wire \mem_wdata_r1[127]~q ;
wire \mem_wdata_r2[127]~q ;
wire \mem_wdata[63]~125_combout ;
wire \mem_wdata_r1[63]~q ;
wire \mem_wdata_r2[63]~q ;
wire \mem_wdata[95]~126_combout ;
wire \mem_wdata_r1[95]~q ;
wire \mem_wdata_r2[95]~q ;
wire \mem_wdata[31]~127_combout ;
wire \mem_wdata_r1[31]~q ;
wire \mem_wdata_r2[31]~q ;
wire \mem_dqs_burst[4]~0_combout ;
wire \dqs_burst_1x_r[4]~q ;
wire \dqs_burst_2x_r1[4]~q ;
wire \mem_dqs_burst[0]~1_combout ;
wire \dqs_burst_1x_r[0]~q ;
wire \dqs_burst_2x_r1[0]~q ;
wire \dqs_burst_2x_r2~0_combout ;
wire \dqs_burst_2x_r2[0]~q ;
wire \dqs_burst_1x_r[5]~q ;
wire \dqs_burst_2x_r1[5]~q ;
wire \dqs_burst_1x_r[1]~q ;
wire \dqs_burst_2x_r1[1]~q ;
wire \dqs_burst_2x_r2~1_combout ;
wire \dqs_burst_2x_r2[1]~q ;
wire \dqs_burst_1x_r[6]~q ;
wire \dqs_burst_2x_r1[6]~q ;
wire \dqs_burst_1x_r[2]~q ;
wire \dqs_burst_2x_r1[2]~q ;
wire \dqs_burst_2x_r2~2_combout ;
wire \dqs_burst_2x_r2[2]~q ;
wire \dqs_burst_1x_r[7]~q ;
wire \dqs_burst_2x_r1[7]~q ;
wire \dqs_burst_1x_r[3]~q ;
wire \dqs_burst_2x_r1[3]~q ;
wire \dqs_burst_2x_r2~3_combout ;
wire \dqs_burst_2x_r2[3]~q ;


dffeas \dqs_burst_sel[0] (
	.clk(mem_clk_2x),
	.d(\dqs_burst_sel~0_combout ),
	.asdata(vcc),
	.clrn(reset_mem_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst_sel[0]~q ),
	.prn(vcc));
defparam \dqs_burst_sel[0] .is_wysiwyg = "true";
defparam \dqs_burst_sel[0] .power_up = "low";

dffeas \dqs_burst_sel[1] (
	.clk(mem_clk_2x),
	.d(\dqs_burst_sel~1_combout ),
	.asdata(vcc),
	.clrn(reset_mem_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst_sel[1]~q ),
	.prn(vcc));
defparam \dqs_burst_sel[1] .is_wysiwyg = "true";
defparam \dqs_burst_sel[1] .power_up = "low";

dffeas \dqs_burst_sel[2] (
	.clk(mem_clk_2x),
	.d(\dqs_burst_sel~2_combout ),
	.asdata(vcc),
	.clrn(reset_mem_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst_sel[2]~q ),
	.prn(vcc));
defparam \dqs_burst_sel[2] .is_wysiwyg = "true";
defparam \dqs_burst_sel[2] .power_up = "low";

dffeas \dqs_burst_sel[3] (
	.clk(mem_clk_2x),
	.d(\dqs_burst_sel~3_combout ),
	.asdata(vcc),
	.clrn(reset_mem_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst_sel[3]~q ),
	.prn(vcc));
defparam \dqs_burst_sel[3] .is_wysiwyg = "true";
defparam \dqs_burst_sel[3] .power_up = "low";

dffeas \dqs_burst2_2x_r2[0] (
	.clk(mem_clk_2x),
	.d(\dqs_burst2_2x_r1[0]~q ),
	.asdata(vcc),
	.clrn(reset_mem_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst2_2x_r2[0]~q ),
	.prn(vcc));
defparam \dqs_burst2_2x_r2[0] .is_wysiwyg = "true";
defparam \dqs_burst2_2x_r2[0] .power_up = "low";

dffeas \dqs_burst2_2x_r3[0] (
	.clk(mem_clk_2x),
	.d(\dqs_burst2_2x_r2[0]~q ),
	.asdata(vcc),
	.clrn(reset_mem_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst2_2x_r3[0]~q ),
	.prn(vcc));
defparam \dqs_burst2_2x_r3[0] .is_wysiwyg = "true";
defparam \dqs_burst2_2x_r3[0] .power_up = "low";

arriaii_lcell_comb \dqs_burst_sel~0 (
	.dataa(!\dqs_burst_sel[0]~q ),
	.datab(!\dqs_burst2_2x_r2[0]~q ),
	.datac(!\dqs_burst2_2x_r3[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dqs_burst_sel~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dqs_burst_sel~0 .extended_lut = "off";
defparam \dqs_burst_sel~0 .lut_mask = 64'h8A8A8A8A8A8A8A8A;
defparam \dqs_burst_sel~0 .shared_arith = "off";

dffeas \dqs_burst2_2x_r2[1] (
	.clk(mem_clk_2x),
	.d(\dqs_burst2_2x_r1[1]~q ),
	.asdata(vcc),
	.clrn(reset_mem_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst2_2x_r2[1]~q ),
	.prn(vcc));
defparam \dqs_burst2_2x_r2[1] .is_wysiwyg = "true";
defparam \dqs_burst2_2x_r2[1] .power_up = "low";

dffeas \dqs_burst2_2x_r3[1] (
	.clk(mem_clk_2x),
	.d(\dqs_burst2_2x_r2[1]~q ),
	.asdata(vcc),
	.clrn(reset_mem_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst2_2x_r3[1]~q ),
	.prn(vcc));
defparam \dqs_burst2_2x_r3[1] .is_wysiwyg = "true";
defparam \dqs_burst2_2x_r3[1] .power_up = "low";

arriaii_lcell_comb \dqs_burst_sel~1 (
	.dataa(!\dqs_burst_sel[1]~q ),
	.datab(!\dqs_burst2_2x_r2[1]~q ),
	.datac(!\dqs_burst2_2x_r3[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dqs_burst_sel~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dqs_burst_sel~1 .extended_lut = "off";
defparam \dqs_burst_sel~1 .lut_mask = 64'h8A8A8A8A8A8A8A8A;
defparam \dqs_burst_sel~1 .shared_arith = "off";

dffeas \dqs_burst2_2x_r2[2] (
	.clk(mem_clk_2x),
	.d(\dqs_burst2_2x_r1[2]~q ),
	.asdata(vcc),
	.clrn(reset_mem_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst2_2x_r2[2]~q ),
	.prn(vcc));
defparam \dqs_burst2_2x_r2[2] .is_wysiwyg = "true";
defparam \dqs_burst2_2x_r2[2] .power_up = "low";

dffeas \dqs_burst2_2x_r3[2] (
	.clk(mem_clk_2x),
	.d(\dqs_burst2_2x_r2[2]~q ),
	.asdata(vcc),
	.clrn(reset_mem_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst2_2x_r3[2]~q ),
	.prn(vcc));
defparam \dqs_burst2_2x_r3[2] .is_wysiwyg = "true";
defparam \dqs_burst2_2x_r3[2] .power_up = "low";

arriaii_lcell_comb \dqs_burst_sel~2 (
	.dataa(!\dqs_burst_sel[2]~q ),
	.datab(!\dqs_burst2_2x_r2[2]~q ),
	.datac(!\dqs_burst2_2x_r3[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dqs_burst_sel~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dqs_burst_sel~2 .extended_lut = "off";
defparam \dqs_burst_sel~2 .lut_mask = 64'h8A8A8A8A8A8A8A8A;
defparam \dqs_burst_sel~2 .shared_arith = "off";

dffeas \dqs_burst2_2x_r2[3] (
	.clk(mem_clk_2x),
	.d(\dqs_burst2_2x_r1[3]~q ),
	.asdata(vcc),
	.clrn(reset_mem_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst2_2x_r2[3]~q ),
	.prn(vcc));
defparam \dqs_burst2_2x_r2[3] .is_wysiwyg = "true";
defparam \dqs_burst2_2x_r2[3] .power_up = "low";

dffeas \dqs_burst2_2x_r3[3] (
	.clk(mem_clk_2x),
	.d(\dqs_burst2_2x_r2[3]~q ),
	.asdata(vcc),
	.clrn(reset_mem_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst2_2x_r3[3]~q ),
	.prn(vcc));
defparam \dqs_burst2_2x_r3[3] .is_wysiwyg = "true";
defparam \dqs_burst2_2x_r3[3] .power_up = "low";

arriaii_lcell_comb \dqs_burst_sel~3 (
	.dataa(!\dqs_burst_sel[3]~q ),
	.datab(!\dqs_burst2_2x_r2[3]~q ),
	.datac(!\dqs_burst2_2x_r3[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dqs_burst_sel~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dqs_burst_sel~3 .extended_lut = "off";
defparam \dqs_burst_sel~3 .lut_mask = 64'h8A8A8A8A8A8A8A8A;
defparam \dqs_burst_sel~3 .shared_arith = "off";

dffeas \dqs_burst2_2x_r1[0] (
	.clk(mem_clk_2x),
	.d(\dqs_burst2_1x_r[0]~q ),
	.asdata(vcc),
	.clrn(reset_mem_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst2_2x_r1[0]~q ),
	.prn(vcc));
defparam \dqs_burst2_2x_r1[0] .is_wysiwyg = "true";
defparam \dqs_burst2_2x_r1[0] .power_up = "low";

dffeas \dqs_burst2_2x_r1[1] (
	.clk(mem_clk_2x),
	.d(\dqs_burst2_1x_r[1]~q ),
	.asdata(vcc),
	.clrn(reset_mem_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst2_2x_r1[1]~q ),
	.prn(vcc));
defparam \dqs_burst2_2x_r1[1] .is_wysiwyg = "true";
defparam \dqs_burst2_2x_r1[1] .power_up = "low";

dffeas \dqs_burst2_2x_r1[2] (
	.clk(mem_clk_2x),
	.d(\dqs_burst2_1x_r[2]~q ),
	.asdata(vcc),
	.clrn(reset_mem_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst2_2x_r1[2]~q ),
	.prn(vcc));
defparam \dqs_burst2_2x_r1[2] .is_wysiwyg = "true";
defparam \dqs_burst2_2x_r1[2] .power_up = "low";

dffeas \dqs_burst2_2x_r1[3] (
	.clk(mem_clk_2x),
	.d(\dqs_burst2_1x_r[3]~q ),
	.asdata(vcc),
	.clrn(reset_mem_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst2_2x_r1[3]~q ),
	.prn(vcc));
defparam \dqs_burst2_2x_r1[3] .is_wysiwyg = "true";
defparam \dqs_burst2_2x_r1[3] .power_up = "low";

dffeas \dqs_burst2_1x_r[0] (
	.clk(phy_clk_1x),
	.d(\mem_dqs_burst[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst2_1x_r[0]~q ),
	.prn(vcc));
defparam \dqs_burst2_1x_r[0] .is_wysiwyg = "true";
defparam \dqs_burst2_1x_r[0] .power_up = "low";

dffeas \dqs_burst2_1x_r[1] (
	.clk(phy_clk_1x),
	.d(\mem_dqs_burst[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst2_1x_r[1]~q ),
	.prn(vcc));
defparam \dqs_burst2_1x_r[1] .is_wysiwyg = "true";
defparam \dqs_burst2_1x_r[1] .power_up = "low";

dffeas \dqs_burst2_1x_r[2] (
	.clk(phy_clk_1x),
	.d(\mem_dqs_burst[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst2_1x_r[2]~q ),
	.prn(vcc));
defparam \dqs_burst2_1x_r[2] .is_wysiwyg = "true";
defparam \dqs_burst2_1x_r[2] .power_up = "low";

dffeas \dqs_burst2_1x_r[3] (
	.clk(phy_clk_1x),
	.d(\mem_dqs_burst[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst2_1x_r[3]~q ),
	.prn(vcc));
defparam \dqs_burst2_1x_r[3] .is_wysiwyg = "true";
defparam \dqs_burst2_1x_r[3] .power_up = "low";

dffeas \wdp_dm_l_2x[0] (
	.clk(write_clk_2x),
	.d(\mem_dm_r2[4]~q ),
	.asdata(\mem_dm_r2[12]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\dm_sel~q ),
	.ena(vcc),
	.q(wdp_dm_l_2x_0),
	.prn(vcc));
defparam \wdp_dm_l_2x[0] .is_wysiwyg = "true";
defparam \wdp_dm_l_2x[0] .power_up = "low";

dffeas \wdp_dm_h_2x[0] (
	.clk(write_clk_2x),
	.d(\mem_dm_r2[0]~q ),
	.asdata(\mem_dm_r2[8]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\dm_sel~q ),
	.ena(vcc),
	.q(wdp_dm_h_2x_0),
	.prn(vcc));
defparam \wdp_dm_h_2x[0] .is_wysiwyg = "true";
defparam \wdp_dm_h_2x[0] .power_up = "low";

dffeas \wdp_dm_l_2x[1] (
	.clk(write_clk_2x),
	.d(\mem_dm_r2[5]~q ),
	.asdata(\mem_dm_r2[13]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\dm_sel~q ),
	.ena(vcc),
	.q(wdp_dm_l_2x_1),
	.prn(vcc));
defparam \wdp_dm_l_2x[1] .is_wysiwyg = "true";
defparam \wdp_dm_l_2x[1] .power_up = "low";

dffeas \wdp_dm_h_2x[1] (
	.clk(write_clk_2x),
	.d(\mem_dm_r2[1]~q ),
	.asdata(\mem_dm_r2[9]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\dm_sel~q ),
	.ena(vcc),
	.q(wdp_dm_h_2x_1),
	.prn(vcc));
defparam \wdp_dm_h_2x[1] .is_wysiwyg = "true";
defparam \wdp_dm_h_2x[1] .power_up = "low";

dffeas \wdp_dm_l_2x[2] (
	.clk(write_clk_2x),
	.d(\mem_dm_r2[6]~q ),
	.asdata(\mem_dm_r2[14]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\dm_sel~q ),
	.ena(vcc),
	.q(wdp_dm_l_2x_2),
	.prn(vcc));
defparam \wdp_dm_l_2x[2] .is_wysiwyg = "true";
defparam \wdp_dm_l_2x[2] .power_up = "low";

dffeas \wdp_dm_h_2x[2] (
	.clk(write_clk_2x),
	.d(\mem_dm_r2[2]~q ),
	.asdata(\mem_dm_r2[10]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\dm_sel~q ),
	.ena(vcc),
	.q(wdp_dm_h_2x_2),
	.prn(vcc));
defparam \wdp_dm_h_2x[2] .is_wysiwyg = "true";
defparam \wdp_dm_h_2x[2] .power_up = "low";

dffeas \wdp_dm_l_2x[3] (
	.clk(write_clk_2x),
	.d(\mem_dm_r2[7]~q ),
	.asdata(\mem_dm_r2[15]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\dm_sel~q ),
	.ena(vcc),
	.q(wdp_dm_l_2x_3),
	.prn(vcc));
defparam \wdp_dm_l_2x[3] .is_wysiwyg = "true";
defparam \wdp_dm_l_2x[3] .power_up = "low";

dffeas \wdp_dm_h_2x[3] (
	.clk(write_clk_2x),
	.d(\mem_dm_r2[3]~q ),
	.asdata(\mem_dm_r2[11]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\dm_sel~q ),
	.ena(vcc),
	.q(wdp_dm_h_2x_3),
	.prn(vcc));
defparam \wdp_dm_h_2x[3] .is_wysiwyg = "true";
defparam \wdp_dm_h_2x[3] .power_up = "low";

dffeas \wdp_wdata_l_2x[0] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[96]~q ),
	.asdata(\mem_wdata_r2[32]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[0]~q ),
	.ena(vcc),
	.q(wdp_wdata_l_2x_0),
	.prn(vcc));
defparam \wdp_wdata_l_2x[0] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[0] .power_up = "low";

dffeas \wdp_wdata_h_2x[0] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[64]~q ),
	.asdata(\mem_wdata_r2[0]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[0]~q ),
	.ena(vcc),
	.q(wdp_wdata_h_2x_0),
	.prn(vcc));
defparam \wdp_wdata_h_2x[0] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[0] .power_up = "low";

dffeas \dq_oe_2x[0] (
	.clk(write_clk_2x),
	.d(\wdata_valid_1x_r2[8]~q ),
	.asdata(\wdata_valid_1x_r2[0]~q ),
	.clrn(reset_write_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[0]~q ),
	.ena(vcc),
	.q(dq_oe_2x_0),
	.prn(vcc));
defparam \dq_oe_2x[0] .is_wysiwyg = "true";
defparam \dq_oe_2x[0] .power_up = "low";

dffeas \wdp_wdata_l_2x[1] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[97]~q ),
	.asdata(\mem_wdata_r2[33]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[0]~q ),
	.ena(vcc),
	.q(wdp_wdata_l_2x_1),
	.prn(vcc));
defparam \wdp_wdata_l_2x[1] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[1] .power_up = "low";

dffeas \wdp_wdata_h_2x[1] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[65]~q ),
	.asdata(\mem_wdata_r2[1]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[0]~q ),
	.ena(vcc),
	.q(wdp_wdata_h_2x_1),
	.prn(vcc));
defparam \wdp_wdata_h_2x[1] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[1] .power_up = "low";

dffeas \wdp_wdata_l_2x[2] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[98]~q ),
	.asdata(\mem_wdata_r2[34]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[0]~q ),
	.ena(vcc),
	.q(wdp_wdata_l_2x_2),
	.prn(vcc));
defparam \wdp_wdata_l_2x[2] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[2] .power_up = "low";

dffeas \wdp_wdata_h_2x[2] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[66]~q ),
	.asdata(\mem_wdata_r2[2]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[0]~q ),
	.ena(vcc),
	.q(wdp_wdata_h_2x_2),
	.prn(vcc));
defparam \wdp_wdata_h_2x[2] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[2] .power_up = "low";

dffeas \wdp_wdata_l_2x[3] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[99]~q ),
	.asdata(\mem_wdata_r2[35]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[0]~q ),
	.ena(vcc),
	.q(wdp_wdata_l_2x_3),
	.prn(vcc));
defparam \wdp_wdata_l_2x[3] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[3] .power_up = "low";

dffeas \wdp_wdata_h_2x[3] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[67]~q ),
	.asdata(\mem_wdata_r2[3]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[0]~q ),
	.ena(vcc),
	.q(wdp_wdata_h_2x_3),
	.prn(vcc));
defparam \wdp_wdata_h_2x[3] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[3] .power_up = "low";

dffeas \wdp_wdata_l_2x[4] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[100]~q ),
	.asdata(\mem_wdata_r2[36]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[1]~q ),
	.ena(vcc),
	.q(wdp_wdata_l_2x_4),
	.prn(vcc));
defparam \wdp_wdata_l_2x[4] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[4] .power_up = "low";

dffeas \wdp_wdata_h_2x[4] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[68]~q ),
	.asdata(\mem_wdata_r2[4]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[1]~q ),
	.ena(vcc),
	.q(wdp_wdata_h_2x_4),
	.prn(vcc));
defparam \wdp_wdata_h_2x[4] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[4] .power_up = "low";

dffeas \dq_oe_2x[1] (
	.clk(write_clk_2x),
	.d(\wdata_valid_1x_r2[9]~q ),
	.asdata(\wdata_valid_1x_r2[1]~q ),
	.clrn(reset_write_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[1]~q ),
	.ena(vcc),
	.q(dq_oe_2x_1),
	.prn(vcc));
defparam \dq_oe_2x[1] .is_wysiwyg = "true";
defparam \dq_oe_2x[1] .power_up = "low";

dffeas \wdp_wdata_l_2x[5] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[101]~q ),
	.asdata(\mem_wdata_r2[37]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[1]~q ),
	.ena(vcc),
	.q(wdp_wdata_l_2x_5),
	.prn(vcc));
defparam \wdp_wdata_l_2x[5] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[5] .power_up = "low";

dffeas \wdp_wdata_h_2x[5] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[69]~q ),
	.asdata(\mem_wdata_r2[5]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[1]~q ),
	.ena(vcc),
	.q(wdp_wdata_h_2x_5),
	.prn(vcc));
defparam \wdp_wdata_h_2x[5] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[5] .power_up = "low";

dffeas \wdp_wdata_l_2x[6] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[102]~q ),
	.asdata(\mem_wdata_r2[38]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[1]~q ),
	.ena(vcc),
	.q(wdp_wdata_l_2x_6),
	.prn(vcc));
defparam \wdp_wdata_l_2x[6] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[6] .power_up = "low";

dffeas \wdp_wdata_h_2x[6] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[70]~q ),
	.asdata(\mem_wdata_r2[6]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[1]~q ),
	.ena(vcc),
	.q(wdp_wdata_h_2x_6),
	.prn(vcc));
defparam \wdp_wdata_h_2x[6] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[6] .power_up = "low";

dffeas \wdp_wdata_l_2x[7] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[103]~q ),
	.asdata(\mem_wdata_r2[39]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[1]~q ),
	.ena(vcc),
	.q(wdp_wdata_l_2x_7),
	.prn(vcc));
defparam \wdp_wdata_l_2x[7] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[7] .power_up = "low";

dffeas \wdp_wdata_h_2x[7] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[71]~q ),
	.asdata(\mem_wdata_r2[7]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[1]~q ),
	.ena(vcc),
	.q(wdp_wdata_h_2x_7),
	.prn(vcc));
defparam \wdp_wdata_h_2x[7] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[7] .power_up = "low";

dffeas \wdp_wdata_l_2x[8] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[104]~q ),
	.asdata(\mem_wdata_r2[40]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[2]~q ),
	.ena(vcc),
	.q(wdp_wdata_l_2x_8),
	.prn(vcc));
defparam \wdp_wdata_l_2x[8] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[8] .power_up = "low";

dffeas \wdp_wdata_h_2x[8] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[72]~q ),
	.asdata(\mem_wdata_r2[8]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[2]~q ),
	.ena(vcc),
	.q(wdp_wdata_h_2x_8),
	.prn(vcc));
defparam \wdp_wdata_h_2x[8] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[8] .power_up = "low";

dffeas \dq_oe_2x[2] (
	.clk(write_clk_2x),
	.d(\wdata_valid_1x_r2[10]~q ),
	.asdata(\wdata_valid_1x_r2[2]~q ),
	.clrn(reset_write_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[2]~q ),
	.ena(vcc),
	.q(dq_oe_2x_2),
	.prn(vcc));
defparam \dq_oe_2x[2] .is_wysiwyg = "true";
defparam \dq_oe_2x[2] .power_up = "low";

dffeas \wdp_wdata_l_2x[9] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[105]~q ),
	.asdata(\mem_wdata_r2[41]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[2]~q ),
	.ena(vcc),
	.q(wdp_wdata_l_2x_9),
	.prn(vcc));
defparam \wdp_wdata_l_2x[9] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[9] .power_up = "low";

dffeas \wdp_wdata_h_2x[9] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[73]~q ),
	.asdata(\mem_wdata_r2[9]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[2]~q ),
	.ena(vcc),
	.q(wdp_wdata_h_2x_9),
	.prn(vcc));
defparam \wdp_wdata_h_2x[9] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[9] .power_up = "low";

dffeas \wdp_wdata_l_2x[10] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[106]~q ),
	.asdata(\mem_wdata_r2[42]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[2]~q ),
	.ena(vcc),
	.q(wdp_wdata_l_2x_10),
	.prn(vcc));
defparam \wdp_wdata_l_2x[10] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[10] .power_up = "low";

dffeas \wdp_wdata_h_2x[10] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[74]~q ),
	.asdata(\mem_wdata_r2[10]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[2]~q ),
	.ena(vcc),
	.q(wdp_wdata_h_2x_10),
	.prn(vcc));
defparam \wdp_wdata_h_2x[10] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[10] .power_up = "low";

dffeas \wdp_wdata_l_2x[11] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[107]~q ),
	.asdata(\mem_wdata_r2[43]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[2]~q ),
	.ena(vcc),
	.q(wdp_wdata_l_2x_11),
	.prn(vcc));
defparam \wdp_wdata_l_2x[11] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[11] .power_up = "low";

dffeas \wdp_wdata_h_2x[11] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[75]~q ),
	.asdata(\mem_wdata_r2[11]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[2]~q ),
	.ena(vcc),
	.q(wdp_wdata_h_2x_11),
	.prn(vcc));
defparam \wdp_wdata_h_2x[11] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[11] .power_up = "low";

dffeas \wdp_wdata_l_2x[12] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[108]~q ),
	.asdata(\mem_wdata_r2[44]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[3]~q ),
	.ena(vcc),
	.q(wdp_wdata_l_2x_12),
	.prn(vcc));
defparam \wdp_wdata_l_2x[12] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[12] .power_up = "low";

dffeas \wdp_wdata_h_2x[12] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[76]~q ),
	.asdata(\mem_wdata_r2[12]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[3]~q ),
	.ena(vcc),
	.q(wdp_wdata_h_2x_12),
	.prn(vcc));
defparam \wdp_wdata_h_2x[12] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[12] .power_up = "low";

dffeas \dq_oe_2x[3] (
	.clk(write_clk_2x),
	.d(\wdata_valid_1x_r2[11]~q ),
	.asdata(\wdata_valid_1x_r2[3]~q ),
	.clrn(reset_write_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[3]~q ),
	.ena(vcc),
	.q(dq_oe_2x_3),
	.prn(vcc));
defparam \dq_oe_2x[3] .is_wysiwyg = "true";
defparam \dq_oe_2x[3] .power_up = "low";

dffeas \wdp_wdata_l_2x[13] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[109]~q ),
	.asdata(\mem_wdata_r2[45]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[3]~q ),
	.ena(vcc),
	.q(wdp_wdata_l_2x_13),
	.prn(vcc));
defparam \wdp_wdata_l_2x[13] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[13] .power_up = "low";

dffeas \wdp_wdata_h_2x[13] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[77]~q ),
	.asdata(\mem_wdata_r2[13]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[3]~q ),
	.ena(vcc),
	.q(wdp_wdata_h_2x_13),
	.prn(vcc));
defparam \wdp_wdata_h_2x[13] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[13] .power_up = "low";

dffeas \wdp_wdata_l_2x[14] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[110]~q ),
	.asdata(\mem_wdata_r2[46]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[3]~q ),
	.ena(vcc),
	.q(wdp_wdata_l_2x_14),
	.prn(vcc));
defparam \wdp_wdata_l_2x[14] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[14] .power_up = "low";

dffeas \wdp_wdata_h_2x[14] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[78]~q ),
	.asdata(\mem_wdata_r2[14]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[3]~q ),
	.ena(vcc),
	.q(wdp_wdata_h_2x_14),
	.prn(vcc));
defparam \wdp_wdata_h_2x[14] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[14] .power_up = "low";

dffeas \wdp_wdata_l_2x[15] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[111]~q ),
	.asdata(\mem_wdata_r2[47]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[3]~q ),
	.ena(vcc),
	.q(wdp_wdata_l_2x_15),
	.prn(vcc));
defparam \wdp_wdata_l_2x[15] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[15] .power_up = "low";

dffeas \wdp_wdata_h_2x[15] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[79]~q ),
	.asdata(\mem_wdata_r2[15]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[3]~q ),
	.ena(vcc),
	.q(wdp_wdata_h_2x_15),
	.prn(vcc));
defparam \wdp_wdata_h_2x[15] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[15] .power_up = "low";

dffeas \wdp_wdata_l_2x[16] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[112]~q ),
	.asdata(\mem_wdata_r2[48]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[4]~q ),
	.ena(vcc),
	.q(wdp_wdata_l_2x_16),
	.prn(vcc));
defparam \wdp_wdata_l_2x[16] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[16] .power_up = "low";

dffeas \wdp_wdata_h_2x[16] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[80]~q ),
	.asdata(\mem_wdata_r2[16]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[4]~q ),
	.ena(vcc),
	.q(wdp_wdata_h_2x_16),
	.prn(vcc));
defparam \wdp_wdata_h_2x[16] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[16] .power_up = "low";

dffeas \dq_oe_2x[4] (
	.clk(write_clk_2x),
	.d(\wdata_valid_1x_r2[12]~q ),
	.asdata(\wdata_valid_1x_r2[4]~q ),
	.clrn(reset_write_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[4]~q ),
	.ena(vcc),
	.q(dq_oe_2x_4),
	.prn(vcc));
defparam \dq_oe_2x[4] .is_wysiwyg = "true";
defparam \dq_oe_2x[4] .power_up = "low";

dffeas \wdp_wdata_l_2x[17] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[113]~q ),
	.asdata(\mem_wdata_r2[49]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[4]~q ),
	.ena(vcc),
	.q(wdp_wdata_l_2x_17),
	.prn(vcc));
defparam \wdp_wdata_l_2x[17] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[17] .power_up = "low";

dffeas \wdp_wdata_h_2x[17] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[81]~q ),
	.asdata(\mem_wdata_r2[17]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[4]~q ),
	.ena(vcc),
	.q(wdp_wdata_h_2x_17),
	.prn(vcc));
defparam \wdp_wdata_h_2x[17] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[17] .power_up = "low";

dffeas \wdp_wdata_l_2x[18] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[114]~q ),
	.asdata(\mem_wdata_r2[50]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[4]~q ),
	.ena(vcc),
	.q(wdp_wdata_l_2x_18),
	.prn(vcc));
defparam \wdp_wdata_l_2x[18] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[18] .power_up = "low";

dffeas \wdp_wdata_h_2x[18] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[82]~q ),
	.asdata(\mem_wdata_r2[18]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[4]~q ),
	.ena(vcc),
	.q(wdp_wdata_h_2x_18),
	.prn(vcc));
defparam \wdp_wdata_h_2x[18] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[18] .power_up = "low";

dffeas \wdp_wdata_l_2x[19] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[115]~q ),
	.asdata(\mem_wdata_r2[51]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[4]~q ),
	.ena(vcc),
	.q(wdp_wdata_l_2x_19),
	.prn(vcc));
defparam \wdp_wdata_l_2x[19] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[19] .power_up = "low";

dffeas \wdp_wdata_h_2x[19] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[83]~q ),
	.asdata(\mem_wdata_r2[19]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[4]~q ),
	.ena(vcc),
	.q(wdp_wdata_h_2x_19),
	.prn(vcc));
defparam \wdp_wdata_h_2x[19] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[19] .power_up = "low";

dffeas \wdp_wdata_l_2x[20] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[116]~q ),
	.asdata(\mem_wdata_r2[52]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[5]~q ),
	.ena(vcc),
	.q(wdp_wdata_l_2x_20),
	.prn(vcc));
defparam \wdp_wdata_l_2x[20] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[20] .power_up = "low";

dffeas \wdp_wdata_h_2x[20] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[84]~q ),
	.asdata(\mem_wdata_r2[20]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[5]~q ),
	.ena(vcc),
	.q(wdp_wdata_h_2x_20),
	.prn(vcc));
defparam \wdp_wdata_h_2x[20] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[20] .power_up = "low";

dffeas \dq_oe_2x[5] (
	.clk(write_clk_2x),
	.d(\wdata_valid_1x_r2[13]~q ),
	.asdata(\wdata_valid_1x_r2[5]~q ),
	.clrn(reset_write_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[5]~q ),
	.ena(vcc),
	.q(dq_oe_2x_5),
	.prn(vcc));
defparam \dq_oe_2x[5] .is_wysiwyg = "true";
defparam \dq_oe_2x[5] .power_up = "low";

dffeas \wdp_wdata_l_2x[21] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[117]~q ),
	.asdata(\mem_wdata_r2[53]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[5]~q ),
	.ena(vcc),
	.q(wdp_wdata_l_2x_21),
	.prn(vcc));
defparam \wdp_wdata_l_2x[21] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[21] .power_up = "low";

dffeas \wdp_wdata_h_2x[21] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[85]~q ),
	.asdata(\mem_wdata_r2[21]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[5]~q ),
	.ena(vcc),
	.q(wdp_wdata_h_2x_21),
	.prn(vcc));
defparam \wdp_wdata_h_2x[21] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[21] .power_up = "low";

dffeas \wdp_wdata_l_2x[22] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[118]~q ),
	.asdata(\mem_wdata_r2[54]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[5]~q ),
	.ena(vcc),
	.q(wdp_wdata_l_2x_22),
	.prn(vcc));
defparam \wdp_wdata_l_2x[22] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[22] .power_up = "low";

dffeas \wdp_wdata_h_2x[22] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[86]~q ),
	.asdata(\mem_wdata_r2[22]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[5]~q ),
	.ena(vcc),
	.q(wdp_wdata_h_2x_22),
	.prn(vcc));
defparam \wdp_wdata_h_2x[22] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[22] .power_up = "low";

dffeas \wdp_wdata_l_2x[23] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[119]~q ),
	.asdata(\mem_wdata_r2[55]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[5]~q ),
	.ena(vcc),
	.q(wdp_wdata_l_2x_23),
	.prn(vcc));
defparam \wdp_wdata_l_2x[23] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[23] .power_up = "low";

dffeas \wdp_wdata_h_2x[23] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[87]~q ),
	.asdata(\mem_wdata_r2[23]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[5]~q ),
	.ena(vcc),
	.q(wdp_wdata_h_2x_23),
	.prn(vcc));
defparam \wdp_wdata_h_2x[23] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[23] .power_up = "low";

dffeas \wdp_wdata_l_2x[24] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[120]~q ),
	.asdata(\mem_wdata_r2[56]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[6]~q ),
	.ena(vcc),
	.q(wdp_wdata_l_2x_24),
	.prn(vcc));
defparam \wdp_wdata_l_2x[24] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[24] .power_up = "low";

dffeas \wdp_wdata_h_2x[24] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[88]~q ),
	.asdata(\mem_wdata_r2[24]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[6]~q ),
	.ena(vcc),
	.q(wdp_wdata_h_2x_24),
	.prn(vcc));
defparam \wdp_wdata_h_2x[24] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[24] .power_up = "low";

dffeas \dq_oe_2x[6] (
	.clk(write_clk_2x),
	.d(\wdata_valid_1x_r2[14]~q ),
	.asdata(\wdata_valid_1x_r2[6]~q ),
	.clrn(reset_write_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[6]~q ),
	.ena(vcc),
	.q(dq_oe_2x_6),
	.prn(vcc));
defparam \dq_oe_2x[6] .is_wysiwyg = "true";
defparam \dq_oe_2x[6] .power_up = "low";

dffeas \wdp_wdata_l_2x[25] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[121]~q ),
	.asdata(\mem_wdata_r2[57]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[6]~q ),
	.ena(vcc),
	.q(wdp_wdata_l_2x_25),
	.prn(vcc));
defparam \wdp_wdata_l_2x[25] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[25] .power_up = "low";

dffeas \wdp_wdata_h_2x[25] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[89]~q ),
	.asdata(\mem_wdata_r2[25]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[6]~q ),
	.ena(vcc),
	.q(wdp_wdata_h_2x_25),
	.prn(vcc));
defparam \wdp_wdata_h_2x[25] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[25] .power_up = "low";

dffeas \wdp_wdata_l_2x[26] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[122]~q ),
	.asdata(\mem_wdata_r2[58]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[6]~q ),
	.ena(vcc),
	.q(wdp_wdata_l_2x_26),
	.prn(vcc));
defparam \wdp_wdata_l_2x[26] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[26] .power_up = "low";

dffeas \wdp_wdata_h_2x[26] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[90]~q ),
	.asdata(\mem_wdata_r2[26]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[6]~q ),
	.ena(vcc),
	.q(wdp_wdata_h_2x_26),
	.prn(vcc));
defparam \wdp_wdata_h_2x[26] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[26] .power_up = "low";

dffeas \wdp_wdata_l_2x[27] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[123]~q ),
	.asdata(\mem_wdata_r2[59]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[6]~q ),
	.ena(vcc),
	.q(wdp_wdata_l_2x_27),
	.prn(vcc));
defparam \wdp_wdata_l_2x[27] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[27] .power_up = "low";

dffeas \wdp_wdata_h_2x[27] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[91]~q ),
	.asdata(\mem_wdata_r2[27]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[6]~q ),
	.ena(vcc),
	.q(wdp_wdata_h_2x_27),
	.prn(vcc));
defparam \wdp_wdata_h_2x[27] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[27] .power_up = "low";

dffeas \wdp_wdata_l_2x[28] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[124]~q ),
	.asdata(\mem_wdata_r2[60]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[7]~q ),
	.ena(vcc),
	.q(wdp_wdata_l_2x_28),
	.prn(vcc));
defparam \wdp_wdata_l_2x[28] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[28] .power_up = "low";

dffeas \wdp_wdata_h_2x[28] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[92]~q ),
	.asdata(\mem_wdata_r2[28]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[7]~q ),
	.ena(vcc),
	.q(wdp_wdata_h_2x_28),
	.prn(vcc));
defparam \wdp_wdata_h_2x[28] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[28] .power_up = "low";

dffeas \dq_oe_2x[7] (
	.clk(write_clk_2x),
	.d(\wdata_valid_1x_r2[15]~q ),
	.asdata(\wdata_valid_1x_r2[7]~q ),
	.clrn(reset_write_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[7]~q ),
	.ena(vcc),
	.q(dq_oe_2x_7),
	.prn(vcc));
defparam \dq_oe_2x[7] .is_wysiwyg = "true";
defparam \dq_oe_2x[7] .power_up = "low";

dffeas \wdp_wdata_l_2x[29] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[125]~q ),
	.asdata(\mem_wdata_r2[61]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[7]~q ),
	.ena(vcc),
	.q(wdp_wdata_l_2x_29),
	.prn(vcc));
defparam \wdp_wdata_l_2x[29] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[29] .power_up = "low";

dffeas \wdp_wdata_h_2x[29] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[93]~q ),
	.asdata(\mem_wdata_r2[29]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[7]~q ),
	.ena(vcc),
	.q(wdp_wdata_h_2x_29),
	.prn(vcc));
defparam \wdp_wdata_h_2x[29] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[29] .power_up = "low";

dffeas \wdp_wdata_l_2x[30] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[126]~q ),
	.asdata(\mem_wdata_r2[62]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[7]~q ),
	.ena(vcc),
	.q(wdp_wdata_l_2x_30),
	.prn(vcc));
defparam \wdp_wdata_l_2x[30] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[30] .power_up = "low";

dffeas \wdp_wdata_h_2x[30] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[94]~q ),
	.asdata(\mem_wdata_r2[30]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[7]~q ),
	.ena(vcc),
	.q(wdp_wdata_h_2x_30),
	.prn(vcc));
defparam \wdp_wdata_h_2x[30] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[30] .power_up = "low";

dffeas \wdp_wdata_l_2x[31] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[127]~q ),
	.asdata(\mem_wdata_r2[63]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[7]~q ),
	.ena(vcc),
	.q(wdp_wdata_l_2x_31),
	.prn(vcc));
defparam \wdp_wdata_l_2x[31] .is_wysiwyg = "true";
defparam \wdp_wdata_l_2x[31] .power_up = "low";

dffeas \wdp_wdata_h_2x[31] (
	.clk(write_clk_2x),
	.d(\mem_wdata_r2[95]~q ),
	.asdata(\mem_wdata_r2[31]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\wdata_sel[7]~q ),
	.ena(vcc),
	.q(wdp_wdata_h_2x_31),
	.prn(vcc));
defparam \wdp_wdata_h_2x[31] .is_wysiwyg = "true";
defparam \wdp_wdata_h_2x[31] .power_up = "low";

dffeas \dqs_burst_2x_r3[0] (
	.clk(mem_clk_2x),
	.d(\dqs_burst_2x_r2[0]~q ),
	.asdata(vcc),
	.clrn(reset_mem_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dqs_burst_2x_r3_0),
	.prn(vcc));
defparam \dqs_burst_2x_r3[0] .is_wysiwyg = "true";
defparam \dqs_burst_2x_r3[0] .power_up = "low";

dffeas \dqs_burst_2x_r3[1] (
	.clk(mem_clk_2x),
	.d(\dqs_burst_2x_r2[1]~q ),
	.asdata(vcc),
	.clrn(reset_mem_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dqs_burst_2x_r3_1),
	.prn(vcc));
defparam \dqs_burst_2x_r3[1] .is_wysiwyg = "true";
defparam \dqs_burst_2x_r3[1] .power_up = "low";

dffeas \dqs_burst_2x_r3[2] (
	.clk(mem_clk_2x),
	.d(\dqs_burst_2x_r2[2]~q ),
	.asdata(vcc),
	.clrn(reset_mem_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dqs_burst_2x_r3_2),
	.prn(vcc));
defparam \dqs_burst_2x_r3[2] .is_wysiwyg = "true";
defparam \dqs_burst_2x_r3[2] .power_up = "low";

dffeas \dqs_burst_2x_r3[3] (
	.clk(mem_clk_2x),
	.d(\dqs_burst_2x_r2[3]~q ),
	.asdata(vcc),
	.clrn(reset_mem_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dqs_burst_2x_r3_3),
	.prn(vcc));
defparam \dqs_burst_2x_r3[3] .is_wysiwyg = "true";
defparam \dqs_burst_2x_r3[3] .power_up = "low";

dffeas \mem_dm_r1[4] (
	.clk(phy_clk_1x),
	.d(afi_dm_4),
	.asdata(dgwb_wdp_ovride1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_wdp_ovride),
	.ena(vcc),
	.q(\mem_dm_r1[4]~q ),
	.prn(vcc));
defparam \mem_dm_r1[4] .is_wysiwyg = "true";
defparam \mem_dm_r1[4] .power_up = "low";

dffeas \mem_dm_r2[4] (
	.clk(phy_clk_1x),
	.d(\mem_dm_r1[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_dm_r2[4]~q ),
	.prn(vcc));
defparam \mem_dm_r2[4] .is_wysiwyg = "true";
defparam \mem_dm_r2[4] .power_up = "low";

dffeas \mem_dm_r1[12] (
	.clk(phy_clk_1x),
	.d(afi_dm_12),
	.asdata(dgwb_wdp_ovride1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_wdp_ovride),
	.ena(vcc),
	.q(\mem_dm_r1[12]~q ),
	.prn(vcc));
defparam \mem_dm_r1[12] .is_wysiwyg = "true";
defparam \mem_dm_r1[12] .power_up = "low";

dffeas \mem_dm_r2[12] (
	.clk(phy_clk_1x),
	.d(\mem_dm_r1[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_dm_r2[12]~q ),
	.prn(vcc));
defparam \mem_dm_r2[12] .is_wysiwyg = "true";
defparam \mem_dm_r2[12] .power_up = "low";

arriaii_lcell_comb \mem_wdata_valid[0]~0 (
	.dataa(!ctl_init_fail),
	.datab(!ctl_init_success),
	.datac(!dgwb_wdp_ovride),
	.datad(!int_wdata_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata_valid[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata_valid[0]~0 .extended_lut = "off";
defparam \mem_wdata_valid[0]~0 .lut_mask = 64'h08FF08FF08FF08FF;
defparam \mem_wdata_valid[0]~0 .shared_arith = "off";

dffeas wdata_dm_1x_r(
	.clk(phy_clk_1x),
	.d(\mem_wdata_valid[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_dm_1x_r~q ),
	.prn(vcc));
defparam wdata_dm_1x_r.is_wysiwyg = "true";
defparam wdata_dm_1x_r.power_up = "low";

dffeas wdata_dm_2x_r1(
	.clk(write_clk_2x),
	.d(\wdata_dm_1x_r~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_dm_2x_r1~q ),
	.prn(vcc));
defparam wdata_dm_2x_r1.is_wysiwyg = "true";
defparam wdata_dm_2x_r1.power_up = "low";

dffeas wdata_dm_2x_r2(
	.clk(write_clk_2x),
	.d(\wdata_dm_2x_r1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_dm_2x_r2~q ),
	.prn(vcc));
defparam wdata_dm_2x_r2.is_wysiwyg = "true";
defparam wdata_dm_2x_r2.power_up = "low";

arriaii_lcell_comb \dm_sel~0 (
	.dataa(!\dm_sel~q ),
	.datab(!\wdata_dm_2x_r1~q ),
	.datac(!\wdata_dm_2x_r2~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dm_sel~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dm_sel~0 .extended_lut = "off";
defparam \dm_sel~0 .lut_mask = 64'h8A8A8A8A8A8A8A8A;
defparam \dm_sel~0 .shared_arith = "off";

dffeas dm_sel(
	.clk(write_clk_2x),
	.d(\dm_sel~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dm_sel~q ),
	.prn(vcc));
defparam dm_sel.is_wysiwyg = "true";
defparam dm_sel.power_up = "low";

dffeas \mem_dm_r1[0] (
	.clk(phy_clk_1x),
	.d(afi_dm_0),
	.asdata(dgwb_wdp_ovride1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_wdp_ovride),
	.ena(vcc),
	.q(\mem_dm_r1[0]~q ),
	.prn(vcc));
defparam \mem_dm_r1[0] .is_wysiwyg = "true";
defparam \mem_dm_r1[0] .power_up = "low";

dffeas \mem_dm_r2[0] (
	.clk(phy_clk_1x),
	.d(\mem_dm_r1[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_dm_r2[0]~q ),
	.prn(vcc));
defparam \mem_dm_r2[0] .is_wysiwyg = "true";
defparam \mem_dm_r2[0] .power_up = "low";

dffeas \mem_dm_r1[8] (
	.clk(phy_clk_1x),
	.d(afi_dm_8),
	.asdata(dgwb_wdp_ovride1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_wdp_ovride),
	.ena(vcc),
	.q(\mem_dm_r1[8]~q ),
	.prn(vcc));
defparam \mem_dm_r1[8] .is_wysiwyg = "true";
defparam \mem_dm_r1[8] .power_up = "low";

dffeas \mem_dm_r2[8] (
	.clk(phy_clk_1x),
	.d(\mem_dm_r1[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_dm_r2[8]~q ),
	.prn(vcc));
defparam \mem_dm_r2[8] .is_wysiwyg = "true";
defparam \mem_dm_r2[8] .power_up = "low";

dffeas \mem_dm_r1[5] (
	.clk(phy_clk_1x),
	.d(afi_dm_5),
	.asdata(dgwb_wdp_ovride1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_wdp_ovride),
	.ena(vcc),
	.q(\mem_dm_r1[5]~q ),
	.prn(vcc));
defparam \mem_dm_r1[5] .is_wysiwyg = "true";
defparam \mem_dm_r1[5] .power_up = "low";

dffeas \mem_dm_r2[5] (
	.clk(phy_clk_1x),
	.d(\mem_dm_r1[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_dm_r2[5]~q ),
	.prn(vcc));
defparam \mem_dm_r2[5] .is_wysiwyg = "true";
defparam \mem_dm_r2[5] .power_up = "low";

dffeas \mem_dm_r1[13] (
	.clk(phy_clk_1x),
	.d(afi_dm_13),
	.asdata(dgwb_wdp_ovride1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_wdp_ovride),
	.ena(vcc),
	.q(\mem_dm_r1[13]~q ),
	.prn(vcc));
defparam \mem_dm_r1[13] .is_wysiwyg = "true";
defparam \mem_dm_r1[13] .power_up = "low";

dffeas \mem_dm_r2[13] (
	.clk(phy_clk_1x),
	.d(\mem_dm_r1[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_dm_r2[13]~q ),
	.prn(vcc));
defparam \mem_dm_r2[13] .is_wysiwyg = "true";
defparam \mem_dm_r2[13] .power_up = "low";

dffeas \mem_dm_r1[1] (
	.clk(phy_clk_1x),
	.d(afi_dm_1),
	.asdata(dgwb_wdp_ovride1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_wdp_ovride),
	.ena(vcc),
	.q(\mem_dm_r1[1]~q ),
	.prn(vcc));
defparam \mem_dm_r1[1] .is_wysiwyg = "true";
defparam \mem_dm_r1[1] .power_up = "low";

dffeas \mem_dm_r2[1] (
	.clk(phy_clk_1x),
	.d(\mem_dm_r1[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_dm_r2[1]~q ),
	.prn(vcc));
defparam \mem_dm_r2[1] .is_wysiwyg = "true";
defparam \mem_dm_r2[1] .power_up = "low";

dffeas \mem_dm_r1[9] (
	.clk(phy_clk_1x),
	.d(afi_dm_9),
	.asdata(dgwb_wdp_ovride1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_wdp_ovride),
	.ena(vcc),
	.q(\mem_dm_r1[9]~q ),
	.prn(vcc));
defparam \mem_dm_r1[9] .is_wysiwyg = "true";
defparam \mem_dm_r1[9] .power_up = "low";

dffeas \mem_dm_r2[9] (
	.clk(phy_clk_1x),
	.d(\mem_dm_r1[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_dm_r2[9]~q ),
	.prn(vcc));
defparam \mem_dm_r2[9] .is_wysiwyg = "true";
defparam \mem_dm_r2[9] .power_up = "low";

dffeas \mem_dm_r1[6] (
	.clk(phy_clk_1x),
	.d(afi_dm_6),
	.asdata(dgwb_wdp_ovride1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_wdp_ovride),
	.ena(vcc),
	.q(\mem_dm_r1[6]~q ),
	.prn(vcc));
defparam \mem_dm_r1[6] .is_wysiwyg = "true";
defparam \mem_dm_r1[6] .power_up = "low";

dffeas \mem_dm_r2[6] (
	.clk(phy_clk_1x),
	.d(\mem_dm_r1[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_dm_r2[6]~q ),
	.prn(vcc));
defparam \mem_dm_r2[6] .is_wysiwyg = "true";
defparam \mem_dm_r2[6] .power_up = "low";

dffeas \mem_dm_r1[14] (
	.clk(phy_clk_1x),
	.d(afi_dm_14),
	.asdata(dgwb_wdp_ovride1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_wdp_ovride),
	.ena(vcc),
	.q(\mem_dm_r1[14]~q ),
	.prn(vcc));
defparam \mem_dm_r1[14] .is_wysiwyg = "true";
defparam \mem_dm_r1[14] .power_up = "low";

dffeas \mem_dm_r2[14] (
	.clk(phy_clk_1x),
	.d(\mem_dm_r1[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_dm_r2[14]~q ),
	.prn(vcc));
defparam \mem_dm_r2[14] .is_wysiwyg = "true";
defparam \mem_dm_r2[14] .power_up = "low";

dffeas \mem_dm_r1[2] (
	.clk(phy_clk_1x),
	.d(afi_dm_2),
	.asdata(dgwb_wdp_ovride1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_wdp_ovride),
	.ena(vcc),
	.q(\mem_dm_r1[2]~q ),
	.prn(vcc));
defparam \mem_dm_r1[2] .is_wysiwyg = "true";
defparam \mem_dm_r1[2] .power_up = "low";

dffeas \mem_dm_r2[2] (
	.clk(phy_clk_1x),
	.d(\mem_dm_r1[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_dm_r2[2]~q ),
	.prn(vcc));
defparam \mem_dm_r2[2] .is_wysiwyg = "true";
defparam \mem_dm_r2[2] .power_up = "low";

dffeas \mem_dm_r1[10] (
	.clk(phy_clk_1x),
	.d(afi_dm_10),
	.asdata(dgwb_wdp_ovride1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_wdp_ovride),
	.ena(vcc),
	.q(\mem_dm_r1[10]~q ),
	.prn(vcc));
defparam \mem_dm_r1[10] .is_wysiwyg = "true";
defparam \mem_dm_r1[10] .power_up = "low";

dffeas \mem_dm_r2[10] (
	.clk(phy_clk_1x),
	.d(\mem_dm_r1[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_dm_r2[10]~q ),
	.prn(vcc));
defparam \mem_dm_r2[10] .is_wysiwyg = "true";
defparam \mem_dm_r2[10] .power_up = "low";

dffeas \mem_dm_r1[7] (
	.clk(phy_clk_1x),
	.d(afi_dm_7),
	.asdata(dgwb_wdp_ovride1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_wdp_ovride),
	.ena(vcc),
	.q(\mem_dm_r1[7]~q ),
	.prn(vcc));
defparam \mem_dm_r1[7] .is_wysiwyg = "true";
defparam \mem_dm_r1[7] .power_up = "low";

dffeas \mem_dm_r2[7] (
	.clk(phy_clk_1x),
	.d(\mem_dm_r1[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_dm_r2[7]~q ),
	.prn(vcc));
defparam \mem_dm_r2[7] .is_wysiwyg = "true";
defparam \mem_dm_r2[7] .power_up = "low";

dffeas \mem_dm_r1[15] (
	.clk(phy_clk_1x),
	.d(afi_dm_15),
	.asdata(dgwb_wdp_ovride1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_wdp_ovride),
	.ena(vcc),
	.q(\mem_dm_r1[15]~q ),
	.prn(vcc));
defparam \mem_dm_r1[15] .is_wysiwyg = "true";
defparam \mem_dm_r1[15] .power_up = "low";

dffeas \mem_dm_r2[15] (
	.clk(phy_clk_1x),
	.d(\mem_dm_r1[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_dm_r2[15]~q ),
	.prn(vcc));
defparam \mem_dm_r2[15] .is_wysiwyg = "true";
defparam \mem_dm_r2[15] .power_up = "low";

dffeas \mem_dm_r1[3] (
	.clk(phy_clk_1x),
	.d(afi_dm_3),
	.asdata(dgwb_wdp_ovride1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_wdp_ovride),
	.ena(vcc),
	.q(\mem_dm_r1[3]~q ),
	.prn(vcc));
defparam \mem_dm_r1[3] .is_wysiwyg = "true";
defparam \mem_dm_r1[3] .power_up = "low";

dffeas \mem_dm_r2[3] (
	.clk(phy_clk_1x),
	.d(\mem_dm_r1[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_dm_r2[3]~q ),
	.prn(vcc));
defparam \mem_dm_r2[3] .is_wysiwyg = "true";
defparam \mem_dm_r2[3] .power_up = "low";

dffeas \mem_dm_r1[11] (
	.clk(phy_clk_1x),
	.d(afi_dm_11),
	.asdata(dgwb_wdp_ovride1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(seq_wdp_ovride),
	.ena(vcc),
	.q(\mem_dm_r1[11]~q ),
	.prn(vcc));
defparam \mem_dm_r1[11] .is_wysiwyg = "true";
defparam \mem_dm_r1[11] .power_up = "low";

dffeas \mem_dm_r2[11] (
	.clk(phy_clk_1x),
	.d(\mem_dm_r1[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_dm_r2[11]~q ),
	.prn(vcc));
defparam \mem_dm_r2[11] .is_wysiwyg = "true";
defparam \mem_dm_r2[11] .power_up = "low";

arriaii_lcell_comb \mem_wdata[96]~0 (
	.dataa(!seq_wdp_ovride),
	.datab(!q_b_96),
	.datac(!dgwb_wdata_120),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[96]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[96]~0 .extended_lut = "off";
defparam \mem_wdata[96]~0 .lut_mask = 64'h2727272727272727;
defparam \mem_wdata[96]~0 .shared_arith = "off";

dffeas \mem_wdata_r1[96] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[96]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[96]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[96] .is_wysiwyg = "true";
defparam \mem_wdata_r1[96] .power_up = "low";

dffeas \mem_wdata_r2[96] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[96]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[96]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[96] .is_wysiwyg = "true";
defparam \mem_wdata_r2[96] .power_up = "low";

arriaii_lcell_comb \mem_wdata[32]~1 (
	.dataa(!seq_wdp_ovride),
	.datab(!q_b_32),
	.datac(!dgwb_wdata_56),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[32]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[32]~1 .extended_lut = "off";
defparam \mem_wdata[32]~1 .lut_mask = 64'h2727272727272727;
defparam \mem_wdata[32]~1 .shared_arith = "off";

dffeas \mem_wdata_r1[32] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[32]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[32]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[32] .is_wysiwyg = "true";
defparam \mem_wdata_r1[32] .power_up = "low";

dffeas \mem_wdata_r2[32] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[32]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[32]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[32] .is_wysiwyg = "true";
defparam \mem_wdata_r2[32] .power_up = "low";

dffeas \wdata_valid_1x_r[0] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_valid[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r[0]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r[0] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r[0] .power_up = "low";

dffeas \wdata_valid_2x_r1[0] (
	.clk(write_clk_2x),
	.d(\wdata_valid_1x_r[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_2x_r1[0]~q ),
	.prn(vcc));
defparam \wdata_valid_2x_r1[0] .is_wysiwyg = "true";
defparam \wdata_valid_2x_r1[0] .power_up = "low";

dffeas \wdata_valid_2x_r2[0] (
	.clk(write_clk_2x),
	.d(\wdata_valid_2x_r1[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_2x_r2[0]~q ),
	.prn(vcc));
defparam \wdata_valid_2x_r2[0] .is_wysiwyg = "true";
defparam \wdata_valid_2x_r2[0] .power_up = "low";

arriaii_lcell_comb \wdata_sel~0 (
	.dataa(!\wdata_sel[0]~q ),
	.datab(!\wdata_valid_2x_r2[0]~q ),
	.datac(!\wdata_valid_2x_r1[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wdata_sel~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wdata_sel~0 .extended_lut = "off";
defparam \wdata_sel~0 .lut_mask = 64'hA2A2A2A2A2A2A2A2;
defparam \wdata_sel~0 .shared_arith = "off";

dffeas \wdata_sel[0] (
	.clk(write_clk_2x),
	.d(\wdata_sel~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_sel[0]~q ),
	.prn(vcc));
defparam \wdata_sel[0] .is_wysiwyg = "true";
defparam \wdata_sel[0] .power_up = "low";

arriaii_lcell_comb \mem_wdata[64]~2 (
	.dataa(!seq_wdp_ovride),
	.datab(!q_b_64),
	.datac(!dgwb_wdata_88),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[64]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[64]~2 .extended_lut = "off";
defparam \mem_wdata[64]~2 .lut_mask = 64'h2727272727272727;
defparam \mem_wdata[64]~2 .shared_arith = "off";

dffeas \mem_wdata_r1[64] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[64]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[64]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[64] .is_wysiwyg = "true";
defparam \mem_wdata_r1[64] .power_up = "low";

dffeas \mem_wdata_r2[64] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[64]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[64]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[64] .is_wysiwyg = "true";
defparam \mem_wdata_r2[64] .power_up = "low";

arriaii_lcell_comb \mem_wdata[0]~3 (
	.dataa(!seq_wdp_ovride),
	.datab(!q_b_0),
	.datac(!dgwb_wdata_24),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[0]~3 .extended_lut = "off";
defparam \mem_wdata[0]~3 .lut_mask = 64'h2727272727272727;
defparam \mem_wdata[0]~3 .shared_arith = "off";

dffeas \mem_wdata_r1[0] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[0]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[0]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[0] .is_wysiwyg = "true";
defparam \mem_wdata_r1[0] .power_up = "low";

dffeas \mem_wdata_r2[0] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[0]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[0] .is_wysiwyg = "true";
defparam \mem_wdata_r2[0] .power_up = "low";

dffeas \wdata_valid_1x_r1[8] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_valid[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r1[8]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r1[8] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r1[8] .power_up = "low";

dffeas \wdata_valid_1x_r2[8] (
	.clk(phy_clk_1x),
	.d(\wdata_valid_1x_r1[8]~q ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r2[8]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r2[8] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r2[8] .power_up = "low";

dffeas \wdata_valid_1x_r1[0] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_valid[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r1[0]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r1[0] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r1[0] .power_up = "low";

dffeas \wdata_valid_1x_r2[0] (
	.clk(phy_clk_1x),
	.d(\wdata_valid_1x_r1[0]~q ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r2[0]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r2[0] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r2[0] .power_up = "low";

arriaii_lcell_comb \mem_wdata[97]~4 (
	.dataa(!seq_wdp_ovride),
	.datab(!q_b_97),
	.datac(!dgwb_wdata_121),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[97]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[97]~4 .extended_lut = "off";
defparam \mem_wdata[97]~4 .lut_mask = 64'h2727272727272727;
defparam \mem_wdata[97]~4 .shared_arith = "off";

dffeas \mem_wdata_r1[97] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[97]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[97]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[97] .is_wysiwyg = "true";
defparam \mem_wdata_r1[97] .power_up = "low";

dffeas \mem_wdata_r2[97] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[97]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[97]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[97] .is_wysiwyg = "true";
defparam \mem_wdata_r2[97] .power_up = "low";

arriaii_lcell_comb \mem_wdata[33]~5 (
	.dataa(!seq_wdp_ovride),
	.datab(!q_b_33),
	.datac(!dgwb_wdata_57),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[33]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[33]~5 .extended_lut = "off";
defparam \mem_wdata[33]~5 .lut_mask = 64'h2727272727272727;
defparam \mem_wdata[33]~5 .shared_arith = "off";

dffeas \mem_wdata_r1[33] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[33]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[33]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[33] .is_wysiwyg = "true";
defparam \mem_wdata_r1[33] .power_up = "low";

dffeas \mem_wdata_r2[33] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[33]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[33]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[33] .is_wysiwyg = "true";
defparam \mem_wdata_r2[33] .power_up = "low";

arriaii_lcell_comb \mem_wdata[65]~6 (
	.dataa(!seq_wdp_ovride),
	.datab(!q_b_65),
	.datac(!dgwb_wdata_89),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[65]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[65]~6 .extended_lut = "off";
defparam \mem_wdata[65]~6 .lut_mask = 64'h2727272727272727;
defparam \mem_wdata[65]~6 .shared_arith = "off";

dffeas \mem_wdata_r1[65] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[65]~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[65]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[65] .is_wysiwyg = "true";
defparam \mem_wdata_r1[65] .power_up = "low";

dffeas \mem_wdata_r2[65] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[65]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[65]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[65] .is_wysiwyg = "true";
defparam \mem_wdata_r2[65] .power_up = "low";

arriaii_lcell_comb \mem_wdata[1]~7 (
	.dataa(!seq_wdp_ovride),
	.datab(!q_b_1),
	.datac(!dgwb_wdata_25),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[1]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[1]~7 .extended_lut = "off";
defparam \mem_wdata[1]~7 .lut_mask = 64'h2727272727272727;
defparam \mem_wdata[1]~7 .shared_arith = "off";

dffeas \mem_wdata_r1[1] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[1]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[1]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[1] .is_wysiwyg = "true";
defparam \mem_wdata_r1[1] .power_up = "low";

dffeas \mem_wdata_r2[1] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[1]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[1] .is_wysiwyg = "true";
defparam \mem_wdata_r2[1] .power_up = "low";

arriaii_lcell_comb \mem_wdata[98]~8 (
	.dataa(!seq_wdp_ovride),
	.datab(!q_b_98),
	.datac(!dgwb_wdata_122),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[98]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[98]~8 .extended_lut = "off";
defparam \mem_wdata[98]~8 .lut_mask = 64'h2727272727272727;
defparam \mem_wdata[98]~8 .shared_arith = "off";

dffeas \mem_wdata_r1[98] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[98]~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[98]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[98] .is_wysiwyg = "true";
defparam \mem_wdata_r1[98] .power_up = "low";

dffeas \mem_wdata_r2[98] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[98]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[98]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[98] .is_wysiwyg = "true";
defparam \mem_wdata_r2[98] .power_up = "low";

arriaii_lcell_comb \mem_wdata[34]~9 (
	.dataa(!seq_wdp_ovride),
	.datab(!q_b_34),
	.datac(!dgwb_wdata_58),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[34]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[34]~9 .extended_lut = "off";
defparam \mem_wdata[34]~9 .lut_mask = 64'h2727272727272727;
defparam \mem_wdata[34]~9 .shared_arith = "off";

dffeas \mem_wdata_r1[34] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[34]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[34]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[34] .is_wysiwyg = "true";
defparam \mem_wdata_r1[34] .power_up = "low";

dffeas \mem_wdata_r2[34] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[34]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[34]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[34] .is_wysiwyg = "true";
defparam \mem_wdata_r2[34] .power_up = "low";

arriaii_lcell_comb \mem_wdata[66]~10 (
	.dataa(!seq_wdp_ovride),
	.datab(!q_b_66),
	.datac(!dgwb_wdata_90),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[66]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[66]~10 .extended_lut = "off";
defparam \mem_wdata[66]~10 .lut_mask = 64'h2727272727272727;
defparam \mem_wdata[66]~10 .shared_arith = "off";

dffeas \mem_wdata_r1[66] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[66]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[66]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[66] .is_wysiwyg = "true";
defparam \mem_wdata_r1[66] .power_up = "low";

dffeas \mem_wdata_r2[66] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[66]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[66]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[66] .is_wysiwyg = "true";
defparam \mem_wdata_r2[66] .power_up = "low";

arriaii_lcell_comb \mem_wdata[2]~11 (
	.dataa(!seq_wdp_ovride),
	.datab(!q_b_2),
	.datac(!dgwb_wdata_26),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[2]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[2]~11 .extended_lut = "off";
defparam \mem_wdata[2]~11 .lut_mask = 64'h2727272727272727;
defparam \mem_wdata[2]~11 .shared_arith = "off";

dffeas \mem_wdata_r1[2] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[2]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[2]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[2] .is_wysiwyg = "true";
defparam \mem_wdata_r1[2] .power_up = "low";

dffeas \mem_wdata_r2[2] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[2]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[2] .is_wysiwyg = "true";
defparam \mem_wdata_r2[2] .power_up = "low";

arriaii_lcell_comb \mem_wdata[99]~12 (
	.dataa(!seq_wdp_ovride),
	.datab(!q_b_99),
	.datac(!dgwb_wdata_123),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[99]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[99]~12 .extended_lut = "off";
defparam \mem_wdata[99]~12 .lut_mask = 64'h2727272727272727;
defparam \mem_wdata[99]~12 .shared_arith = "off";

dffeas \mem_wdata_r1[99] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[99]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[99]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[99] .is_wysiwyg = "true";
defparam \mem_wdata_r1[99] .power_up = "low";

dffeas \mem_wdata_r2[99] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[99]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[99]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[99] .is_wysiwyg = "true";
defparam \mem_wdata_r2[99] .power_up = "low";

arriaii_lcell_comb \mem_wdata[35]~13 (
	.dataa(!seq_wdp_ovride),
	.datab(!q_b_35),
	.datac(!dgwb_wdata_59),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[35]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[35]~13 .extended_lut = "off";
defparam \mem_wdata[35]~13 .lut_mask = 64'h2727272727272727;
defparam \mem_wdata[35]~13 .shared_arith = "off";

dffeas \mem_wdata_r1[35] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[35]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[35]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[35] .is_wysiwyg = "true";
defparam \mem_wdata_r1[35] .power_up = "low";

dffeas \mem_wdata_r2[35] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[35]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[35]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[35] .is_wysiwyg = "true";
defparam \mem_wdata_r2[35] .power_up = "low";

arriaii_lcell_comb \mem_wdata[67]~14 (
	.dataa(!seq_wdp_ovride),
	.datab(!q_b_67),
	.datac(!dgwb_wdata_91),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[67]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[67]~14 .extended_lut = "off";
defparam \mem_wdata[67]~14 .lut_mask = 64'h2727272727272727;
defparam \mem_wdata[67]~14 .shared_arith = "off";

dffeas \mem_wdata_r1[67] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[67]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[67]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[67] .is_wysiwyg = "true";
defparam \mem_wdata_r1[67] .power_up = "low";

dffeas \mem_wdata_r2[67] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[67]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[67]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[67] .is_wysiwyg = "true";
defparam \mem_wdata_r2[67] .power_up = "low";

arriaii_lcell_comb \mem_wdata[3]~15 (
	.dataa(!seq_wdp_ovride),
	.datab(!q_b_3),
	.datac(!dgwb_wdata_27),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[3]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[3]~15 .extended_lut = "off";
defparam \mem_wdata[3]~15 .lut_mask = 64'h2727272727272727;
defparam \mem_wdata[3]~15 .shared_arith = "off";

dffeas \mem_wdata_r1[3] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[3]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[3]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[3] .is_wysiwyg = "true";
defparam \mem_wdata_r1[3] .power_up = "low";

dffeas \mem_wdata_r2[3] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[3]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[3] .is_wysiwyg = "true";
defparam \mem_wdata_r2[3] .power_up = "low";

arriaii_lcell_comb \mem_wdata[100]~16 (
	.dataa(!seq_wdp_ovride),
	.datab(!q_b_100),
	.datac(!dgwb_wdata_124),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[100]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[100]~16 .extended_lut = "off";
defparam \mem_wdata[100]~16 .lut_mask = 64'h2727272727272727;
defparam \mem_wdata[100]~16 .shared_arith = "off";

dffeas \mem_wdata_r1[100] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[100]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[100]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[100] .is_wysiwyg = "true";
defparam \mem_wdata_r1[100] .power_up = "low";

dffeas \mem_wdata_r2[100] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[100]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[100]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[100] .is_wysiwyg = "true";
defparam \mem_wdata_r2[100] .power_up = "low";

arriaii_lcell_comb \mem_wdata[36]~17 (
	.dataa(!seq_wdp_ovride),
	.datab(!q_b_36),
	.datac(!dgwb_wdata_60),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[36]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[36]~17 .extended_lut = "off";
defparam \mem_wdata[36]~17 .lut_mask = 64'h2727272727272727;
defparam \mem_wdata[36]~17 .shared_arith = "off";

dffeas \mem_wdata_r1[36] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[36]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[36]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[36] .is_wysiwyg = "true";
defparam \mem_wdata_r1[36] .power_up = "low";

dffeas \mem_wdata_r2[36] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[36]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[36]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[36] .is_wysiwyg = "true";
defparam \mem_wdata_r2[36] .power_up = "low";

dffeas \wdata_valid_1x_r[1] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_valid[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r[1]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r[1] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r[1] .power_up = "low";

dffeas \wdata_valid_2x_r1[1] (
	.clk(write_clk_2x),
	.d(\wdata_valid_1x_r[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_2x_r1[1]~q ),
	.prn(vcc));
defparam \wdata_valid_2x_r1[1] .is_wysiwyg = "true";
defparam \wdata_valid_2x_r1[1] .power_up = "low";

dffeas \wdata_valid_2x_r2[1] (
	.clk(write_clk_2x),
	.d(\wdata_valid_2x_r1[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_2x_r2[1]~q ),
	.prn(vcc));
defparam \wdata_valid_2x_r2[1] .is_wysiwyg = "true";
defparam \wdata_valid_2x_r2[1] .power_up = "low";

arriaii_lcell_comb \wdata_sel~1 (
	.dataa(!\wdata_sel[1]~q ),
	.datab(!\wdata_valid_2x_r2[1]~q ),
	.datac(!\wdata_valid_2x_r1[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wdata_sel~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wdata_sel~1 .extended_lut = "off";
defparam \wdata_sel~1 .lut_mask = 64'hA2A2A2A2A2A2A2A2;
defparam \wdata_sel~1 .shared_arith = "off";

dffeas \wdata_sel[1] (
	.clk(write_clk_2x),
	.d(\wdata_sel~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_sel[1]~q ),
	.prn(vcc));
defparam \wdata_sel[1] .is_wysiwyg = "true";
defparam \wdata_sel[1] .power_up = "low";

arriaii_lcell_comb \mem_wdata[68]~18 (
	.dataa(!seq_wdp_ovride),
	.datab(!q_b_68),
	.datac(!dgwb_wdata_92),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[68]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[68]~18 .extended_lut = "off";
defparam \mem_wdata[68]~18 .lut_mask = 64'h2727272727272727;
defparam \mem_wdata[68]~18 .shared_arith = "off";

dffeas \mem_wdata_r1[68] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[68]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[68]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[68] .is_wysiwyg = "true";
defparam \mem_wdata_r1[68] .power_up = "low";

dffeas \mem_wdata_r2[68] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[68]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[68]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[68] .is_wysiwyg = "true";
defparam \mem_wdata_r2[68] .power_up = "low";

arriaii_lcell_comb \mem_wdata[4]~19 (
	.dataa(!seq_wdp_ovride),
	.datab(!q_b_4),
	.datac(!dgwb_wdata_28),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[4]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[4]~19 .extended_lut = "off";
defparam \mem_wdata[4]~19 .lut_mask = 64'h2727272727272727;
defparam \mem_wdata[4]~19 .shared_arith = "off";

dffeas \mem_wdata_r1[4] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[4]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[4]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[4] .is_wysiwyg = "true";
defparam \mem_wdata_r1[4] .power_up = "low";

dffeas \mem_wdata_r2[4] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[4]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[4] .is_wysiwyg = "true";
defparam \mem_wdata_r2[4] .power_up = "low";

dffeas \wdata_valid_1x_r1[9] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_valid[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r1[9]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r1[9] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r1[9] .power_up = "low";

dffeas \wdata_valid_1x_r2[9] (
	.clk(phy_clk_1x),
	.d(\wdata_valid_1x_r1[9]~q ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r2[9]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r2[9] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r2[9] .power_up = "low";

dffeas \wdata_valid_1x_r1[1] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_valid[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r1[1]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r1[1] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r1[1] .power_up = "low";

dffeas \wdata_valid_1x_r2[1] (
	.clk(phy_clk_1x),
	.d(\wdata_valid_1x_r1[1]~q ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r2[1]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r2[1] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r2[1] .power_up = "low";

arriaii_lcell_comb \mem_wdata[101]~20 (
	.dataa(!seq_wdp_ovride),
	.datab(!q_b_101),
	.datac(!dgwb_wdata_125),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[101]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[101]~20 .extended_lut = "off";
defparam \mem_wdata[101]~20 .lut_mask = 64'h2727272727272727;
defparam \mem_wdata[101]~20 .shared_arith = "off";

dffeas \mem_wdata_r1[101] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[101]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[101]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[101] .is_wysiwyg = "true";
defparam \mem_wdata_r1[101] .power_up = "low";

dffeas \mem_wdata_r2[101] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[101]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[101]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[101] .is_wysiwyg = "true";
defparam \mem_wdata_r2[101] .power_up = "low";

arriaii_lcell_comb \mem_wdata[37]~21 (
	.dataa(!seq_wdp_ovride),
	.datab(!q_b_37),
	.datac(!dgwb_wdata_61),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[37]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[37]~21 .extended_lut = "off";
defparam \mem_wdata[37]~21 .lut_mask = 64'h2727272727272727;
defparam \mem_wdata[37]~21 .shared_arith = "off";

dffeas \mem_wdata_r1[37] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[37]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[37]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[37] .is_wysiwyg = "true";
defparam \mem_wdata_r1[37] .power_up = "low";

dffeas \mem_wdata_r2[37] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[37]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[37]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[37] .is_wysiwyg = "true";
defparam \mem_wdata_r2[37] .power_up = "low";

arriaii_lcell_comb \mem_wdata[69]~22 (
	.dataa(!seq_wdp_ovride),
	.datab(!q_b_69),
	.datac(!dgwb_wdata_93),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[69]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[69]~22 .extended_lut = "off";
defparam \mem_wdata[69]~22 .lut_mask = 64'h2727272727272727;
defparam \mem_wdata[69]~22 .shared_arith = "off";

dffeas \mem_wdata_r1[69] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[69]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[69]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[69] .is_wysiwyg = "true";
defparam \mem_wdata_r1[69] .power_up = "low";

dffeas \mem_wdata_r2[69] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[69]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[69]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[69] .is_wysiwyg = "true";
defparam \mem_wdata_r2[69] .power_up = "low";

arriaii_lcell_comb \mem_wdata[5]~23 (
	.dataa(!seq_wdp_ovride),
	.datab(!q_b_5),
	.datac(!dgwb_wdata_29),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[5]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[5]~23 .extended_lut = "off";
defparam \mem_wdata[5]~23 .lut_mask = 64'h2727272727272727;
defparam \mem_wdata[5]~23 .shared_arith = "off";

dffeas \mem_wdata_r1[5] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[5]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[5]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[5] .is_wysiwyg = "true";
defparam \mem_wdata_r1[5] .power_up = "low";

dffeas \mem_wdata_r2[5] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[5]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[5] .is_wysiwyg = "true";
defparam \mem_wdata_r2[5] .power_up = "low";

arriaii_lcell_comb \mem_wdata[102]~24 (
	.dataa(!seq_wdp_ovride),
	.datab(!q_b_102),
	.datac(!dgwb_wdata_126),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[102]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[102]~24 .extended_lut = "off";
defparam \mem_wdata[102]~24 .lut_mask = 64'h2727272727272727;
defparam \mem_wdata[102]~24 .shared_arith = "off";

dffeas \mem_wdata_r1[102] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[102]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[102]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[102] .is_wysiwyg = "true";
defparam \mem_wdata_r1[102] .power_up = "low";

dffeas \mem_wdata_r2[102] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[102]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[102]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[102] .is_wysiwyg = "true";
defparam \mem_wdata_r2[102] .power_up = "low";

arriaii_lcell_comb \mem_wdata[38]~25 (
	.dataa(!seq_wdp_ovride),
	.datab(!q_b_38),
	.datac(!dgwb_wdata_62),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[38]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[38]~25 .extended_lut = "off";
defparam \mem_wdata[38]~25 .lut_mask = 64'h2727272727272727;
defparam \mem_wdata[38]~25 .shared_arith = "off";

dffeas \mem_wdata_r1[38] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[38]~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[38]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[38] .is_wysiwyg = "true";
defparam \mem_wdata_r1[38] .power_up = "low";

dffeas \mem_wdata_r2[38] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[38]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[38]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[38] .is_wysiwyg = "true";
defparam \mem_wdata_r2[38] .power_up = "low";

arriaii_lcell_comb \mem_wdata[70]~26 (
	.dataa(!seq_wdp_ovride),
	.datab(!q_b_70),
	.datac(!dgwb_wdata_94),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[70]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[70]~26 .extended_lut = "off";
defparam \mem_wdata[70]~26 .lut_mask = 64'h2727272727272727;
defparam \mem_wdata[70]~26 .shared_arith = "off";

dffeas \mem_wdata_r1[70] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[70]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[70]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[70] .is_wysiwyg = "true";
defparam \mem_wdata_r1[70] .power_up = "low";

dffeas \mem_wdata_r2[70] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[70]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[70]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[70] .is_wysiwyg = "true";
defparam \mem_wdata_r2[70] .power_up = "low";

arriaii_lcell_comb \mem_wdata[6]~27 (
	.dataa(!seq_wdp_ovride),
	.datab(!q_b_6),
	.datac(!dgwb_wdata_30),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[6]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[6]~27 .extended_lut = "off";
defparam \mem_wdata[6]~27 .lut_mask = 64'h2727272727272727;
defparam \mem_wdata[6]~27 .shared_arith = "off";

dffeas \mem_wdata_r1[6] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[6]~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[6]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[6] .is_wysiwyg = "true";
defparam \mem_wdata_r1[6] .power_up = "low";

dffeas \mem_wdata_r2[6] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[6]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[6] .is_wysiwyg = "true";
defparam \mem_wdata_r2[6] .power_up = "low";

arriaii_lcell_comb \mem_wdata[103]~28 (
	.dataa(!seq_wdp_ovride),
	.datab(!q_b_103),
	.datac(!dgwb_wdata_127),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[103]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[103]~28 .extended_lut = "off";
defparam \mem_wdata[103]~28 .lut_mask = 64'h2727272727272727;
defparam \mem_wdata[103]~28 .shared_arith = "off";

dffeas \mem_wdata_r1[103] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[103]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[103]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[103] .is_wysiwyg = "true";
defparam \mem_wdata_r1[103] .power_up = "low";

dffeas \mem_wdata_r2[103] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[103]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[103]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[103] .is_wysiwyg = "true";
defparam \mem_wdata_r2[103] .power_up = "low";

arriaii_lcell_comb \mem_wdata[39]~29 (
	.dataa(!seq_wdp_ovride),
	.datab(!q_b_39),
	.datac(!dgwb_wdata_63),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[39]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[39]~29 .extended_lut = "off";
defparam \mem_wdata[39]~29 .lut_mask = 64'h2727272727272727;
defparam \mem_wdata[39]~29 .shared_arith = "off";

dffeas \mem_wdata_r1[39] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[39]~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[39]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[39] .is_wysiwyg = "true";
defparam \mem_wdata_r1[39] .power_up = "low";

dffeas \mem_wdata_r2[39] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[39]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[39]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[39] .is_wysiwyg = "true";
defparam \mem_wdata_r2[39] .power_up = "low";

arriaii_lcell_comb \mem_wdata[71]~30 (
	.dataa(!seq_wdp_ovride),
	.datab(!q_b_71),
	.datac(!dgwb_wdata_95),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[71]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[71]~30 .extended_lut = "off";
defparam \mem_wdata[71]~30 .lut_mask = 64'h2727272727272727;
defparam \mem_wdata[71]~30 .shared_arith = "off";

dffeas \mem_wdata_r1[71] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[71]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[71]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[71] .is_wysiwyg = "true";
defparam \mem_wdata_r1[71] .power_up = "low";

dffeas \mem_wdata_r2[71] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[71]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[71]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[71] .is_wysiwyg = "true";
defparam \mem_wdata_r2[71] .power_up = "low";

arriaii_lcell_comb \mem_wdata[7]~31 (
	.dataa(!seq_wdp_ovride),
	.datab(!q_b_7),
	.datac(!dgwb_wdata_31),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[7]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[7]~31 .extended_lut = "off";
defparam \mem_wdata[7]~31 .lut_mask = 64'h2727272727272727;
defparam \mem_wdata[7]~31 .shared_arith = "off";

dffeas \mem_wdata_r1[7] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[7]~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[7]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[7] .is_wysiwyg = "true";
defparam \mem_wdata_r1[7] .power_up = "low";

dffeas \mem_wdata_r2[7] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[7]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[7] .is_wysiwyg = "true";
defparam \mem_wdata_r2[7] .power_up = "low";

arriaii_lcell_comb \mem_wdata[104]~32 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_120),
	.datac(!q_b_104),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[104]~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[104]~32 .extended_lut = "off";
defparam \mem_wdata[104]~32 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[104]~32 .shared_arith = "off";

dffeas \mem_wdata_r1[104] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[104]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[104]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[104] .is_wysiwyg = "true";
defparam \mem_wdata_r1[104] .power_up = "low";

dffeas \mem_wdata_r2[104] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[104]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[104]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[104] .is_wysiwyg = "true";
defparam \mem_wdata_r2[104] .power_up = "low";

arriaii_lcell_comb \mem_wdata[40]~33 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_56),
	.datac(!q_b_40),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[40]~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[40]~33 .extended_lut = "off";
defparam \mem_wdata[40]~33 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[40]~33 .shared_arith = "off";

dffeas \mem_wdata_r1[40] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[40]~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[40]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[40] .is_wysiwyg = "true";
defparam \mem_wdata_r1[40] .power_up = "low";

dffeas \mem_wdata_r2[40] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[40]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[40]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[40] .is_wysiwyg = "true";
defparam \mem_wdata_r2[40] .power_up = "low";

dffeas \wdata_valid_1x_r[2] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_valid[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r[2]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r[2] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r[2] .power_up = "low";

dffeas \wdata_valid_2x_r1[2] (
	.clk(write_clk_2x),
	.d(\wdata_valid_1x_r[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_2x_r1[2]~q ),
	.prn(vcc));
defparam \wdata_valid_2x_r1[2] .is_wysiwyg = "true";
defparam \wdata_valid_2x_r1[2] .power_up = "low";

dffeas \wdata_valid_2x_r2[2] (
	.clk(write_clk_2x),
	.d(\wdata_valid_2x_r1[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_2x_r2[2]~q ),
	.prn(vcc));
defparam \wdata_valid_2x_r2[2] .is_wysiwyg = "true";
defparam \wdata_valid_2x_r2[2] .power_up = "low";

arriaii_lcell_comb \wdata_sel~2 (
	.dataa(!\wdata_sel[2]~q ),
	.datab(!\wdata_valid_2x_r2[2]~q ),
	.datac(!\wdata_valid_2x_r1[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wdata_sel~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wdata_sel~2 .extended_lut = "off";
defparam \wdata_sel~2 .lut_mask = 64'hA2A2A2A2A2A2A2A2;
defparam \wdata_sel~2 .shared_arith = "off";

dffeas \wdata_sel[2] (
	.clk(write_clk_2x),
	.d(\wdata_sel~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_sel[2]~q ),
	.prn(vcc));
defparam \wdata_sel[2] .is_wysiwyg = "true";
defparam \wdata_sel[2] .power_up = "low";

arriaii_lcell_comb \mem_wdata[72]~34 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_88),
	.datac(!q_b_72),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[72]~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[72]~34 .extended_lut = "off";
defparam \mem_wdata[72]~34 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[72]~34 .shared_arith = "off";

dffeas \mem_wdata_r1[72] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[72]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[72]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[72] .is_wysiwyg = "true";
defparam \mem_wdata_r1[72] .power_up = "low";

dffeas \mem_wdata_r2[72] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[72]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[72]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[72] .is_wysiwyg = "true";
defparam \mem_wdata_r2[72] .power_up = "low";

arriaii_lcell_comb \mem_wdata[8]~35 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_24),
	.datac(!q_b_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[8]~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[8]~35 .extended_lut = "off";
defparam \mem_wdata[8]~35 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[8]~35 .shared_arith = "off";

dffeas \mem_wdata_r1[8] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[8]~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[8]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[8] .is_wysiwyg = "true";
defparam \mem_wdata_r1[8] .power_up = "low";

dffeas \mem_wdata_r2[8] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[8]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[8] .is_wysiwyg = "true";
defparam \mem_wdata_r2[8] .power_up = "low";

dffeas \wdata_valid_1x_r1[10] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_valid[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r1[10]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r1[10] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r1[10] .power_up = "low";

dffeas \wdata_valid_1x_r2[10] (
	.clk(phy_clk_1x),
	.d(\wdata_valid_1x_r1[10]~q ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r2[10]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r2[10] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r2[10] .power_up = "low";

dffeas \wdata_valid_1x_r1[2] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_valid[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r1[2]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r1[2] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r1[2] .power_up = "low";

dffeas \wdata_valid_1x_r2[2] (
	.clk(phy_clk_1x),
	.d(\wdata_valid_1x_r1[2]~q ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r2[2]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r2[2] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r2[2] .power_up = "low";

arriaii_lcell_comb \mem_wdata[105]~36 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_121),
	.datac(!q_b_105),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[105]~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[105]~36 .extended_lut = "off";
defparam \mem_wdata[105]~36 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[105]~36 .shared_arith = "off";

dffeas \mem_wdata_r1[105] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[105]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[105]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[105] .is_wysiwyg = "true";
defparam \mem_wdata_r1[105] .power_up = "low";

dffeas \mem_wdata_r2[105] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[105]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[105]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[105] .is_wysiwyg = "true";
defparam \mem_wdata_r2[105] .power_up = "low";

arriaii_lcell_comb \mem_wdata[41]~37 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_57),
	.datac(!q_b_41),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[41]~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[41]~37 .extended_lut = "off";
defparam \mem_wdata[41]~37 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[41]~37 .shared_arith = "off";

dffeas \mem_wdata_r1[41] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[41]~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[41]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[41] .is_wysiwyg = "true";
defparam \mem_wdata_r1[41] .power_up = "low";

dffeas \mem_wdata_r2[41] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[41]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[41]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[41] .is_wysiwyg = "true";
defparam \mem_wdata_r2[41] .power_up = "low";

arriaii_lcell_comb \mem_wdata[73]~38 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_89),
	.datac(!q_b_73),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[73]~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[73]~38 .extended_lut = "off";
defparam \mem_wdata[73]~38 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[73]~38 .shared_arith = "off";

dffeas \mem_wdata_r1[73] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[73]~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[73]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[73] .is_wysiwyg = "true";
defparam \mem_wdata_r1[73] .power_up = "low";

dffeas \mem_wdata_r2[73] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[73]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[73]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[73] .is_wysiwyg = "true";
defparam \mem_wdata_r2[73] .power_up = "low";

arriaii_lcell_comb \mem_wdata[9]~39 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_25),
	.datac(!q_b_9),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[9]~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[9]~39 .extended_lut = "off";
defparam \mem_wdata[9]~39 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[9]~39 .shared_arith = "off";

dffeas \mem_wdata_r1[9] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[9]~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[9]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[9] .is_wysiwyg = "true";
defparam \mem_wdata_r1[9] .power_up = "low";

dffeas \mem_wdata_r2[9] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[9]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[9] .is_wysiwyg = "true";
defparam \mem_wdata_r2[9] .power_up = "low";

arriaii_lcell_comb \mem_wdata[106]~40 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_122),
	.datac(!q_b_106),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[106]~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[106]~40 .extended_lut = "off";
defparam \mem_wdata[106]~40 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[106]~40 .shared_arith = "off";

dffeas \mem_wdata_r1[106] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[106]~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[106]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[106] .is_wysiwyg = "true";
defparam \mem_wdata_r1[106] .power_up = "low";

dffeas \mem_wdata_r2[106] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[106]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[106]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[106] .is_wysiwyg = "true";
defparam \mem_wdata_r2[106] .power_up = "low";

arriaii_lcell_comb \mem_wdata[42]~41 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_58),
	.datac(!q_b_42),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[42]~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[42]~41 .extended_lut = "off";
defparam \mem_wdata[42]~41 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[42]~41 .shared_arith = "off";

dffeas \mem_wdata_r1[42] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[42]~41_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[42]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[42] .is_wysiwyg = "true";
defparam \mem_wdata_r1[42] .power_up = "low";

dffeas \mem_wdata_r2[42] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[42]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[42]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[42] .is_wysiwyg = "true";
defparam \mem_wdata_r2[42] .power_up = "low";

arriaii_lcell_comb \mem_wdata[74]~42 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_90),
	.datac(!q_b_74),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[74]~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[74]~42 .extended_lut = "off";
defparam \mem_wdata[74]~42 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[74]~42 .shared_arith = "off";

dffeas \mem_wdata_r1[74] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[74]~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[74]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[74] .is_wysiwyg = "true";
defparam \mem_wdata_r1[74] .power_up = "low";

dffeas \mem_wdata_r2[74] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[74]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[74]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[74] .is_wysiwyg = "true";
defparam \mem_wdata_r2[74] .power_up = "low";

arriaii_lcell_comb \mem_wdata[10]~43 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_26),
	.datac(!q_b_10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[10]~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[10]~43 .extended_lut = "off";
defparam \mem_wdata[10]~43 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[10]~43 .shared_arith = "off";

dffeas \mem_wdata_r1[10] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[10]~43_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[10]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[10] .is_wysiwyg = "true";
defparam \mem_wdata_r1[10] .power_up = "low";

dffeas \mem_wdata_r2[10] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[10]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[10] .is_wysiwyg = "true";
defparam \mem_wdata_r2[10] .power_up = "low";

arriaii_lcell_comb \mem_wdata[107]~44 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_123),
	.datac(!q_b_107),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[107]~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[107]~44 .extended_lut = "off";
defparam \mem_wdata[107]~44 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[107]~44 .shared_arith = "off";

dffeas \mem_wdata_r1[107] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[107]~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[107]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[107] .is_wysiwyg = "true";
defparam \mem_wdata_r1[107] .power_up = "low";

dffeas \mem_wdata_r2[107] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[107]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[107]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[107] .is_wysiwyg = "true";
defparam \mem_wdata_r2[107] .power_up = "low";

arriaii_lcell_comb \mem_wdata[43]~45 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_59),
	.datac(!q_b_43),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[43]~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[43]~45 .extended_lut = "off";
defparam \mem_wdata[43]~45 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[43]~45 .shared_arith = "off";

dffeas \mem_wdata_r1[43] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[43]~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[43]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[43] .is_wysiwyg = "true";
defparam \mem_wdata_r1[43] .power_up = "low";

dffeas \mem_wdata_r2[43] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[43]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[43]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[43] .is_wysiwyg = "true";
defparam \mem_wdata_r2[43] .power_up = "low";

arriaii_lcell_comb \mem_wdata[75]~46 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_91),
	.datac(!q_b_75),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[75]~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[75]~46 .extended_lut = "off";
defparam \mem_wdata[75]~46 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[75]~46 .shared_arith = "off";

dffeas \mem_wdata_r1[75] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[75]~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[75]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[75] .is_wysiwyg = "true";
defparam \mem_wdata_r1[75] .power_up = "low";

dffeas \mem_wdata_r2[75] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[75]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[75]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[75] .is_wysiwyg = "true";
defparam \mem_wdata_r2[75] .power_up = "low";

arriaii_lcell_comb \mem_wdata[11]~47 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_27),
	.datac(!q_b_11),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[11]~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[11]~47 .extended_lut = "off";
defparam \mem_wdata[11]~47 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[11]~47 .shared_arith = "off";

dffeas \mem_wdata_r1[11] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[11]~47_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[11]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[11] .is_wysiwyg = "true";
defparam \mem_wdata_r1[11] .power_up = "low";

dffeas \mem_wdata_r2[11] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[11]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[11] .is_wysiwyg = "true";
defparam \mem_wdata_r2[11] .power_up = "low";

arriaii_lcell_comb \mem_wdata[108]~48 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_124),
	.datac(!q_b_108),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[108]~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[108]~48 .extended_lut = "off";
defparam \mem_wdata[108]~48 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[108]~48 .shared_arith = "off";

dffeas \mem_wdata_r1[108] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[108]~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[108]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[108] .is_wysiwyg = "true";
defparam \mem_wdata_r1[108] .power_up = "low";

dffeas \mem_wdata_r2[108] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[108]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[108]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[108] .is_wysiwyg = "true";
defparam \mem_wdata_r2[108] .power_up = "low";

arriaii_lcell_comb \mem_wdata[44]~49 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_60),
	.datac(!q_b_44),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[44]~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[44]~49 .extended_lut = "off";
defparam \mem_wdata[44]~49 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[44]~49 .shared_arith = "off";

dffeas \mem_wdata_r1[44] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[44]~49_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[44]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[44] .is_wysiwyg = "true";
defparam \mem_wdata_r1[44] .power_up = "low";

dffeas \mem_wdata_r2[44] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[44]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[44]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[44] .is_wysiwyg = "true";
defparam \mem_wdata_r2[44] .power_up = "low";

dffeas \wdata_valid_1x_r[3] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_valid[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r[3]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r[3] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r[3] .power_up = "low";

dffeas \wdata_valid_2x_r1[3] (
	.clk(write_clk_2x),
	.d(\wdata_valid_1x_r[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_2x_r1[3]~q ),
	.prn(vcc));
defparam \wdata_valid_2x_r1[3] .is_wysiwyg = "true";
defparam \wdata_valid_2x_r1[3] .power_up = "low";

dffeas \wdata_valid_2x_r2[3] (
	.clk(write_clk_2x),
	.d(\wdata_valid_2x_r1[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_2x_r2[3]~q ),
	.prn(vcc));
defparam \wdata_valid_2x_r2[3] .is_wysiwyg = "true";
defparam \wdata_valid_2x_r2[3] .power_up = "low";

arriaii_lcell_comb \wdata_sel~3 (
	.dataa(!\wdata_sel[3]~q ),
	.datab(!\wdata_valid_2x_r2[3]~q ),
	.datac(!\wdata_valid_2x_r1[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wdata_sel~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wdata_sel~3 .extended_lut = "off";
defparam \wdata_sel~3 .lut_mask = 64'hA2A2A2A2A2A2A2A2;
defparam \wdata_sel~3 .shared_arith = "off";

dffeas \wdata_sel[3] (
	.clk(write_clk_2x),
	.d(\wdata_sel~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_sel[3]~q ),
	.prn(vcc));
defparam \wdata_sel[3] .is_wysiwyg = "true";
defparam \wdata_sel[3] .power_up = "low";

arriaii_lcell_comb \mem_wdata[76]~50 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_92),
	.datac(!q_b_76),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[76]~50_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[76]~50 .extended_lut = "off";
defparam \mem_wdata[76]~50 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[76]~50 .shared_arith = "off";

dffeas \mem_wdata_r1[76] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[76]~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[76]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[76] .is_wysiwyg = "true";
defparam \mem_wdata_r1[76] .power_up = "low";

dffeas \mem_wdata_r2[76] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[76]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[76]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[76] .is_wysiwyg = "true";
defparam \mem_wdata_r2[76] .power_up = "low";

arriaii_lcell_comb \mem_wdata[12]~51 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_28),
	.datac(!q_b_12),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[12]~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[12]~51 .extended_lut = "off";
defparam \mem_wdata[12]~51 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[12]~51 .shared_arith = "off";

dffeas \mem_wdata_r1[12] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[12]~51_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[12]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[12] .is_wysiwyg = "true";
defparam \mem_wdata_r1[12] .power_up = "low";

dffeas \mem_wdata_r2[12] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[12]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[12] .is_wysiwyg = "true";
defparam \mem_wdata_r2[12] .power_up = "low";

dffeas \wdata_valid_1x_r1[11] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_valid[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r1[11]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r1[11] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r1[11] .power_up = "low";

dffeas \wdata_valid_1x_r2[11] (
	.clk(phy_clk_1x),
	.d(\wdata_valid_1x_r1[11]~q ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r2[11]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r2[11] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r2[11] .power_up = "low";

dffeas \wdata_valid_1x_r1[3] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_valid[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r1[3]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r1[3] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r1[3] .power_up = "low";

dffeas \wdata_valid_1x_r2[3] (
	.clk(phy_clk_1x),
	.d(\wdata_valid_1x_r1[3]~q ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r2[3]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r2[3] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r2[3] .power_up = "low";

arriaii_lcell_comb \mem_wdata[109]~52 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_125),
	.datac(!q_b_109),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[109]~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[109]~52 .extended_lut = "off";
defparam \mem_wdata[109]~52 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[109]~52 .shared_arith = "off";

dffeas \mem_wdata_r1[109] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[109]~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[109]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[109] .is_wysiwyg = "true";
defparam \mem_wdata_r1[109] .power_up = "low";

dffeas \mem_wdata_r2[109] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[109]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[109]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[109] .is_wysiwyg = "true";
defparam \mem_wdata_r2[109] .power_up = "low";

arriaii_lcell_comb \mem_wdata[45]~53 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_61),
	.datac(!q_b_45),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[45]~53_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[45]~53 .extended_lut = "off";
defparam \mem_wdata[45]~53 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[45]~53 .shared_arith = "off";

dffeas \mem_wdata_r1[45] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[45]~53_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[45]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[45] .is_wysiwyg = "true";
defparam \mem_wdata_r1[45] .power_up = "low";

dffeas \mem_wdata_r2[45] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[45]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[45]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[45] .is_wysiwyg = "true";
defparam \mem_wdata_r2[45] .power_up = "low";

arriaii_lcell_comb \mem_wdata[77]~54 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_93),
	.datac(!q_b_77),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[77]~54_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[77]~54 .extended_lut = "off";
defparam \mem_wdata[77]~54 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[77]~54 .shared_arith = "off";

dffeas \mem_wdata_r1[77] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[77]~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[77]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[77] .is_wysiwyg = "true";
defparam \mem_wdata_r1[77] .power_up = "low";

dffeas \mem_wdata_r2[77] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[77]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[77]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[77] .is_wysiwyg = "true";
defparam \mem_wdata_r2[77] .power_up = "low";

arriaii_lcell_comb \mem_wdata[13]~55 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_29),
	.datac(!q_b_13),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[13]~55_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[13]~55 .extended_lut = "off";
defparam \mem_wdata[13]~55 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[13]~55 .shared_arith = "off";

dffeas \mem_wdata_r1[13] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[13]~55_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[13]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[13] .is_wysiwyg = "true";
defparam \mem_wdata_r1[13] .power_up = "low";

dffeas \mem_wdata_r2[13] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[13]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[13] .is_wysiwyg = "true";
defparam \mem_wdata_r2[13] .power_up = "low";

arriaii_lcell_comb \mem_wdata[110]~56 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_126),
	.datac(!q_b_110),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[110]~56_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[110]~56 .extended_lut = "off";
defparam \mem_wdata[110]~56 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[110]~56 .shared_arith = "off";

dffeas \mem_wdata_r1[110] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[110]~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[110]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[110] .is_wysiwyg = "true";
defparam \mem_wdata_r1[110] .power_up = "low";

dffeas \mem_wdata_r2[110] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[110]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[110]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[110] .is_wysiwyg = "true";
defparam \mem_wdata_r2[110] .power_up = "low";

arriaii_lcell_comb \mem_wdata[46]~57 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_62),
	.datac(!q_b_46),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[46]~57_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[46]~57 .extended_lut = "off";
defparam \mem_wdata[46]~57 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[46]~57 .shared_arith = "off";

dffeas \mem_wdata_r1[46] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[46]~57_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[46]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[46] .is_wysiwyg = "true";
defparam \mem_wdata_r1[46] .power_up = "low";

dffeas \mem_wdata_r2[46] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[46]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[46]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[46] .is_wysiwyg = "true";
defparam \mem_wdata_r2[46] .power_up = "low";

arriaii_lcell_comb \mem_wdata[78]~58 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_94),
	.datac(!q_b_78),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[78]~58_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[78]~58 .extended_lut = "off";
defparam \mem_wdata[78]~58 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[78]~58 .shared_arith = "off";

dffeas \mem_wdata_r1[78] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[78]~58_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[78]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[78] .is_wysiwyg = "true";
defparam \mem_wdata_r1[78] .power_up = "low";

dffeas \mem_wdata_r2[78] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[78]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[78]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[78] .is_wysiwyg = "true";
defparam \mem_wdata_r2[78] .power_up = "low";

arriaii_lcell_comb \mem_wdata[14]~59 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_30),
	.datac(!q_b_14),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[14]~59_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[14]~59 .extended_lut = "off";
defparam \mem_wdata[14]~59 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[14]~59 .shared_arith = "off";

dffeas \mem_wdata_r1[14] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[14]~59_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[14]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[14] .is_wysiwyg = "true";
defparam \mem_wdata_r1[14] .power_up = "low";

dffeas \mem_wdata_r2[14] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[14]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[14] .is_wysiwyg = "true";
defparam \mem_wdata_r2[14] .power_up = "low";

arriaii_lcell_comb \mem_wdata[111]~60 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_127),
	.datac(!q_b_111),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[111]~60_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[111]~60 .extended_lut = "off";
defparam \mem_wdata[111]~60 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[111]~60 .shared_arith = "off";

dffeas \mem_wdata_r1[111] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[111]~60_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[111]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[111] .is_wysiwyg = "true";
defparam \mem_wdata_r1[111] .power_up = "low";

dffeas \mem_wdata_r2[111] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[111]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[111]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[111] .is_wysiwyg = "true";
defparam \mem_wdata_r2[111] .power_up = "low";

arriaii_lcell_comb \mem_wdata[47]~61 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_63),
	.datac(!q_b_47),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[47]~61_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[47]~61 .extended_lut = "off";
defparam \mem_wdata[47]~61 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[47]~61 .shared_arith = "off";

dffeas \mem_wdata_r1[47] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[47]~61_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[47]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[47] .is_wysiwyg = "true";
defparam \mem_wdata_r1[47] .power_up = "low";

dffeas \mem_wdata_r2[47] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[47]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[47]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[47] .is_wysiwyg = "true";
defparam \mem_wdata_r2[47] .power_up = "low";

arriaii_lcell_comb \mem_wdata[79]~62 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_95),
	.datac(!q_b_79),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[79]~62_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[79]~62 .extended_lut = "off";
defparam \mem_wdata[79]~62 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[79]~62 .shared_arith = "off";

dffeas \mem_wdata_r1[79] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[79]~62_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[79]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[79] .is_wysiwyg = "true";
defparam \mem_wdata_r1[79] .power_up = "low";

dffeas \mem_wdata_r2[79] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[79]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[79]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[79] .is_wysiwyg = "true";
defparam \mem_wdata_r2[79] .power_up = "low";

arriaii_lcell_comb \mem_wdata[15]~63 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_31),
	.datac(!q_b_15),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[15]~63_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[15]~63 .extended_lut = "off";
defparam \mem_wdata[15]~63 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[15]~63 .shared_arith = "off";

dffeas \mem_wdata_r1[15] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[15]~63_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[15]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[15] .is_wysiwyg = "true";
defparam \mem_wdata_r1[15] .power_up = "low";

dffeas \mem_wdata_r2[15] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[15]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[15] .is_wysiwyg = "true";
defparam \mem_wdata_r2[15] .power_up = "low";

arriaii_lcell_comb \mem_wdata[112]~64 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_120),
	.datac(!q_b_112),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[112]~64_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[112]~64 .extended_lut = "off";
defparam \mem_wdata[112]~64 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[112]~64 .shared_arith = "off";

dffeas \mem_wdata_r1[112] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[112]~64_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[112]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[112] .is_wysiwyg = "true";
defparam \mem_wdata_r1[112] .power_up = "low";

dffeas \mem_wdata_r2[112] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[112]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[112]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[112] .is_wysiwyg = "true";
defparam \mem_wdata_r2[112] .power_up = "low";

arriaii_lcell_comb \mem_wdata[48]~65 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_56),
	.datac(!q_b_48),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[48]~65_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[48]~65 .extended_lut = "off";
defparam \mem_wdata[48]~65 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[48]~65 .shared_arith = "off";

dffeas \mem_wdata_r1[48] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[48]~65_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[48]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[48] .is_wysiwyg = "true";
defparam \mem_wdata_r1[48] .power_up = "low";

dffeas \mem_wdata_r2[48] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[48]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[48]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[48] .is_wysiwyg = "true";
defparam \mem_wdata_r2[48] .power_up = "low";

dffeas \wdata_valid_1x_r[4] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_valid[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r[4]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r[4] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r[4] .power_up = "low";

dffeas \wdata_valid_2x_r1[4] (
	.clk(write_clk_2x),
	.d(\wdata_valid_1x_r[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_2x_r1[4]~q ),
	.prn(vcc));
defparam \wdata_valid_2x_r1[4] .is_wysiwyg = "true";
defparam \wdata_valid_2x_r1[4] .power_up = "low";

dffeas \wdata_valid_2x_r2[4] (
	.clk(write_clk_2x),
	.d(\wdata_valid_2x_r1[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_2x_r2[4]~q ),
	.prn(vcc));
defparam \wdata_valid_2x_r2[4] .is_wysiwyg = "true";
defparam \wdata_valid_2x_r2[4] .power_up = "low";

arriaii_lcell_comb \wdata_sel~4 (
	.dataa(!\wdata_sel[4]~q ),
	.datab(!\wdata_valid_2x_r2[4]~q ),
	.datac(!\wdata_valid_2x_r1[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wdata_sel~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wdata_sel~4 .extended_lut = "off";
defparam \wdata_sel~4 .lut_mask = 64'hA2A2A2A2A2A2A2A2;
defparam \wdata_sel~4 .shared_arith = "off";

dffeas \wdata_sel[4] (
	.clk(write_clk_2x),
	.d(\wdata_sel~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_sel[4]~q ),
	.prn(vcc));
defparam \wdata_sel[4] .is_wysiwyg = "true";
defparam \wdata_sel[4] .power_up = "low";

arriaii_lcell_comb \mem_wdata[80]~66 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_88),
	.datac(!q_b_80),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[80]~66_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[80]~66 .extended_lut = "off";
defparam \mem_wdata[80]~66 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[80]~66 .shared_arith = "off";

dffeas \mem_wdata_r1[80] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[80]~66_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[80]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[80] .is_wysiwyg = "true";
defparam \mem_wdata_r1[80] .power_up = "low";

dffeas \mem_wdata_r2[80] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[80]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[80]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[80] .is_wysiwyg = "true";
defparam \mem_wdata_r2[80] .power_up = "low";

arriaii_lcell_comb \mem_wdata[16]~67 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_24),
	.datac(!q_b_16),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[16]~67_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[16]~67 .extended_lut = "off";
defparam \mem_wdata[16]~67 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[16]~67 .shared_arith = "off";

dffeas \mem_wdata_r1[16] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[16]~67_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[16]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[16] .is_wysiwyg = "true";
defparam \mem_wdata_r1[16] .power_up = "low";

dffeas \mem_wdata_r2[16] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[16]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[16]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[16] .is_wysiwyg = "true";
defparam \mem_wdata_r2[16] .power_up = "low";

dffeas \wdata_valid_1x_r1[12] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_valid[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r1[12]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r1[12] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r1[12] .power_up = "low";

dffeas \wdata_valid_1x_r2[12] (
	.clk(phy_clk_1x),
	.d(\wdata_valid_1x_r1[12]~q ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r2[12]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r2[12] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r2[12] .power_up = "low";

dffeas \wdata_valid_1x_r1[4] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_valid[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r1[4]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r1[4] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r1[4] .power_up = "low";

dffeas \wdata_valid_1x_r2[4] (
	.clk(phy_clk_1x),
	.d(\wdata_valid_1x_r1[4]~q ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r2[4]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r2[4] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r2[4] .power_up = "low";

arriaii_lcell_comb \mem_wdata[113]~68 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_121),
	.datac(!q_b_113),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[113]~68_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[113]~68 .extended_lut = "off";
defparam \mem_wdata[113]~68 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[113]~68 .shared_arith = "off";

dffeas \mem_wdata_r1[113] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[113]~68_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[113]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[113] .is_wysiwyg = "true";
defparam \mem_wdata_r1[113] .power_up = "low";

dffeas \mem_wdata_r2[113] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[113]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[113]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[113] .is_wysiwyg = "true";
defparam \mem_wdata_r2[113] .power_up = "low";

arriaii_lcell_comb \mem_wdata[49]~69 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_57),
	.datac(!q_b_49),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[49]~69_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[49]~69 .extended_lut = "off";
defparam \mem_wdata[49]~69 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[49]~69 .shared_arith = "off";

dffeas \mem_wdata_r1[49] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[49]~69_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[49]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[49] .is_wysiwyg = "true";
defparam \mem_wdata_r1[49] .power_up = "low";

dffeas \mem_wdata_r2[49] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[49]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[49]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[49] .is_wysiwyg = "true";
defparam \mem_wdata_r2[49] .power_up = "low";

arriaii_lcell_comb \mem_wdata[81]~70 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_89),
	.datac(!q_b_81),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[81]~70_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[81]~70 .extended_lut = "off";
defparam \mem_wdata[81]~70 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[81]~70 .shared_arith = "off";

dffeas \mem_wdata_r1[81] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[81]~70_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[81]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[81] .is_wysiwyg = "true";
defparam \mem_wdata_r1[81] .power_up = "low";

dffeas \mem_wdata_r2[81] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[81]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[81]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[81] .is_wysiwyg = "true";
defparam \mem_wdata_r2[81] .power_up = "low";

arriaii_lcell_comb \mem_wdata[17]~71 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_25),
	.datac(!q_b_17),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[17]~71_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[17]~71 .extended_lut = "off";
defparam \mem_wdata[17]~71 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[17]~71 .shared_arith = "off";

dffeas \mem_wdata_r1[17] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[17]~71_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[17]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[17] .is_wysiwyg = "true";
defparam \mem_wdata_r1[17] .power_up = "low";

dffeas \mem_wdata_r2[17] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[17]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[17]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[17] .is_wysiwyg = "true";
defparam \mem_wdata_r2[17] .power_up = "low";

arriaii_lcell_comb \mem_wdata[114]~72 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_122),
	.datac(!q_b_114),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[114]~72_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[114]~72 .extended_lut = "off";
defparam \mem_wdata[114]~72 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[114]~72 .shared_arith = "off";

dffeas \mem_wdata_r1[114] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[114]~72_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[114]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[114] .is_wysiwyg = "true";
defparam \mem_wdata_r1[114] .power_up = "low";

dffeas \mem_wdata_r2[114] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[114]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[114]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[114] .is_wysiwyg = "true";
defparam \mem_wdata_r2[114] .power_up = "low";

arriaii_lcell_comb \mem_wdata[50]~73 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_58),
	.datac(!q_b_50),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[50]~73_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[50]~73 .extended_lut = "off";
defparam \mem_wdata[50]~73 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[50]~73 .shared_arith = "off";

dffeas \mem_wdata_r1[50] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[50]~73_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[50]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[50] .is_wysiwyg = "true";
defparam \mem_wdata_r1[50] .power_up = "low";

dffeas \mem_wdata_r2[50] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[50]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[50]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[50] .is_wysiwyg = "true";
defparam \mem_wdata_r2[50] .power_up = "low";

arriaii_lcell_comb \mem_wdata[82]~74 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_90),
	.datac(!q_b_82),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[82]~74_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[82]~74 .extended_lut = "off";
defparam \mem_wdata[82]~74 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[82]~74 .shared_arith = "off";

dffeas \mem_wdata_r1[82] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[82]~74_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[82]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[82] .is_wysiwyg = "true";
defparam \mem_wdata_r1[82] .power_up = "low";

dffeas \mem_wdata_r2[82] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[82]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[82]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[82] .is_wysiwyg = "true";
defparam \mem_wdata_r2[82] .power_up = "low";

arriaii_lcell_comb \mem_wdata[18]~75 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_26),
	.datac(!q_b_18),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[18]~75_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[18]~75 .extended_lut = "off";
defparam \mem_wdata[18]~75 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[18]~75 .shared_arith = "off";

dffeas \mem_wdata_r1[18] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[18]~75_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[18]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[18] .is_wysiwyg = "true";
defparam \mem_wdata_r1[18] .power_up = "low";

dffeas \mem_wdata_r2[18] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[18]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[18]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[18] .is_wysiwyg = "true";
defparam \mem_wdata_r2[18] .power_up = "low";

arriaii_lcell_comb \mem_wdata[115]~76 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_123),
	.datac(!q_b_115),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[115]~76_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[115]~76 .extended_lut = "off";
defparam \mem_wdata[115]~76 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[115]~76 .shared_arith = "off";

dffeas \mem_wdata_r1[115] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[115]~76_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[115]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[115] .is_wysiwyg = "true";
defparam \mem_wdata_r1[115] .power_up = "low";

dffeas \mem_wdata_r2[115] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[115]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[115]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[115] .is_wysiwyg = "true";
defparam \mem_wdata_r2[115] .power_up = "low";

arriaii_lcell_comb \mem_wdata[51]~77 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_59),
	.datac(!q_b_51),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[51]~77_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[51]~77 .extended_lut = "off";
defparam \mem_wdata[51]~77 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[51]~77 .shared_arith = "off";

dffeas \mem_wdata_r1[51] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[51]~77_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[51]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[51] .is_wysiwyg = "true";
defparam \mem_wdata_r1[51] .power_up = "low";

dffeas \mem_wdata_r2[51] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[51]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[51]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[51] .is_wysiwyg = "true";
defparam \mem_wdata_r2[51] .power_up = "low";

arriaii_lcell_comb \mem_wdata[83]~78 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_91),
	.datac(!q_b_83),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[83]~78_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[83]~78 .extended_lut = "off";
defparam \mem_wdata[83]~78 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[83]~78 .shared_arith = "off";

dffeas \mem_wdata_r1[83] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[83]~78_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[83]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[83] .is_wysiwyg = "true";
defparam \mem_wdata_r1[83] .power_up = "low";

dffeas \mem_wdata_r2[83] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[83]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[83]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[83] .is_wysiwyg = "true";
defparam \mem_wdata_r2[83] .power_up = "low";

arriaii_lcell_comb \mem_wdata[19]~79 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_27),
	.datac(!q_b_19),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[19]~79_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[19]~79 .extended_lut = "off";
defparam \mem_wdata[19]~79 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[19]~79 .shared_arith = "off";

dffeas \mem_wdata_r1[19] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[19]~79_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[19]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[19] .is_wysiwyg = "true";
defparam \mem_wdata_r1[19] .power_up = "low";

dffeas \mem_wdata_r2[19] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[19]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[19]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[19] .is_wysiwyg = "true";
defparam \mem_wdata_r2[19] .power_up = "low";

arriaii_lcell_comb \mem_wdata[116]~80 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_124),
	.datac(!q_b_116),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[116]~80_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[116]~80 .extended_lut = "off";
defparam \mem_wdata[116]~80 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[116]~80 .shared_arith = "off";

dffeas \mem_wdata_r1[116] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[116]~80_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[116]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[116] .is_wysiwyg = "true";
defparam \mem_wdata_r1[116] .power_up = "low";

dffeas \mem_wdata_r2[116] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[116]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[116]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[116] .is_wysiwyg = "true";
defparam \mem_wdata_r2[116] .power_up = "low";

arriaii_lcell_comb \mem_wdata[52]~81 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_60),
	.datac(!q_b_52),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[52]~81_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[52]~81 .extended_lut = "off";
defparam \mem_wdata[52]~81 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[52]~81 .shared_arith = "off";

dffeas \mem_wdata_r1[52] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[52]~81_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[52]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[52] .is_wysiwyg = "true";
defparam \mem_wdata_r1[52] .power_up = "low";

dffeas \mem_wdata_r2[52] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[52]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[52]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[52] .is_wysiwyg = "true";
defparam \mem_wdata_r2[52] .power_up = "low";

dffeas \wdata_valid_1x_r[5] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_valid[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r[5]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r[5] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r[5] .power_up = "low";

dffeas \wdata_valid_2x_r1[5] (
	.clk(write_clk_2x),
	.d(\wdata_valid_1x_r[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_2x_r1[5]~q ),
	.prn(vcc));
defparam \wdata_valid_2x_r1[5] .is_wysiwyg = "true";
defparam \wdata_valid_2x_r1[5] .power_up = "low";

dffeas \wdata_valid_2x_r2[5] (
	.clk(write_clk_2x),
	.d(\wdata_valid_2x_r1[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_2x_r2[5]~q ),
	.prn(vcc));
defparam \wdata_valid_2x_r2[5] .is_wysiwyg = "true";
defparam \wdata_valid_2x_r2[5] .power_up = "low";

arriaii_lcell_comb \wdata_sel~5 (
	.dataa(!\wdata_sel[5]~q ),
	.datab(!\wdata_valid_2x_r2[5]~q ),
	.datac(!\wdata_valid_2x_r1[5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wdata_sel~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wdata_sel~5 .extended_lut = "off";
defparam \wdata_sel~5 .lut_mask = 64'hA2A2A2A2A2A2A2A2;
defparam \wdata_sel~5 .shared_arith = "off";

dffeas \wdata_sel[5] (
	.clk(write_clk_2x),
	.d(\wdata_sel~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_sel[5]~q ),
	.prn(vcc));
defparam \wdata_sel[5] .is_wysiwyg = "true";
defparam \wdata_sel[5] .power_up = "low";

arriaii_lcell_comb \mem_wdata[84]~82 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_92),
	.datac(!q_b_84),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[84]~82_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[84]~82 .extended_lut = "off";
defparam \mem_wdata[84]~82 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[84]~82 .shared_arith = "off";

dffeas \mem_wdata_r1[84] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[84]~82_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[84]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[84] .is_wysiwyg = "true";
defparam \mem_wdata_r1[84] .power_up = "low";

dffeas \mem_wdata_r2[84] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[84]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[84]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[84] .is_wysiwyg = "true";
defparam \mem_wdata_r2[84] .power_up = "low";

arriaii_lcell_comb \mem_wdata[20]~83 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_28),
	.datac(!q_b_20),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[20]~83_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[20]~83 .extended_lut = "off";
defparam \mem_wdata[20]~83 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[20]~83 .shared_arith = "off";

dffeas \mem_wdata_r1[20] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[20]~83_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[20]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[20] .is_wysiwyg = "true";
defparam \mem_wdata_r1[20] .power_up = "low";

dffeas \mem_wdata_r2[20] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[20]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[20]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[20] .is_wysiwyg = "true";
defparam \mem_wdata_r2[20] .power_up = "low";

dffeas \wdata_valid_1x_r1[13] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_valid[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r1[13]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r1[13] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r1[13] .power_up = "low";

dffeas \wdata_valid_1x_r2[13] (
	.clk(phy_clk_1x),
	.d(\wdata_valid_1x_r1[13]~q ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r2[13]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r2[13] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r2[13] .power_up = "low";

dffeas \wdata_valid_1x_r1[5] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_valid[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r1[5]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r1[5] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r1[5] .power_up = "low";

dffeas \wdata_valid_1x_r2[5] (
	.clk(phy_clk_1x),
	.d(\wdata_valid_1x_r1[5]~q ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r2[5]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r2[5] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r2[5] .power_up = "low";

arriaii_lcell_comb \mem_wdata[117]~84 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_125),
	.datac(!q_b_117),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[117]~84_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[117]~84 .extended_lut = "off";
defparam \mem_wdata[117]~84 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[117]~84 .shared_arith = "off";

dffeas \mem_wdata_r1[117] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[117]~84_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[117]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[117] .is_wysiwyg = "true";
defparam \mem_wdata_r1[117] .power_up = "low";

dffeas \mem_wdata_r2[117] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[117]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[117]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[117] .is_wysiwyg = "true";
defparam \mem_wdata_r2[117] .power_up = "low";

arriaii_lcell_comb \mem_wdata[53]~85 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_61),
	.datac(!q_b_53),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[53]~85_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[53]~85 .extended_lut = "off";
defparam \mem_wdata[53]~85 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[53]~85 .shared_arith = "off";

dffeas \mem_wdata_r1[53] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[53]~85_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[53]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[53] .is_wysiwyg = "true";
defparam \mem_wdata_r1[53] .power_up = "low";

dffeas \mem_wdata_r2[53] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[53]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[53]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[53] .is_wysiwyg = "true";
defparam \mem_wdata_r2[53] .power_up = "low";

arriaii_lcell_comb \mem_wdata[85]~86 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_93),
	.datac(!q_b_85),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[85]~86_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[85]~86 .extended_lut = "off";
defparam \mem_wdata[85]~86 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[85]~86 .shared_arith = "off";

dffeas \mem_wdata_r1[85] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[85]~86_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[85]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[85] .is_wysiwyg = "true";
defparam \mem_wdata_r1[85] .power_up = "low";

dffeas \mem_wdata_r2[85] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[85]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[85]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[85] .is_wysiwyg = "true";
defparam \mem_wdata_r2[85] .power_up = "low";

arriaii_lcell_comb \mem_wdata[21]~87 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_29),
	.datac(!q_b_21),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[21]~87_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[21]~87 .extended_lut = "off";
defparam \mem_wdata[21]~87 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[21]~87 .shared_arith = "off";

dffeas \mem_wdata_r1[21] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[21]~87_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[21]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[21] .is_wysiwyg = "true";
defparam \mem_wdata_r1[21] .power_up = "low";

dffeas \mem_wdata_r2[21] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[21]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[21]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[21] .is_wysiwyg = "true";
defparam \mem_wdata_r2[21] .power_up = "low";

arriaii_lcell_comb \mem_wdata[118]~88 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_126),
	.datac(!q_b_118),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[118]~88_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[118]~88 .extended_lut = "off";
defparam \mem_wdata[118]~88 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[118]~88 .shared_arith = "off";

dffeas \mem_wdata_r1[118] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[118]~88_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[118]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[118] .is_wysiwyg = "true";
defparam \mem_wdata_r1[118] .power_up = "low";

dffeas \mem_wdata_r2[118] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[118]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[118]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[118] .is_wysiwyg = "true";
defparam \mem_wdata_r2[118] .power_up = "low";

arriaii_lcell_comb \mem_wdata[54]~89 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_62),
	.datac(!q_b_54),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[54]~89_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[54]~89 .extended_lut = "off";
defparam \mem_wdata[54]~89 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[54]~89 .shared_arith = "off";

dffeas \mem_wdata_r1[54] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[54]~89_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[54]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[54] .is_wysiwyg = "true";
defparam \mem_wdata_r1[54] .power_up = "low";

dffeas \mem_wdata_r2[54] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[54]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[54]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[54] .is_wysiwyg = "true";
defparam \mem_wdata_r2[54] .power_up = "low";

arriaii_lcell_comb \mem_wdata[86]~90 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_94),
	.datac(!q_b_86),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[86]~90_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[86]~90 .extended_lut = "off";
defparam \mem_wdata[86]~90 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[86]~90 .shared_arith = "off";

dffeas \mem_wdata_r1[86] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[86]~90_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[86]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[86] .is_wysiwyg = "true";
defparam \mem_wdata_r1[86] .power_up = "low";

dffeas \mem_wdata_r2[86] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[86]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[86]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[86] .is_wysiwyg = "true";
defparam \mem_wdata_r2[86] .power_up = "low";

arriaii_lcell_comb \mem_wdata[22]~91 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_30),
	.datac(!q_b_22),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[22]~91_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[22]~91 .extended_lut = "off";
defparam \mem_wdata[22]~91 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[22]~91 .shared_arith = "off";

dffeas \mem_wdata_r1[22] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[22]~91_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[22]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[22] .is_wysiwyg = "true";
defparam \mem_wdata_r1[22] .power_up = "low";

dffeas \mem_wdata_r2[22] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[22]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[22]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[22] .is_wysiwyg = "true";
defparam \mem_wdata_r2[22] .power_up = "low";

arriaii_lcell_comb \mem_wdata[119]~92 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_127),
	.datac(!q_b_119),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[119]~92_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[119]~92 .extended_lut = "off";
defparam \mem_wdata[119]~92 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[119]~92 .shared_arith = "off";

dffeas \mem_wdata_r1[119] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[119]~92_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[119]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[119] .is_wysiwyg = "true";
defparam \mem_wdata_r1[119] .power_up = "low";

dffeas \mem_wdata_r2[119] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[119]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[119]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[119] .is_wysiwyg = "true";
defparam \mem_wdata_r2[119] .power_up = "low";

arriaii_lcell_comb \mem_wdata[55]~93 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_63),
	.datac(!q_b_55),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[55]~93_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[55]~93 .extended_lut = "off";
defparam \mem_wdata[55]~93 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[55]~93 .shared_arith = "off";

dffeas \mem_wdata_r1[55] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[55]~93_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[55]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[55] .is_wysiwyg = "true";
defparam \mem_wdata_r1[55] .power_up = "low";

dffeas \mem_wdata_r2[55] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[55]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[55]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[55] .is_wysiwyg = "true";
defparam \mem_wdata_r2[55] .power_up = "low";

arriaii_lcell_comb \mem_wdata[87]~94 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_95),
	.datac(!q_b_87),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[87]~94_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[87]~94 .extended_lut = "off";
defparam \mem_wdata[87]~94 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[87]~94 .shared_arith = "off";

dffeas \mem_wdata_r1[87] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[87]~94_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[87]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[87] .is_wysiwyg = "true";
defparam \mem_wdata_r1[87] .power_up = "low";

dffeas \mem_wdata_r2[87] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[87]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[87]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[87] .is_wysiwyg = "true";
defparam \mem_wdata_r2[87] .power_up = "low";

arriaii_lcell_comb \mem_wdata[23]~95 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_31),
	.datac(!q_b_23),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[23]~95_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[23]~95 .extended_lut = "off";
defparam \mem_wdata[23]~95 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[23]~95 .shared_arith = "off";

dffeas \mem_wdata_r1[23] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[23]~95_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[23]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[23] .is_wysiwyg = "true";
defparam \mem_wdata_r1[23] .power_up = "low";

dffeas \mem_wdata_r2[23] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[23]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[23]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[23] .is_wysiwyg = "true";
defparam \mem_wdata_r2[23] .power_up = "low";

arriaii_lcell_comb \mem_wdata[120]~96 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_120),
	.datac(!q_b_120),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[120]~96_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[120]~96 .extended_lut = "off";
defparam \mem_wdata[120]~96 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[120]~96 .shared_arith = "off";

dffeas \mem_wdata_r1[120] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[120]~96_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[120]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[120] .is_wysiwyg = "true";
defparam \mem_wdata_r1[120] .power_up = "low";

dffeas \mem_wdata_r2[120] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[120]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[120]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[120] .is_wysiwyg = "true";
defparam \mem_wdata_r2[120] .power_up = "low";

arriaii_lcell_comb \mem_wdata[56]~97 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_56),
	.datac(!q_b_56),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[56]~97_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[56]~97 .extended_lut = "off";
defparam \mem_wdata[56]~97 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[56]~97 .shared_arith = "off";

dffeas \mem_wdata_r1[56] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[56]~97_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[56]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[56] .is_wysiwyg = "true";
defparam \mem_wdata_r1[56] .power_up = "low";

dffeas \mem_wdata_r2[56] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[56]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[56]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[56] .is_wysiwyg = "true";
defparam \mem_wdata_r2[56] .power_up = "low";

dffeas \wdata_valid_1x_r[6] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_valid[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r[6]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r[6] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r[6] .power_up = "low";

dffeas \wdata_valid_2x_r1[6] (
	.clk(write_clk_2x),
	.d(\wdata_valid_1x_r[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_2x_r1[6]~q ),
	.prn(vcc));
defparam \wdata_valid_2x_r1[6] .is_wysiwyg = "true";
defparam \wdata_valid_2x_r1[6] .power_up = "low";

dffeas \wdata_valid_2x_r2[6] (
	.clk(write_clk_2x),
	.d(\wdata_valid_2x_r1[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_2x_r2[6]~q ),
	.prn(vcc));
defparam \wdata_valid_2x_r2[6] .is_wysiwyg = "true";
defparam \wdata_valid_2x_r2[6] .power_up = "low";

arriaii_lcell_comb \wdata_sel~6 (
	.dataa(!\wdata_sel[6]~q ),
	.datab(!\wdata_valid_2x_r2[6]~q ),
	.datac(!\wdata_valid_2x_r1[6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wdata_sel~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wdata_sel~6 .extended_lut = "off";
defparam \wdata_sel~6 .lut_mask = 64'hA2A2A2A2A2A2A2A2;
defparam \wdata_sel~6 .shared_arith = "off";

dffeas \wdata_sel[6] (
	.clk(write_clk_2x),
	.d(\wdata_sel~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_sel[6]~q ),
	.prn(vcc));
defparam \wdata_sel[6] .is_wysiwyg = "true";
defparam \wdata_sel[6] .power_up = "low";

arriaii_lcell_comb \mem_wdata[88]~98 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_88),
	.datac(!q_b_88),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[88]~98_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[88]~98 .extended_lut = "off";
defparam \mem_wdata[88]~98 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[88]~98 .shared_arith = "off";

dffeas \mem_wdata_r1[88] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[88]~98_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[88]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[88] .is_wysiwyg = "true";
defparam \mem_wdata_r1[88] .power_up = "low";

dffeas \mem_wdata_r2[88] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[88]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[88]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[88] .is_wysiwyg = "true";
defparam \mem_wdata_r2[88] .power_up = "low";

arriaii_lcell_comb \mem_wdata[24]~99 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_24),
	.datac(!q_b_24),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[24]~99_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[24]~99 .extended_lut = "off";
defparam \mem_wdata[24]~99 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[24]~99 .shared_arith = "off";

dffeas \mem_wdata_r1[24] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[24]~99_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[24]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[24] .is_wysiwyg = "true";
defparam \mem_wdata_r1[24] .power_up = "low";

dffeas \mem_wdata_r2[24] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[24]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[24]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[24] .is_wysiwyg = "true";
defparam \mem_wdata_r2[24] .power_up = "low";

dffeas \wdata_valid_1x_r1[14] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_valid[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r1[14]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r1[14] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r1[14] .power_up = "low";

dffeas \wdata_valid_1x_r2[14] (
	.clk(phy_clk_1x),
	.d(\wdata_valid_1x_r1[14]~q ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r2[14]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r2[14] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r2[14] .power_up = "low";

dffeas \wdata_valid_1x_r1[6] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_valid[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r1[6]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r1[6] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r1[6] .power_up = "low";

dffeas \wdata_valid_1x_r2[6] (
	.clk(phy_clk_1x),
	.d(\wdata_valid_1x_r1[6]~q ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r2[6]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r2[6] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r2[6] .power_up = "low";

arriaii_lcell_comb \mem_wdata[121]~100 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_121),
	.datac(!q_b_121),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[121]~100_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[121]~100 .extended_lut = "off";
defparam \mem_wdata[121]~100 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[121]~100 .shared_arith = "off";

dffeas \mem_wdata_r1[121] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[121]~100_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[121]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[121] .is_wysiwyg = "true";
defparam \mem_wdata_r1[121] .power_up = "low";

dffeas \mem_wdata_r2[121] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[121]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[121]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[121] .is_wysiwyg = "true";
defparam \mem_wdata_r2[121] .power_up = "low";

arriaii_lcell_comb \mem_wdata[57]~101 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_57),
	.datac(!q_b_57),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[57]~101_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[57]~101 .extended_lut = "off";
defparam \mem_wdata[57]~101 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[57]~101 .shared_arith = "off";

dffeas \mem_wdata_r1[57] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[57]~101_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[57]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[57] .is_wysiwyg = "true";
defparam \mem_wdata_r1[57] .power_up = "low";

dffeas \mem_wdata_r2[57] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[57]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[57]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[57] .is_wysiwyg = "true";
defparam \mem_wdata_r2[57] .power_up = "low";

arriaii_lcell_comb \mem_wdata[89]~102 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_89),
	.datac(!q_b_89),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[89]~102_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[89]~102 .extended_lut = "off";
defparam \mem_wdata[89]~102 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[89]~102 .shared_arith = "off";

dffeas \mem_wdata_r1[89] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[89]~102_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[89]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[89] .is_wysiwyg = "true";
defparam \mem_wdata_r1[89] .power_up = "low";

dffeas \mem_wdata_r2[89] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[89]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[89]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[89] .is_wysiwyg = "true";
defparam \mem_wdata_r2[89] .power_up = "low";

arriaii_lcell_comb \mem_wdata[25]~103 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_25),
	.datac(!q_b_25),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[25]~103_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[25]~103 .extended_lut = "off";
defparam \mem_wdata[25]~103 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[25]~103 .shared_arith = "off";

dffeas \mem_wdata_r1[25] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[25]~103_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[25]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[25] .is_wysiwyg = "true";
defparam \mem_wdata_r1[25] .power_up = "low";

dffeas \mem_wdata_r2[25] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[25]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[25]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[25] .is_wysiwyg = "true";
defparam \mem_wdata_r2[25] .power_up = "low";

arriaii_lcell_comb \mem_wdata[122]~104 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_122),
	.datac(!q_b_122),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[122]~104_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[122]~104 .extended_lut = "off";
defparam \mem_wdata[122]~104 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[122]~104 .shared_arith = "off";

dffeas \mem_wdata_r1[122] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[122]~104_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[122]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[122] .is_wysiwyg = "true";
defparam \mem_wdata_r1[122] .power_up = "low";

dffeas \mem_wdata_r2[122] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[122]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[122]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[122] .is_wysiwyg = "true";
defparam \mem_wdata_r2[122] .power_up = "low";

arriaii_lcell_comb \mem_wdata[58]~105 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_58),
	.datac(!q_b_58),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[58]~105_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[58]~105 .extended_lut = "off";
defparam \mem_wdata[58]~105 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[58]~105 .shared_arith = "off";

dffeas \mem_wdata_r1[58] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[58]~105_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[58]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[58] .is_wysiwyg = "true";
defparam \mem_wdata_r1[58] .power_up = "low";

dffeas \mem_wdata_r2[58] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[58]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[58]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[58] .is_wysiwyg = "true";
defparam \mem_wdata_r2[58] .power_up = "low";

arriaii_lcell_comb \mem_wdata[90]~106 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_90),
	.datac(!q_b_90),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[90]~106_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[90]~106 .extended_lut = "off";
defparam \mem_wdata[90]~106 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[90]~106 .shared_arith = "off";

dffeas \mem_wdata_r1[90] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[90]~106_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[90]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[90] .is_wysiwyg = "true";
defparam \mem_wdata_r1[90] .power_up = "low";

dffeas \mem_wdata_r2[90] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[90]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[90]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[90] .is_wysiwyg = "true";
defparam \mem_wdata_r2[90] .power_up = "low";

arriaii_lcell_comb \mem_wdata[26]~107 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_26),
	.datac(!q_b_26),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[26]~107_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[26]~107 .extended_lut = "off";
defparam \mem_wdata[26]~107 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[26]~107 .shared_arith = "off";

dffeas \mem_wdata_r1[26] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[26]~107_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[26]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[26] .is_wysiwyg = "true";
defparam \mem_wdata_r1[26] .power_up = "low";

dffeas \mem_wdata_r2[26] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[26]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[26]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[26] .is_wysiwyg = "true";
defparam \mem_wdata_r2[26] .power_up = "low";

arriaii_lcell_comb \mem_wdata[123]~108 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_123),
	.datac(!q_b_123),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[123]~108_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[123]~108 .extended_lut = "off";
defparam \mem_wdata[123]~108 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[123]~108 .shared_arith = "off";

dffeas \mem_wdata_r1[123] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[123]~108_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[123]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[123] .is_wysiwyg = "true";
defparam \mem_wdata_r1[123] .power_up = "low";

dffeas \mem_wdata_r2[123] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[123]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[123]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[123] .is_wysiwyg = "true";
defparam \mem_wdata_r2[123] .power_up = "low";

arriaii_lcell_comb \mem_wdata[59]~109 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_59),
	.datac(!q_b_59),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[59]~109_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[59]~109 .extended_lut = "off";
defparam \mem_wdata[59]~109 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[59]~109 .shared_arith = "off";

dffeas \mem_wdata_r1[59] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[59]~109_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[59]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[59] .is_wysiwyg = "true";
defparam \mem_wdata_r1[59] .power_up = "low";

dffeas \mem_wdata_r2[59] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[59]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[59]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[59] .is_wysiwyg = "true";
defparam \mem_wdata_r2[59] .power_up = "low";

arriaii_lcell_comb \mem_wdata[91]~110 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_91),
	.datac(!q_b_91),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[91]~110_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[91]~110 .extended_lut = "off";
defparam \mem_wdata[91]~110 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[91]~110 .shared_arith = "off";

dffeas \mem_wdata_r1[91] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[91]~110_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[91]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[91] .is_wysiwyg = "true";
defparam \mem_wdata_r1[91] .power_up = "low";

dffeas \mem_wdata_r2[91] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[91]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[91]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[91] .is_wysiwyg = "true";
defparam \mem_wdata_r2[91] .power_up = "low";

arriaii_lcell_comb \mem_wdata[27]~111 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_27),
	.datac(!q_b_27),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[27]~111_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[27]~111 .extended_lut = "off";
defparam \mem_wdata[27]~111 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[27]~111 .shared_arith = "off";

dffeas \mem_wdata_r1[27] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[27]~111_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[27]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[27] .is_wysiwyg = "true";
defparam \mem_wdata_r1[27] .power_up = "low";

dffeas \mem_wdata_r2[27] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[27]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[27]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[27] .is_wysiwyg = "true";
defparam \mem_wdata_r2[27] .power_up = "low";

arriaii_lcell_comb \mem_wdata[124]~112 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_124),
	.datac(!q_b_124),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[124]~112_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[124]~112 .extended_lut = "off";
defparam \mem_wdata[124]~112 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[124]~112 .shared_arith = "off";

dffeas \mem_wdata_r1[124] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[124]~112_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[124]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[124] .is_wysiwyg = "true";
defparam \mem_wdata_r1[124] .power_up = "low";

dffeas \mem_wdata_r2[124] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[124]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[124]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[124] .is_wysiwyg = "true";
defparam \mem_wdata_r2[124] .power_up = "low";

arriaii_lcell_comb \mem_wdata[60]~113 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_60),
	.datac(!q_b_60),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[60]~113_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[60]~113 .extended_lut = "off";
defparam \mem_wdata[60]~113 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[60]~113 .shared_arith = "off";

dffeas \mem_wdata_r1[60] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[60]~113_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[60]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[60] .is_wysiwyg = "true";
defparam \mem_wdata_r1[60] .power_up = "low";

dffeas \mem_wdata_r2[60] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[60]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[60]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[60] .is_wysiwyg = "true";
defparam \mem_wdata_r2[60] .power_up = "low";

dffeas \wdata_valid_1x_r[7] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_valid[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r[7]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r[7] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r[7] .power_up = "low";

dffeas \wdata_valid_2x_r1[7] (
	.clk(write_clk_2x),
	.d(\wdata_valid_1x_r[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_2x_r1[7]~q ),
	.prn(vcc));
defparam \wdata_valid_2x_r1[7] .is_wysiwyg = "true";
defparam \wdata_valid_2x_r1[7] .power_up = "low";

dffeas \wdata_valid_2x_r2[7] (
	.clk(write_clk_2x),
	.d(\wdata_valid_2x_r1[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_2x_r2[7]~q ),
	.prn(vcc));
defparam \wdata_valid_2x_r2[7] .is_wysiwyg = "true";
defparam \wdata_valid_2x_r2[7] .power_up = "low";

arriaii_lcell_comb \wdata_sel~7 (
	.dataa(!\wdata_sel[7]~q ),
	.datab(!\wdata_valid_2x_r2[7]~q ),
	.datac(!\wdata_valid_2x_r1[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wdata_sel~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wdata_sel~7 .extended_lut = "off";
defparam \wdata_sel~7 .lut_mask = 64'hA2A2A2A2A2A2A2A2;
defparam \wdata_sel~7 .shared_arith = "off";

dffeas \wdata_sel[7] (
	.clk(write_clk_2x),
	.d(\wdata_sel~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_sel[7]~q ),
	.prn(vcc));
defparam \wdata_sel[7] .is_wysiwyg = "true";
defparam \wdata_sel[7] .power_up = "low";

arriaii_lcell_comb \mem_wdata[92]~114 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_92),
	.datac(!q_b_92),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[92]~114_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[92]~114 .extended_lut = "off";
defparam \mem_wdata[92]~114 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[92]~114 .shared_arith = "off";

dffeas \mem_wdata_r1[92] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[92]~114_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[92]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[92] .is_wysiwyg = "true";
defparam \mem_wdata_r1[92] .power_up = "low";

dffeas \mem_wdata_r2[92] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[92]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[92]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[92] .is_wysiwyg = "true";
defparam \mem_wdata_r2[92] .power_up = "low";

arriaii_lcell_comb \mem_wdata[28]~115 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_28),
	.datac(!q_b_28),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[28]~115_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[28]~115 .extended_lut = "off";
defparam \mem_wdata[28]~115 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[28]~115 .shared_arith = "off";

dffeas \mem_wdata_r1[28] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[28]~115_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[28]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[28] .is_wysiwyg = "true";
defparam \mem_wdata_r1[28] .power_up = "low";

dffeas \mem_wdata_r2[28] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[28]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[28]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[28] .is_wysiwyg = "true";
defparam \mem_wdata_r2[28] .power_up = "low";

dffeas \wdata_valid_1x_r1[15] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_valid[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r1[15]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r1[15] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r1[15] .power_up = "low";

dffeas \wdata_valid_1x_r2[15] (
	.clk(phy_clk_1x),
	.d(\wdata_valid_1x_r1[15]~q ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r2[15]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r2[15] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r2[15] .power_up = "low";

dffeas \wdata_valid_1x_r1[7] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_valid[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r1[7]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r1[7] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r1[7] .power_up = "low";

dffeas \wdata_valid_1x_r2[7] (
	.clk(phy_clk_1x),
	.d(\wdata_valid_1x_r1[7]~q ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wdata_valid_1x_r2[7]~q ),
	.prn(vcc));
defparam \wdata_valid_1x_r2[7] .is_wysiwyg = "true";
defparam \wdata_valid_1x_r2[7] .power_up = "low";

arriaii_lcell_comb \mem_wdata[125]~116 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_125),
	.datac(!q_b_125),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[125]~116_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[125]~116 .extended_lut = "off";
defparam \mem_wdata[125]~116 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[125]~116 .shared_arith = "off";

dffeas \mem_wdata_r1[125] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[125]~116_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[125]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[125] .is_wysiwyg = "true";
defparam \mem_wdata_r1[125] .power_up = "low";

dffeas \mem_wdata_r2[125] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[125]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[125]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[125] .is_wysiwyg = "true";
defparam \mem_wdata_r2[125] .power_up = "low";

arriaii_lcell_comb \mem_wdata[61]~117 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_61),
	.datac(!q_b_61),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[61]~117_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[61]~117 .extended_lut = "off";
defparam \mem_wdata[61]~117 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[61]~117 .shared_arith = "off";

dffeas \mem_wdata_r1[61] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[61]~117_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[61]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[61] .is_wysiwyg = "true";
defparam \mem_wdata_r1[61] .power_up = "low";

dffeas \mem_wdata_r2[61] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[61]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[61]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[61] .is_wysiwyg = "true";
defparam \mem_wdata_r2[61] .power_up = "low";

arriaii_lcell_comb \mem_wdata[93]~118 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_93),
	.datac(!q_b_93),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[93]~118_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[93]~118 .extended_lut = "off";
defparam \mem_wdata[93]~118 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[93]~118 .shared_arith = "off";

dffeas \mem_wdata_r1[93] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[93]~118_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[93]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[93] .is_wysiwyg = "true";
defparam \mem_wdata_r1[93] .power_up = "low";

dffeas \mem_wdata_r2[93] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[93]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[93]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[93] .is_wysiwyg = "true";
defparam \mem_wdata_r2[93] .power_up = "low";

arriaii_lcell_comb \mem_wdata[29]~119 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_29),
	.datac(!q_b_29),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[29]~119_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[29]~119 .extended_lut = "off";
defparam \mem_wdata[29]~119 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[29]~119 .shared_arith = "off";

dffeas \mem_wdata_r1[29] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[29]~119_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[29]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[29] .is_wysiwyg = "true";
defparam \mem_wdata_r1[29] .power_up = "low";

dffeas \mem_wdata_r2[29] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[29]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[29]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[29] .is_wysiwyg = "true";
defparam \mem_wdata_r2[29] .power_up = "low";

arriaii_lcell_comb \mem_wdata[126]~120 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_126),
	.datac(!q_b_126),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[126]~120_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[126]~120 .extended_lut = "off";
defparam \mem_wdata[126]~120 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[126]~120 .shared_arith = "off";

dffeas \mem_wdata_r1[126] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[126]~120_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[126]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[126] .is_wysiwyg = "true";
defparam \mem_wdata_r1[126] .power_up = "low";

dffeas \mem_wdata_r2[126] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[126]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[126]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[126] .is_wysiwyg = "true";
defparam \mem_wdata_r2[126] .power_up = "low";

arriaii_lcell_comb \mem_wdata[62]~121 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_62),
	.datac(!q_b_62),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[62]~121_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[62]~121 .extended_lut = "off";
defparam \mem_wdata[62]~121 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[62]~121 .shared_arith = "off";

dffeas \mem_wdata_r1[62] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[62]~121_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[62]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[62] .is_wysiwyg = "true";
defparam \mem_wdata_r1[62] .power_up = "low";

dffeas \mem_wdata_r2[62] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[62]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[62]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[62] .is_wysiwyg = "true";
defparam \mem_wdata_r2[62] .power_up = "low";

arriaii_lcell_comb \mem_wdata[94]~122 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_94),
	.datac(!q_b_94),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[94]~122_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[94]~122 .extended_lut = "off";
defparam \mem_wdata[94]~122 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[94]~122 .shared_arith = "off";

dffeas \mem_wdata_r1[94] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[94]~122_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[94]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[94] .is_wysiwyg = "true";
defparam \mem_wdata_r1[94] .power_up = "low";

dffeas \mem_wdata_r2[94] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[94]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[94]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[94] .is_wysiwyg = "true";
defparam \mem_wdata_r2[94] .power_up = "low";

arriaii_lcell_comb \mem_wdata[30]~123 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_30),
	.datac(!q_b_30),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[30]~123_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[30]~123 .extended_lut = "off";
defparam \mem_wdata[30]~123 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[30]~123 .shared_arith = "off";

dffeas \mem_wdata_r1[30] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[30]~123_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[30]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[30] .is_wysiwyg = "true";
defparam \mem_wdata_r1[30] .power_up = "low";

dffeas \mem_wdata_r2[30] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[30]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[30]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[30] .is_wysiwyg = "true";
defparam \mem_wdata_r2[30] .power_up = "low";

arriaii_lcell_comb \mem_wdata[127]~124 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_127),
	.datac(!q_b_127),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[127]~124_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[127]~124 .extended_lut = "off";
defparam \mem_wdata[127]~124 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[127]~124 .shared_arith = "off";

dffeas \mem_wdata_r1[127] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[127]~124_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[127]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[127] .is_wysiwyg = "true";
defparam \mem_wdata_r1[127] .power_up = "low";

dffeas \mem_wdata_r2[127] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[127]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[127]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[127] .is_wysiwyg = "true";
defparam \mem_wdata_r2[127] .power_up = "low";

arriaii_lcell_comb \mem_wdata[63]~125 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_63),
	.datac(!q_b_63),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[63]~125_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[63]~125 .extended_lut = "off";
defparam \mem_wdata[63]~125 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[63]~125 .shared_arith = "off";

dffeas \mem_wdata_r1[63] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[63]~125_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[63]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[63] .is_wysiwyg = "true";
defparam \mem_wdata_r1[63] .power_up = "low";

dffeas \mem_wdata_r2[63] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[63]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[63]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[63] .is_wysiwyg = "true";
defparam \mem_wdata_r2[63] .power_up = "low";

arriaii_lcell_comb \mem_wdata[95]~126 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_95),
	.datac(!q_b_95),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[95]~126_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[95]~126 .extended_lut = "off";
defparam \mem_wdata[95]~126 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[95]~126 .shared_arith = "off";

dffeas \mem_wdata_r1[95] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[95]~126_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[95]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[95] .is_wysiwyg = "true";
defparam \mem_wdata_r1[95] .power_up = "low";

dffeas \mem_wdata_r2[95] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[95]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[95]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[95] .is_wysiwyg = "true";
defparam \mem_wdata_r2[95] .power_up = "low";

arriaii_lcell_comb \mem_wdata[31]~127 (
	.dataa(!seq_wdp_ovride),
	.datab(!dgwb_wdata_31),
	.datac(!q_b_31),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_wdata[31]~127_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_wdata[31]~127 .extended_lut = "off";
defparam \mem_wdata[31]~127 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \mem_wdata[31]~127 .shared_arith = "off";

dffeas \mem_wdata_r1[31] (
	.clk(phy_clk_1x),
	.d(\mem_wdata[31]~127_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r1[31]~q ),
	.prn(vcc));
defparam \mem_wdata_r1[31] .is_wysiwyg = "true";
defparam \mem_wdata_r1[31] .power_up = "low";

dffeas \mem_wdata_r2[31] (
	.clk(phy_clk_1x),
	.d(\mem_wdata_r1[31]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_wdata_r2[31]~q ),
	.prn(vcc));
defparam \mem_wdata_r2[31] .is_wysiwyg = "true";
defparam \mem_wdata_r2[31] .power_up = "low";

arriaii_lcell_comb \mem_dqs_burst[4]~0 (
	.dataa(!ctl_init_fail),
	.datab(!ctl_init_success),
	.datac(!dgwb_wdp_ovride),
	.datad(!int_dqs_burst),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_dqs_burst[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_dqs_burst[4]~0 .extended_lut = "off";
defparam \mem_dqs_burst[4]~0 .lut_mask = 64'h08FF08FF08FF08FF;
defparam \mem_dqs_burst[4]~0 .shared_arith = "off";

dffeas \dqs_burst_1x_r[4] (
	.clk(phy_clk_1x),
	.d(\mem_dqs_burst[4]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst_1x_r[4]~q ),
	.prn(vcc));
defparam \dqs_burst_1x_r[4] .is_wysiwyg = "true";
defparam \dqs_burst_1x_r[4] .power_up = "low";

dffeas \dqs_burst_2x_r1[4] (
	.clk(mem_clk_2x),
	.d(\dqs_burst_1x_r[4]~q ),
	.asdata(vcc),
	.clrn(reset_mem_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst_2x_r1[4]~q ),
	.prn(vcc));
defparam \dqs_burst_2x_r1[4] .is_wysiwyg = "true";
defparam \dqs_burst_2x_r1[4] .power_up = "low";

arriaii_lcell_comb \mem_dqs_burst[0]~1 (
	.dataa(!ctl_init_fail),
	.datab(!ctl_init_success),
	.datac(!dgwb_wdp_ovride),
	.datad(!int_dqs_burst_hr),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_dqs_burst[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_dqs_burst[0]~1 .extended_lut = "off";
defparam \mem_dqs_burst[0]~1 .lut_mask = 64'h08FF08FF08FF08FF;
defparam \mem_dqs_burst[0]~1 .shared_arith = "off";

dffeas \dqs_burst_1x_r[0] (
	.clk(phy_clk_1x),
	.d(\mem_dqs_burst[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst_1x_r[0]~q ),
	.prn(vcc));
defparam \dqs_burst_1x_r[0] .is_wysiwyg = "true";
defparam \dqs_burst_1x_r[0] .power_up = "low";

dffeas \dqs_burst_2x_r1[0] (
	.clk(mem_clk_2x),
	.d(\dqs_burst_1x_r[0]~q ),
	.asdata(vcc),
	.clrn(reset_mem_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst_2x_r1[0]~q ),
	.prn(vcc));
defparam \dqs_burst_2x_r1[0] .is_wysiwyg = "true";
defparam \dqs_burst_2x_r1[0] .power_up = "low";

arriaii_lcell_comb \dqs_burst_2x_r2~0 (
	.dataa(!\dqs_burst_sel[0]~q ),
	.datab(!\dqs_burst_2x_r1[4]~q ),
	.datac(!\dqs_burst_2x_r1[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dqs_burst_2x_r2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dqs_burst_2x_r2~0 .extended_lut = "off";
defparam \dqs_burst_2x_r2~0 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \dqs_burst_2x_r2~0 .shared_arith = "off";

dffeas \dqs_burst_2x_r2[0] (
	.clk(mem_clk_2x),
	.d(\dqs_burst_2x_r2~0_combout ),
	.asdata(vcc),
	.clrn(reset_mem_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst_2x_r2[0]~q ),
	.prn(vcc));
defparam \dqs_burst_2x_r2[0] .is_wysiwyg = "true";
defparam \dqs_burst_2x_r2[0] .power_up = "low";

dffeas \dqs_burst_1x_r[5] (
	.clk(phy_clk_1x),
	.d(\mem_dqs_burst[4]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst_1x_r[5]~q ),
	.prn(vcc));
defparam \dqs_burst_1x_r[5] .is_wysiwyg = "true";
defparam \dqs_burst_1x_r[5] .power_up = "low";

dffeas \dqs_burst_2x_r1[5] (
	.clk(mem_clk_2x),
	.d(\dqs_burst_1x_r[5]~q ),
	.asdata(vcc),
	.clrn(reset_mem_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst_2x_r1[5]~q ),
	.prn(vcc));
defparam \dqs_burst_2x_r1[5] .is_wysiwyg = "true";
defparam \dqs_burst_2x_r1[5] .power_up = "low";

dffeas \dqs_burst_1x_r[1] (
	.clk(phy_clk_1x),
	.d(\mem_dqs_burst[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst_1x_r[1]~q ),
	.prn(vcc));
defparam \dqs_burst_1x_r[1] .is_wysiwyg = "true";
defparam \dqs_burst_1x_r[1] .power_up = "low";

dffeas \dqs_burst_2x_r1[1] (
	.clk(mem_clk_2x),
	.d(\dqs_burst_1x_r[1]~q ),
	.asdata(vcc),
	.clrn(reset_mem_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst_2x_r1[1]~q ),
	.prn(vcc));
defparam \dqs_burst_2x_r1[1] .is_wysiwyg = "true";
defparam \dqs_burst_2x_r1[1] .power_up = "low";

arriaii_lcell_comb \dqs_burst_2x_r2~1 (
	.dataa(!\dqs_burst_sel[1]~q ),
	.datab(!\dqs_burst_2x_r1[5]~q ),
	.datac(!\dqs_burst_2x_r1[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dqs_burst_2x_r2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dqs_burst_2x_r2~1 .extended_lut = "off";
defparam \dqs_burst_2x_r2~1 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \dqs_burst_2x_r2~1 .shared_arith = "off";

dffeas \dqs_burst_2x_r2[1] (
	.clk(mem_clk_2x),
	.d(\dqs_burst_2x_r2~1_combout ),
	.asdata(vcc),
	.clrn(reset_mem_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst_2x_r2[1]~q ),
	.prn(vcc));
defparam \dqs_burst_2x_r2[1] .is_wysiwyg = "true";
defparam \dqs_burst_2x_r2[1] .power_up = "low";

dffeas \dqs_burst_1x_r[6] (
	.clk(phy_clk_1x),
	.d(\mem_dqs_burst[4]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst_1x_r[6]~q ),
	.prn(vcc));
defparam \dqs_burst_1x_r[6] .is_wysiwyg = "true";
defparam \dqs_burst_1x_r[6] .power_up = "low";

dffeas \dqs_burst_2x_r1[6] (
	.clk(mem_clk_2x),
	.d(\dqs_burst_1x_r[6]~q ),
	.asdata(vcc),
	.clrn(reset_mem_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst_2x_r1[6]~q ),
	.prn(vcc));
defparam \dqs_burst_2x_r1[6] .is_wysiwyg = "true";
defparam \dqs_burst_2x_r1[6] .power_up = "low";

dffeas \dqs_burst_1x_r[2] (
	.clk(phy_clk_1x),
	.d(\mem_dqs_burst[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst_1x_r[2]~q ),
	.prn(vcc));
defparam \dqs_burst_1x_r[2] .is_wysiwyg = "true";
defparam \dqs_burst_1x_r[2] .power_up = "low";

dffeas \dqs_burst_2x_r1[2] (
	.clk(mem_clk_2x),
	.d(\dqs_burst_1x_r[2]~q ),
	.asdata(vcc),
	.clrn(reset_mem_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst_2x_r1[2]~q ),
	.prn(vcc));
defparam \dqs_burst_2x_r1[2] .is_wysiwyg = "true";
defparam \dqs_burst_2x_r1[2] .power_up = "low";

arriaii_lcell_comb \dqs_burst_2x_r2~2 (
	.dataa(!\dqs_burst_sel[2]~q ),
	.datab(!\dqs_burst_2x_r1[6]~q ),
	.datac(!\dqs_burst_2x_r1[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dqs_burst_2x_r2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dqs_burst_2x_r2~2 .extended_lut = "off";
defparam \dqs_burst_2x_r2~2 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \dqs_burst_2x_r2~2 .shared_arith = "off";

dffeas \dqs_burst_2x_r2[2] (
	.clk(mem_clk_2x),
	.d(\dqs_burst_2x_r2~2_combout ),
	.asdata(vcc),
	.clrn(reset_mem_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst_2x_r2[2]~q ),
	.prn(vcc));
defparam \dqs_burst_2x_r2[2] .is_wysiwyg = "true";
defparam \dqs_burst_2x_r2[2] .power_up = "low";

dffeas \dqs_burst_1x_r[7] (
	.clk(phy_clk_1x),
	.d(\mem_dqs_burst[4]~0_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst_1x_r[7]~q ),
	.prn(vcc));
defparam \dqs_burst_1x_r[7] .is_wysiwyg = "true";
defparam \dqs_burst_1x_r[7] .power_up = "low";

dffeas \dqs_burst_2x_r1[7] (
	.clk(mem_clk_2x),
	.d(\dqs_burst_1x_r[7]~q ),
	.asdata(vcc),
	.clrn(reset_mem_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst_2x_r1[7]~q ),
	.prn(vcc));
defparam \dqs_burst_2x_r1[7] .is_wysiwyg = "true";
defparam \dqs_burst_2x_r1[7] .power_up = "low";

dffeas \dqs_burst_1x_r[3] (
	.clk(phy_clk_1x),
	.d(\mem_dqs_burst[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset_phy_clk_1x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst_1x_r[3]~q ),
	.prn(vcc));
defparam \dqs_burst_1x_r[3] .is_wysiwyg = "true";
defparam \dqs_burst_1x_r[3] .power_up = "low";

dffeas \dqs_burst_2x_r1[3] (
	.clk(mem_clk_2x),
	.d(\dqs_burst_1x_r[3]~q ),
	.asdata(vcc),
	.clrn(reset_mem_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst_2x_r1[3]~q ),
	.prn(vcc));
defparam \dqs_burst_2x_r1[3] .is_wysiwyg = "true";
defparam \dqs_burst_2x_r1[3] .power_up = "low";

arriaii_lcell_comb \dqs_burst_2x_r2~3 (
	.dataa(!\dqs_burst_sel[3]~q ),
	.datab(!\dqs_burst_2x_r1[7]~q ),
	.datac(!\dqs_burst_2x_r1[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dqs_burst_2x_r2~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dqs_burst_2x_r2~3 .extended_lut = "off";
defparam \dqs_burst_2x_r2~3 .lut_mask = 64'h1B1B1B1B1B1B1B1B;
defparam \dqs_burst_2x_r2~3 .shared_arith = "off";

dffeas \dqs_burst_2x_r2[3] (
	.clk(mem_clk_2x),
	.d(\dqs_burst_2x_r2~3_combout ),
	.asdata(vcc),
	.clrn(reset_mem_clk_2x_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dqs_burst_2x_r2[3]~q ),
	.prn(vcc));
defparam \dqs_burst_2x_r2[3] .is_wysiwyg = "true";
defparam \dqs_burst_2x_r2[3] .power_up = "low";

endmodule
