-- Copyright (C) 1991-2011 Altera Corporation
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs for
-- use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- Quartus II 11.0 Build 157 04/27/2011
LIBRARY IEEE;
use IEEE.STD_LOGIC_1164.all;

package STRATIXV_HSSI_COMPONENTS is

component stratixv_channel_pll
	generic
	(
		avmm_group_channel_index			:	integer	:= 0;
		output_clock_frequency				:	string	:= "0 ps";
		reference_clock_frequency			:	string	:= "0 ps";
		sim_use_fast_model					:	string	:= "true";
		use_default_base_address			:	string	:= "true";
		user_base_address					:	integer	:= 0;
		bbpd_salatch_offset_ctrl_clk0		:	string	:= "clk0_offset_0mv";
		bbpd_salatch_offset_ctrl_clk180		:	string	:= "clk180_offset_0mv";
		bbpd_salatch_offset_ctrl_clk270		:	string	:= "clk270_offset_0mv";
		bbpd_salatch_offset_ctrl_clk90		:	string	:= "clk90_offset_0mv";
		bbpd_salatch_sel					:	string	:= "normal";
		bypass_cp_rgla						:	string	:= "false";
		cdr_atb_select						:	string	:= "atb_disable";
		cgb_clk_enable						:	string	:= "false";
		charge_pump_current_test			:	string	:= "enable_ch_pump_normal";
		clklow_fref_to_ppm_div_sel			:	integer	:= 1;
		clock_monitor						:	string	:= "lpbk_data";
		diag_rev_lpbk						:	string	:= "false";
		eye_monitor_bbpd_data_ctrl			:	string	:= "cdr_data";
		fast_lock_mode						:	string	:= "false";
		fb_sel								:	string	:= "vcoclk";
		gpon_lock2ref_ctrl					:	string	:= "lck2ref";
		hs_levshift_power_supply_setting	:	integer	:= 1;
		ignore_phslock						:	string	:= "false";
		l_counter_pd_clock_disable			:	string	:= "false";
		m_counter							:	integer	:= 25;
		pcie_freq_control					:	string	:= "pcie_100mhz";
		pd_charge_pump_current_ctrl			:	integer	:= 5;
		pd_l_counter						:	integer	:= 1;
		pfd_charge_pump_current_ctrl		:	integer	:= 20;
		pfd_l_counter						:	integer	:= 1;
		powerdown							:	string	:= "false";
		ref_clk_div							:	integer	:= 1;
		regulator_volt_inc					:	string	:= "volt_inc_0pct";
		replica_bias_ctrl					:	string	:= "true";
		reverse_serial_lpbk					:	string	:= "false";
		ripple_cap_ctrl						:	string	:= "none";
		rxpll_pd_bw_ctrl					:	integer	:= 300;
		rxpll_pfd_bw_ctrl					:	integer	:= 3200;
		txpll_hclk_driver_enable			:	string	:= "false";
		vco_overange_ref					:	string	:= "off";
		vco_range_ctrl_en					:	string	:= "false"
	);
	port
	(
		avmmaddress							:	in		std_logic_vector(10 downto 0);
		avmmbyteen							:	in		std_logic;
		avmmclk								:	in		std_logic;
		avmmread							:	in		std_logic;
		avmmrstn							:	in		std_logic;
		avmmwrite							:	in		std_logic;
		avmmwritedata						:	in		std_logic_vector(15 downto 0);
		clk270eye							:   in		std_logic;
		clk270beyerm						:	in		std_logic;
		clk90eye							:   in		std_logic;
		clk90beyerm							:	in		std_logic;
		clkindeser							:	in		std_logic;
		crurstb								:   in		std_logic;
		deeye								:   in		std_logic;
		deeyerm								:   in		std_logic;
		doeye								:   in		std_logic;
		doeyerm								:   in		std_logic;
		earlyeios							:   in		std_logic;
		extclk								:	in		std_logic;
		extfbctrla							:	in		std_logic;
		extfbctrlb							:	in		std_logic;
		gpblck2refb							:	in		std_logic;
		lpbkpreen							:	in		std_logic;
		ltd									:	in		std_logic;
		ltr									:	in		std_logic;
		occalen								:	in		std_logic;
		pciel								:	in		std_logic;
		pciem								:	in		std_logic;
		pciesw								:	in		std_logic_vector(1 downto 0);
		ppmlock								:	in		std_logic;
		refclk								:	in		std_logic;
		rstn								:	in		std_logic;
		rxp									:	in		std_logic;
		sd									:	in		std_logic;
		avmmreaddata						:	out		std_logic_vector(15 downto 0);
		blockselect							:	out		std_logic;
		ck0pd								:	out		std_logic;
		ck180pd								:	out		std_logic;
		ck270pd								:	out		std_logic;
		ck90pd								:	out		std_logic;
		clk270bcdr							:	out		std_logic;
		clk270bdes							:	out		std_logic;
		clk90bcdr							:	out		std_logic;
		clk90bdes							:	out		std_logic;
		clkcdr								:	out		std_logic;
		clklow								:	out		std_logic;
		decdr								:	out		std_logic;
		deven								:	out		std_logic;
		docdr								:	out		std_logic;
		dodd								:	out		std_logic;
		fref								:	out		std_logic;
		pdof								:	out		std_logic_vector(3 downto 0);
		pfdmodelock							:	out		std_logic;
		rxlpbdp								:	out		std_logic;
		rxlpbp								:	out		std_logic;
		rxplllock							:	out		std_logic;
		txpllhclk							:	out		std_logic;
		txrlpbk								:	out		std_logic;
		vctrloverrange						:	out		std_logic
	);
end component;

component stratixv_atx_pll
	generic
	(
         avmm_group_channel_index                :  integer  := 0 ;
         output_clock_frequency                  :  string   := "" ;
         reference_clock_frequency               :  string   := "" ;
         use_default_base_address                :  string   := "true" ;
         user_base_address0                      :  integer  := 0 ;
         user_base_address1                      :  integer  := 0 ;
         user_base_address2                      :  integer  := 0 ;
         cp_current_ctrl                         :  integer  := 300 ;
         cp_current_test                         :  string   := "enable_ch_pump_normal" ;
         cp_hs_levshift_power_supply_setting     :  integer  := 1 ;
         cp_replica_bias_ctrl                    :  string   := "disable_replica_bias_ctrl" ;
         cp_rgla_bypass                          :  string   := "false" ;
         cp_rgla_volt_inc                        :  string   := "boost_30pct" ;
         l_counter                               :  integer  := 1 ;
         lcpll_atb_select                        :  string   := "atb_disable" ;
         lcpll_d2a_sel                           :  string   := "volt_1p02v" ;
         lcpll_hclk_driver_enable                :  string   := "driver_off" ;
         lcvco_gear_sel                          :  string   := "high_gear" ;
         lcvco_sel                               :  string   := "high_freq_14g" ;
         lpf_ripple_cap_ctrl                     :  string   := "none" ;
         lpf_rxpll_pfd_bw_ctrl                   :  integer  := 2400 ;
         m_counter                               :  integer  := 4 ;
         ref_clk_div                             :  integer  := 1 ;
         refclk_sel                              :  string   := "refclk" ;
         vreg1_lcvco_volt_inc                    :  string   := "volt_1p1v" ;
         vreg1_vccehlow                          :  string   := "normal_operation" ;
         vreg2_lcpll_volt_sel                    :  string   := "vreg2_volt_1p0v" ;
         vreg3_lcpll_volt_sel                    :  string   := "vreg3_volt_1p0v"
	);
	port
	(
           avmmaddress        :     in   std_logic_vector( 10 downto 0 );
           avmmbyteen         :     in   std_logic_vector( 1 downto 0 );
           avmmclk            :     in   std_logic;
           avmmread           :     in   std_logic;
           avmmrstn           :     in   std_logic;
           avmmwrite          :     in   std_logic;
           avmmwritedata      :     in   std_logic_vector( 15 downto 0 );
           avmmreaddata       :     out  std_logic_vector( 15 downto 0 );
           blockselect        :     out  std_logic;
           ch0rcsrlc          :     in   std_logic_vector( 31 downto 0 );
           ch1rcsrlc          :     in   std_logic_vector( 31 downto 0 );
           ch2rcsrlc          :     in   std_logic_vector( 31 downto 0 );
           cmurstn            :     in   std_logic;
           cmurstnlpf         :     in   std_logic;
           extfbclk           :     in   std_logic;
           iqclklc            :     in   std_logic;
           pldclklc           :     in   std_logic;
           pllfbswblc         :     in   std_logic;
           pllfbswtlc         :     in   std_logic;
           refclklc           :     in   std_logic;
           clk010g            :     out  std_logic;
           clk025g            :     out  std_logic;
           clk18010g          :     out  std_logic;
           clk18025g          :     out  std_logic;
           clk33cmu           :     out  std_logic;
           clklowcmu          :     out  std_logic;
           frefcmu            :     out  std_logic;
           iqclkatt           :     out  std_logic;
           pfdmodelockcmu     :     out  std_logic;
           pldclkatt          :     out  std_logic;
           refclkatt          :     out  std_logic;
           txpllhclk          :     out  std_logic
	);
end component;


component    stratixv_hssi_10g_rx_pcs
    generic    (
        prot_mode    :    string    :=    "disable_mode";
        sup_mode    :    string    :=    "full_mode";
        dis_signal_ok    :    string    :=    "dis_signal_ok_dis";
        gb_rx_idwidth    :    string    :=    "idwidth_32";
        gb_rx_odwidth    :    string    :=    "odwidth_66";
        bit_reverse    :    string    :=    "bit_reverse_dis";
        gb_sel_mode    :    string    :=    "internal";
        lpbk_mode    :    string    :=    "lpbk_dis";
        test_mode    :    string    :=    "test_off";
        blksync_bypass    :    string    :=    "blksync_bypass_dis";
        blksync_pipeln    :    string    :=    "blksync_pipeln_dis";
        blksync_knum_sh_cnt_prelock    :    string    :=    "int";
        blksync_knum_sh_cnt_postlock    :    string    :=    "int";
        blksync_enum_invalid_sh_cnt    :    string    :=    "int";
        blksync_bitslip_wait_cnt    :    string    :=    "int";
        bitslip_wait_cnt_user    :    string    :=    "int";
        blksync_bitslip_type    :    string    :=    "bitslip_comb";
        blksync_bitslip_wait_type    :    string    :=    "bitslip_match";
        dispchk_bypass    :    string    :=    "dispchk_bypass_dis";
        dispchk_rd_level    :    string    :=    "dispchk_rd_level_min";
        dispchk_rd_level_user    :    string    :=    "int";
        dispchk_pipeln    :    string    :=    "dispchk_pipeln_dis";
        descrm_bypass    :    string    :=    "descrm_bypass_en";
        descrm_mode    :    string    :=    "async";
        frmsync_bypass    :    string    :=    "frmsync_bypass_dis";
        frmsync_pipeln    :    string    :=    "frmsync_pipeln_dis";
        frmsync_mfrm_length    :    string    :=    "int";
        frmsync_mfrm_length_user    :    string    :=    "int";
        frmsync_knum_sync    :    string    :=    "int";
        frmsync_enum_sync    :    string    :=    "int";
        frmsync_enum_scrm    :    string    :=    "int";
        frmsync_flag_type    :    string    :=    "all_framing_words";
        dec_64b66b_10g_mode    :    string    :=    "dec_64b66b_10g_mode_en";
        dec_64b66b_rxsm_bypass    :    string    :=    "dec_64b66b_rxsm_bypass_dis";
        rx_sm_bypass    :    string    :=    "rx_sm_bypass_dis";
        rx_sm_pipeln    :    string    :=    "rx_sm_pipeln_dis";
        rx_sm_hiber    :    string    :=    "rx_sm_hiber_en";
        ber_xus_timer_window    :    string    :=    "int";
        ber_bit_err_total_cnt    :    string    :=    "int";
        crcchk_bypass    :    string    :=    "crcchk_bypass_dis";
        crcchk_pipeln    :    string    :=    "crcchk_pipeln_dis";
        crcflag_pipeln    :    string    :=    "crcflag_pipeln_dis";
        crcchk_init    :    string    :=    "crcchk_init_user_setting";
        crcchk_init_user    :    bit_vector    :=    B"11111111111111111111111111111111";
        crcchk_inv    :    string    :=    "crcchk_inv_dis";
        force_align    :    string    :=    "force_align_dis";
        align_del    :    string    :=    "align_del_en";
        control_del    :    bit_vector    :=    B"11110000";
        rxfifo_mode    :    string    :=    "phase_comp";
        master_clk_sel    :    string    :=    "master_rx_pma_clk";
        rd_clk_sel    :    string    :=    "rd_rx_pma_clk";
        gbexp_clken    :    string    :=    "gbexp_clk_dis";
        prbs_clken    :    string    :=    "prbs_clk_dis";
        blksync_clken    :    string    :=    "blksync_clk_dis";
        dispchk_clken    :    string    :=    "dispchk_clk_dis";
        descrm_clken    :    string    :=    "descrm_clk_dis";
        frmsync_clken    :    string    :=    "frmsync_clk_dis";
        dec64b66b_clken    :    string    :=    "dec64b66b_clk_dis";
        ber_clken    :    string    :=    "ber_clk_dis";
        rand_clken    :    string    :=    "rand_clk_dis";
        crcchk_clken    :    string    :=    "crcchk_clk_dis";
        wrfifo_clken    :    string    :=    "wrfifo_clk_dis";
        rdfifo_clken    :    string    :=    "rdfifo_clk_dis";
        rxfifo_pempty    :    string    :=    "pempty_default";
        rxfifo_pfull    :    string    :=    "pfull_default";
        rxfifo_full    :    string    :=    "full_default";
        rxfifo_empty    :    string    :=    "pempty_default";
        bitslip_mode    :    string    :=    "bitslip_dis";
        fast_path    :    string    :=    "fast_path_dis";
        stretch_num_stages    :    string    :=    "zero_stage";
        stretch_en    :    string    :=    "stretch_en";
        iqtxrx_clkout_sel    :    string    :=    "iq_rx_clk_out";
        channel_number    :    integer    :=    0;
        frmgen_diag_word    :    bit_vector    :=    B"0000000000000000011001000000000000000000000000000000000000000000";
        frmgen_scrm_word    :    bit_vector    :=    B"0000000000000000001010000000000000000000000000000000000000000000";
        frmgen_skip_word    :    bit_vector    :=    B"0000000000000000000111100001111000011110000111100001111000011110";
        frmgen_sync_word    :    bit_vector    :=    B"0000000000000000011110001111011001111000111101100111100011110110";
        test_bus_mode    :    string    :=    "tx"
    );
    port    (
        bercount    :    out    std_logic_vector(5 downto 0);
        errorblockcount    :    out    std_logic_vector(7 downto 0);
        pcsstatus    :    out    std_logic_vector(0 downto 0);
        randomerrorcount    :    out    std_logic_vector(15 downto 0);
        prbserrorlatch    :    out    std_logic_vector(0 downto 0);
        txpmaclk    :    in    std_logic_vector(0 downto 0);
        rxpmaclk    :    in    std_logic_vector(0 downto 0);
        pmaclkdiv33txorrx    :    in    std_logic_vector(0 downto 0);
        rxpmadatavalid    :    in    std_logic_vector(0 downto 0);
        hardresetn    :    in    std_logic_vector(0 downto 0);
        rxpldclk    :    in    std_logic_vector(0 downto 0);
        rxpldrstn    :    in    std_logic_vector(0 downto 0);
        refclkdig    :    in    std_logic_vector(0 downto 0);
        rxalignen    :    in    std_logic_vector(0 downto 0);
        rxalignclr    :    in    std_logic_vector(0 downto 0);
        rxrden    :    in    std_logic_vector(0 downto 0);
        rxdisparityclr    :    in    std_logic_vector(0 downto 0);
        rxclrerrorblockcount    :    in    std_logic_vector(0 downto 0);
        rxclrbercount    :    in    std_logic_vector(0 downto 0);
        rxbitslip    :    in    std_logic_vector(0 downto 0);
        rxprbserrorclr    :    in    std_logic_vector(0 downto 0);
        rxclkout    :    out    std_logic_vector(0 downto 0);
        rxclkiqout    :    out    std_logic_vector(0 downto 0);
        rxdatavalid    :    out    std_logic_vector(0 downto 0);
        rxfifoempty    :    out    std_logic_vector(0 downto 0);
        rxfifopartialempty    :    out    std_logic_vector(0 downto 0);
        rxfifopartialfull    :    out    std_logic_vector(0 downto 0);
        rxfifofull    :    out    std_logic_vector(0 downto 0);
        rxalignval    :    out    std_logic_vector(0 downto 0);
        rxblocklock    :    out    std_logic_vector(0 downto 0);
        rxsyncheadererror    :    out    std_logic_vector(0 downto 0);
        rxhighber    :    out    std_logic_vector(0 downto 0);
        rxframelock    :    out    std_logic_vector(0 downto 0);
        rxrdpossts    :    out    std_logic_vector(0 downto 0);
        rxrdnegsts    :    out    std_logic_vector(0 downto 0);
        rxskipinserted    :    out    std_logic_vector(0 downto 0);
        rxrxframe    :    out    std_logic_vector(0 downto 0);
        rxpayloadinserted    :    out    std_logic_vector(0 downto 0);
        rxsyncworderror    :    out    std_logic_vector(0 downto 0);
        rxscramblererror    :    out    std_logic_vector(0 downto 0);
        rxskipworderror    :    out    std_logic_vector(0 downto 0);
        rxdiagnosticerror    :    out    std_logic_vector(0 downto 0);
        rxmetaframeerror    :    out    std_logic_vector(0 downto 0);
        rxcrc32error    :    out    std_logic_vector(0 downto 0);
        rxdiagnosticstatus    :    out    std_logic_vector(1 downto 0);
        rxdata    :    out    std_logic_vector(63 downto 0);
        rxcontrol    :    out    std_logic_vector(9 downto 0);
        accumdisparity    :    out    std_logic_vector(8 downto 0);
        loopbackdatain    :    in    std_logic_vector(39 downto 0);
        rxpmadata    :    in    std_logic_vector(39 downto 0);
        rxtestdata    :    out    std_logic_vector(19 downto 0);
        syncdatain    :    out    std_logic_vector(0 downto 0)
    );
end component; --stratixv_hssi_10g_rx_pcs


component    stratixv_hssi_10g_tx_pcs
    generic    (
        prot_mode    :    string    :=    "disable_mode";
        sup_mode    :    string    :=    "full_mode";
        ctrl_plane_bonding    :    string    :=    "individual";
        master_clk_sel    :    string    :=    "master_tx_pma_clk";
        wr_clk_sel    :    string    :=    "wr_tx_pma_clk";
        wrfifo_clken    :    string    :=    "wrfifo_clk_dis";
        rdfifo_clken    :    string    :=    "rdfifo_clk_dis";
        frmgen_clken    :    string    :=    "frmgen_clk_dis";
        crcgen_clken    :    string    :=    "crcgen_clk_dis";
        enc64b66b_txsm_clken    :    string    :=    "enc64b66b_txsm_clk_dis";
        scrm_clken    :    string    :=    "scrm_clk_dis";
        dispgen_clken    :    string    :=    "dispgen_clk_dis";
        prbs_clken    :    string    :=    "prbs_clk_dis";
        sqwgen_clken    :    string    :=    "sqwgen_clk_dis";
        gbred_clken    :    string    :=    "gbred_clk_dis";
        gb_tx_idwidth    :    string    :=    "idwidth_50";
        gb_tx_odwidth    :    string    :=    "odwidth_32";
        txfifo_mode    :    string    :=    "phase_comp";
        txfifo_pempty    :    string    :=    "pempty_default";
        txfifo_pfull    :    string    :=    "pfull_default";
        txfifo_empty    :    string    :=    "empty_default";
        txfifo_full    :    string    :=    "full_default";
        frmgen_bypass    :    string    :=    "frmgen_bypass_dis";
        frmgen_pipeln    :    string    :=    "frmgen_pipeln_dis";
        frmgen_mfrm_length    :    string    :=    "frmgen_mfrm_length_min";
        frmgen_mfrm_length_user    :    string    :=    "int";
        frmgen_pyld_ins    :    string    :=    "frmgen_pyld_ins_dis";
        sh_err    :    string    :=    "sh_err_dis";
        frmgen_burst    :    string    :=    "frmgen_burst_dis";
        frmgen_wordslip    :    string    :=    "frmgen_wordslip_dis";
        crcgen_bypass    :    string    :=    "crcgen_bypass_dis";
        crcgen_init    :    string    :=    "crcgen_init_user_setting";
        crcgen_init_user    :    bit_vector    :=    B"11111111111111111111111111111111";
        crcgen_inv    :    string    :=    "crcgen_inv_dis";
        crcgen_err    :    string    :=    "crcgen_err_dis";
        enc_64b66b_10g_mode    :    string    :=    "enc_64b66b_10g_mode_en";
        enc_64b66b_txsm_bypass    :    string    :=    "enc_64b66b_txsm_bypass_dis";
        tx_sm_bypass    :    string    :=    "tx_sm_bypass_dis";
        tx_sm_pipeln    :    string    :=    "tx_sm_pipeln_dis";
        scrm_bypass    :    string    :=    "scrm_bypass_dis";
        test_mode    :    string    :=    "test_off";
        pseudo_random    :    string    :=    "all_0";
        pseudo_seed_a    :    string    :=    "pseudo_seed_a_user_setting";
        pseudo_seed_a_user    :    bit_vector    :=    B"1111111111111111111111111111111111111111111111111111111111";
        pseudo_seed_b    :    string    :=    "pseudo_seed_b_user_setting";
        pseudo_seed_b_user    :    bit_vector    :=    B"1111111111111111111111111111111111111111111111111111111111";
        bit_reverse    :    string    :=    "bit_reverse_dis";
        scrm_seed    :    string    :=    "scram_seed_user_setting";
        scrm_seed_user    :    bit_vector    :=    B"1111111111111111111111111111111111111111111111111111111111";
        scrm_mode    :    string    :=    "async";
        dispgen_bypass    :    string    :=    "dispgen_bypass_dis";
        dispgen_err    :    string    :=    "dispgen_err_dis";
        dispgen_pipeln    :    string    :=    "dispgen_pipeln_dis";
        gb_sel_mode    :    string    :=    "internal";
        sq_wave    :    string    :=    "sq_wave_4";
        bitslip_en    :    string    :=    "bitslip_dis";
        fastpath    :    string    :=    "fastpath_dis";
        distup_bypass_pipeln    :    string    :=    "distup_bypass_pipeln_dis";
        distup_master    :    string    :=    "distup_master_en";
        distdwn_bypass_pipeln    :    string    :=    "distdwn_bypass_pipeln_dis";
        distdwn_master    :    string    :=    "distdwn_master_en";
        compin_sel    :    string    :=    "compin_master";
        comp_cnt    :    string    :=    "comp_cnt_00";
        indv    :    string    :=    "indv_en";
        stretch_num_stages    :    string    :=    "zero_stage";
        stretch_en    :    string    :=    "stretch_en";
        iqtxrx_clkout_sel    :    string    :=    "iq_tx_pma_clk";
        channel_number    :    integer    :=    0;
        frmgen_sync_word    :    bit_vector    :=    B"0000000000000000011110001111011001111000111101100111100011110110";
        frmgen_scrm_word    :    bit_vector    :=    B"0000000000000000001010000000000000000000000000000000000000000000";
        frmgen_skip_word    :    bit_vector    :=    B"0000000000000000000111100001111000011110000111100001111000011110";
        frmgen_diag_word    :    bit_vector    :=    B"0000000000000000011001000000000000000000000000000000000000000000";
        test_bus_mode    :    string    :=    "tx";
        lpm_type    :    string    :=    "stratixv_hssi_10g_tx_pcs"
    );
    port    (
        txpmaclk    :    in    std_logic_vector(0 downto 0);
        pmaclkdiv33lc    :    in    std_logic_vector(0 downto 0);
        hardresetn    :    in    std_logic_vector(0 downto 0);
        txpldclk    :    in    std_logic_vector(0 downto 0);
        txpldrstn    :    in    std_logic_vector(0 downto 0);
        refclkdig    :    in    std_logic_vector(0 downto 0);
        txdatavalid    :    in    std_logic_vector(0 downto 0);
        txbitslip    :    in    std_logic_vector(6 downto 0);
        txdiagnosticstatus    :    in    std_logic_vector(1 downto 0);
        txwordslip    :    in    std_logic_vector(0 downto 0);
        txbursten    :    in    std_logic_vector(0 downto 0);
        txdisparityclr    :    in    std_logic_vector(0 downto 0);
        txclkout    :    out    std_logic_vector(0 downto 0);
        txclkiqout    :    out    std_logic_vector(0 downto 0);
        txfifoempty    :    out    std_logic_vector(0 downto 0);
        txfifopartialempty    :    out    std_logic_vector(0 downto 0);
        txfifopartialfull    :    out    std_logic_vector(0 downto 0);
        txfifofull    :    out    std_logic_vector(0 downto 0);
        txframe    :    out    std_logic_vector(0 downto 0);
        txburstenexe    :    out    std_logic_vector(0 downto 0);
        txwordslipexe    :    out    std_logic_vector(0 downto 0);
        distupindv    :    in    std_logic_vector(0 downto 0);
        distdwnindv    :    in    std_logic_vector(0 downto 0);
        distupinwren    :    in    std_logic_vector(0 downto 0);
        distdwninwren    :    in    std_logic_vector(0 downto 0);
        distupinrden    :    in    std_logic_vector(0 downto 0);
        distdwninrden    :    in    std_logic_vector(0 downto 0);
        distupoutdv    :    out    std_logic_vector(0 downto 0);
        distdwnoutdv    :    out    std_logic_vector(0 downto 0);
        distupoutwren    :    out    std_logic_vector(0 downto 0);
        distdwnoutwren    :    out    std_logic_vector(0 downto 0);
        distupoutrden    :    out    std_logic_vector(0 downto 0);
        distdwnoutrden    :    out    std_logic_vector(0 downto 0);
        txtestdata    :    out    std_logic_vector(19 downto 0);
        txdata    :    in    std_logic_vector(63 downto 0);
        txcontrol    :    in    std_logic_vector(8 downto 0);
        loopbackdataout    :    out    std_logic_vector(39 downto 0);
        txpmadata    :    out    std_logic_vector(39 downto 0);
        syncdatain    :    out    std_logic_vector(0 downto 0)
    );
end component; --stratixv_hssi_10g_tx_pcs


component    stratixv_hssi_8g_pcs_aggregate
    generic    (
        xaui_sm_operation    :    string    :=    "en_xaui_sm";
        dskw_sm_operation    :    string    :=    "dskw_xaui_sm";
        data_agg_bonding    :    string    :=    "agg_disable";
        prot_mode_tx    :    string    :=    "pipe_g1_tx";
        pcs_dw_datapath    :    string    :=    "sw_data_path";
        dskw_control    :    string    :=    "dskw_write_control";
        refclkdig_sel    :    string    :=    "dis_refclk_dig_sel"
    );
    port    (
        refclkdig    :    in    std_logic_vector(0 downto 0);
        scanmoden    :    in    std_logic_vector(0 downto 0);
        scanshiftn    :    in    std_logic_vector(0 downto 0);
        txpmaclk    :    in    std_logic_vector(0 downto 0);
        rcvdclkch0    :    in    std_logic_vector(0 downto 0);
        rcvdclkch1    :    in    std_logic_vector(0 downto 0);
        hardrst    :    in    std_logic_vector(0 downto 0);
        txpcsrst    :    in    std_logic_vector(0 downto 0);
        rxpcsrst    :    in    std_logic_vector(0 downto 0);
        dprioagg    :    in    std_logic_vector(63 downto 0);
        rcvdclkout    :    out    std_logic_vector(0 downto 0);
        rcvdclkouttop    :    out    std_logic_vector(0 downto 0);
        rcvdclkoutbot    :    out    std_logic_vector(0 downto 0);
        rdenablesynctopch1    :    in    std_logic_vector(0 downto 0);
        txdatatctopch1    :    in    std_logic_vector(7 downto 0);
        txctltctopch1    :    in    std_logic_vector(0 downto 0);
        syncstatustopch1    :    in    std_logic_vector(0 downto 0);
        rdaligntopch1    :    in    std_logic_vector(1 downto 0);
        aligndetsynctopch1    :    in    std_logic_vector(1 downto 0);
        fifordintopch1    :    in    std_logic_vector(0 downto 0);
        alignstatussynctopch1    :    in    std_logic_vector(0 downto 0);
        cgcomprddintopch1    :    in    std_logic_vector(1 downto 0);
        cgcompwrintopch1    :    in    std_logic_vector(1 downto 0);
        delcondmetintopch1    :    in    std_logic_vector(0 downto 0);
        fifoovrintopch1    :    in    std_logic_vector(0 downto 0);
        latencycompintopch1    :    in    std_logic_vector(0 downto 0);
        insertincompleteintopch1    :    in    std_logic_vector(0 downto 0);
        decdatatopch1    :    in    std_logic_vector(7 downto 0);
        decctltopch1    :    in    std_logic_vector(0 downto 0);
        decdatavalidtopch1    :    in    std_logic_vector(0 downto 0);
        runningdisptopch1    :    in    std_logic_vector(1 downto 0);
        txdatatstopch1    :    out    std_logic_vector(7 downto 0);
        txctltstopch1    :    out    std_logic_vector(0 downto 0);
        fiforstrdqdtopch1    :    out    std_logic_vector(0 downto 0);
        endskwqdtopch1    :    out    std_logic_vector(0 downto 0);
        endskwrdptrstopch1    :    out    std_logic_vector(0 downto 0);
        alignstatustopch1    :    out    std_logic_vector(0 downto 0);
        alignstatussync0topch1    :    out    std_logic_vector(0 downto 0);
        fifordoutcomp0topch1    :    out    std_logic_vector(0 downto 0);
        cgcomprddalltopch1    :    out    std_logic_vector(0 downto 0);
        cgcompwralltopch1    :    out    std_logic_vector(0 downto 0);
        delcondmet0topch1    :    out    std_logic_vector(0 downto 0);
        insertincomplete0topch1    :    out    std_logic_vector(0 downto 0);
        fifoovr0topch1    :    out    std_logic_vector(0 downto 0);
        latencycomp0topch1    :    out    std_logic_vector(0 downto 0);
        rxdatarstopch1    :    out    std_logic_vector(7 downto 0);
        rxctlrstopch1    :    out    std_logic_vector(0 downto 0);
        rdenablesynctopch0    :    in    std_logic_vector(0 downto 0);
        txdatatctopch0    :    in    std_logic_vector(7 downto 0);
        txctltctopch0    :    in    std_logic_vector(0 downto 0);
        syncstatustopch0    :    in    std_logic_vector(0 downto 0);
        rdaligntopch0    :    in    std_logic_vector(1 downto 0);
        aligndetsynctopch0    :    in    std_logic_vector(1 downto 0);
        fifordintopch0    :    in    std_logic_vector(0 downto 0);
        alignstatussynctopch0    :    in    std_logic_vector(0 downto 0);
        cgcomprddintopch0    :    in    std_logic_vector(1 downto 0);
        cgcompwrintopch0    :    in    std_logic_vector(1 downto 0);
        delcondmetintopch0    :    in    std_logic_vector(0 downto 0);
        fifoovrintopch0    :    in    std_logic_vector(0 downto 0);
        latencycompintopch0    :    in    std_logic_vector(0 downto 0);
        insertincompleteintopch0    :    in    std_logic_vector(0 downto 0);
        decdatatopch0    :    in    std_logic_vector(7 downto 0);
        decctltopch0    :    in    std_logic_vector(0 downto 0);
        decdatavalidtopch0    :    in    std_logic_vector(0 downto 0);
        runningdisptopch0    :    in    std_logic_vector(1 downto 0);
        txdatatstopch0    :    out    std_logic_vector(7 downto 0);
        txctltstopch0    :    out    std_logic_vector(0 downto 0);
        fiforstrdqdtopch0    :    out    std_logic_vector(0 downto 0);
        endskwqdtopch0    :    out    std_logic_vector(0 downto 0);
        endskwrdptrstopch0    :    out    std_logic_vector(0 downto 0);
        alignstatustopch0    :    out    std_logic_vector(0 downto 0);
        alignstatussync0topch0    :    out    std_logic_vector(0 downto 0);
        fifordoutcomp0topch0    :    out    std_logic_vector(0 downto 0);
        cgcomprddalltopch0    :    out    std_logic_vector(0 downto 0);
        cgcompwralltopch0    :    out    std_logic_vector(0 downto 0);
        delcondmet0topch0    :    out    std_logic_vector(0 downto 0);
        insertincomplete0topch0    :    out    std_logic_vector(0 downto 0);
        fifoovr0topch0    :    out    std_logic_vector(0 downto 0);
        latencycomp0topch0    :    out    std_logic_vector(0 downto 0);
        rxdatarstopch0    :    out    std_logic_vector(7 downto 0);
        rxctlrstopch0    :    out    std_logic_vector(0 downto 0);
        rdenablesyncch2    :    in    std_logic_vector(0 downto 0);
        txdatatcch2    :    in    std_logic_vector(7 downto 0);
        txctltcch2    :    in    std_logic_vector(0 downto 0);
        syncstatusch2    :    in    std_logic_vector(0 downto 0);
        rdalignch2    :    in    std_logic_vector(1 downto 0);
        aligndetsyncch2    :    in    std_logic_vector(1 downto 0);
        fifordinch2    :    in    std_logic_vector(0 downto 0);
        alignstatussyncch2    :    in    std_logic_vector(0 downto 0);
        cgcomprddinch2    :    in    std_logic_vector(1 downto 0);
        cgcompwrinch2    :    in    std_logic_vector(1 downto 0);
        delcondmetinch2    :    in    std_logic_vector(0 downto 0);
        fifoovrinch2    :    in    std_logic_vector(0 downto 0);
        latencycompinch2    :    in    std_logic_vector(0 downto 0);
        insertincompleteinch2    :    in    std_logic_vector(0 downto 0);
        decdatach2    :    in    std_logic_vector(7 downto 0);
        decctlch2    :    in    std_logic_vector(0 downto 0);
        decdatavalidch2    :    in    std_logic_vector(0 downto 0);
        runningdispch2    :    in    std_logic_vector(1 downto 0);
        txdatatsch2    :    out    std_logic_vector(7 downto 0);
        txctltsch2    :    out    std_logic_vector(0 downto 0);
        fiforstrdqdch2    :    out    std_logic_vector(0 downto 0);
        endskwqdch2    :    out    std_logic_vector(0 downto 0);
        endskwrdptrsch2    :    out    std_logic_vector(0 downto 0);
        alignstatusch2    :    out    std_logic_vector(0 downto 0);
        alignstatussync0ch2    :    out    std_logic_vector(0 downto 0);
        fifordoutcomp0ch2    :    out    std_logic_vector(0 downto 0);
        cgcomprddallch2    :    out    std_logic_vector(0 downto 0);
        cgcompwrallch2    :    out    std_logic_vector(0 downto 0);
        delcondmet0ch2    :    out    std_logic_vector(0 downto 0);
        insertincomplete0ch2    :    out    std_logic_vector(0 downto 0);
        fifoovr0ch2    :    out    std_logic_vector(0 downto 0);
        latencycomp0ch2    :    out    std_logic_vector(0 downto 0);
        rxdatarsch2    :    out    std_logic_vector(7 downto 0);
        rxctlrsch2    :    out    std_logic_vector(0 downto 0);
        rdenablesyncch1    :    in    std_logic_vector(0 downto 0);
        txdatatcch1    :    in    std_logic_vector(7 downto 0);
        txctltcch1    :    in    std_logic_vector(0 downto 0);
        syncstatusch1    :    in    std_logic_vector(0 downto 0);
        rdalignch1    :    in    std_logic_vector(1 downto 0);
        aligndetsyncch1    :    in    std_logic_vector(1 downto 0);
        fifordinch1    :    in    std_logic_vector(0 downto 0);
        alignstatussyncch1    :    in    std_logic_vector(0 downto 0);
        cgcomprddinch1    :    in    std_logic_vector(1 downto 0);
        cgcompwrinch1    :    in    std_logic_vector(1 downto 0);
        delcondmetinch1    :    in    std_logic_vector(0 downto 0);
        fifoovrinch1    :    in    std_logic_vector(0 downto 0);
        latencycompinch1    :    in    std_logic_vector(0 downto 0);
        insertincompleteinch1    :    in    std_logic_vector(0 downto 0);
        decdatach1    :    in    std_logic_vector(7 downto 0);
        decctlch1    :    in    std_logic_vector(0 downto 0);
        decdatavalidch1    :    in    std_logic_vector(0 downto 0);
        runningdispch1    :    in    std_logic_vector(1 downto 0);
        txdatatsch1    :    out    std_logic_vector(7 downto 0);
        txctltsch1    :    out    std_logic_vector(0 downto 0);
        fiforstrdqdch1    :    out    std_logic_vector(0 downto 0);
        endskwqdch1    :    out    std_logic_vector(0 downto 0);
        endskwrdptrsch1    :    out    std_logic_vector(0 downto 0);
        alignstatusch1    :    out    std_logic_vector(0 downto 0);
        alignstatussync0ch1    :    out    std_logic_vector(0 downto 0);
        fifordoutcomp0ch1    :    out    std_logic_vector(0 downto 0);
        cgcomprddallch1    :    out    std_logic_vector(0 downto 0);
        cgcompwrallch1    :    out    std_logic_vector(0 downto 0);
        delcondmet0ch1    :    out    std_logic_vector(0 downto 0);
        insertincomplete0ch1    :    out    std_logic_vector(0 downto 0);
        fifoovr0ch1    :    out    std_logic_vector(0 downto 0);
        latencycomp0ch1    :    out    std_logic_vector(0 downto 0);
        rxdatarsch1    :    out    std_logic_vector(7 downto 0);
        rxctlrsch1    :    out    std_logic_vector(0 downto 0);
        rdenablesyncch0    :    in    std_logic_vector(0 downto 0);
        txdatatcch0    :    in    std_logic_vector(7 downto 0);
        txctltcch0    :    in    std_logic_vector(0 downto 0);
        syncstatusch0    :    in    std_logic_vector(0 downto 0);
        rdalignch0    :    in    std_logic_vector(1 downto 0);
        aligndetsyncch0    :    in    std_logic_vector(1 downto 0);
        fifordinch0    :    in    std_logic_vector(0 downto 0);
        alignstatussyncch0    :    in    std_logic_vector(0 downto 0);
        cgcomprddinch0    :    in    std_logic_vector(1 downto 0);
        cgcompwrinch0    :    in    std_logic_vector(1 downto 0);
        delcondmetinch0    :    in    std_logic_vector(0 downto 0);
        fifoovrinch0    :    in    std_logic_vector(0 downto 0);
        latencycompinch0    :    in    std_logic_vector(0 downto 0);
        insertincompleteinch0    :    in    std_logic_vector(0 downto 0);
        decdatach0    :    in    std_logic_vector(7 downto 0);
        decctlch0    :    in    std_logic_vector(0 downto 0);
        decdatavalidch0    :    in    std_logic_vector(0 downto 0);
        runningdispch0    :    in    std_logic_vector(1 downto 0);
        txdatatsch0    :    out    std_logic_vector(7 downto 0);
        txctltsch0    :    out    std_logic_vector(0 downto 0);
        fiforstrdqdch0    :    out    std_logic_vector(0 downto 0);
        endskwqdch0    :    out    std_logic_vector(0 downto 0);
        endskwrdptrsch0    :    out    std_logic_vector(0 downto 0);
        alignstatusch0    :    out    std_logic_vector(0 downto 0);
        alignstatussync0ch0    :    out    std_logic_vector(0 downto 0);
        fifordoutcomp0ch0    :    out    std_logic_vector(0 downto 0);
        cgcomprddallch0    :    out    std_logic_vector(0 downto 0);
        cgcompwrallch0    :    out    std_logic_vector(0 downto 0);
        delcondmet0ch0    :    out    std_logic_vector(0 downto 0);
        insertincomplete0ch0    :    out    std_logic_vector(0 downto 0);
        fifoovr0ch0    :    out    std_logic_vector(0 downto 0);
        latencycomp0ch0    :    out    std_logic_vector(0 downto 0);
        rxdatarsch0    :    out    std_logic_vector(7 downto 0);
        rxctlrsch0    :    out    std_logic_vector(0 downto 0);
        rdenablesyncbotch2    :    in    std_logic_vector(0 downto 0);
        txdatatcbotch2    :    in    std_logic_vector(7 downto 0);
        txctltcbotch2    :    in    std_logic_vector(0 downto 0);
        syncstatusbotch2    :    in    std_logic_vector(0 downto 0);
        rdalignbotch2    :    in    std_logic_vector(1 downto 0);
        aligndetsyncbotch2    :    in    std_logic_vector(1 downto 0);
        fifordinbotch2    :    in    std_logic_vector(0 downto 0);
        alignstatussyncbotch2    :    in    std_logic_vector(0 downto 0);
        cgcomprddinbotch2    :    in    std_logic_vector(1 downto 0);
        cgcompwrinbotch2    :    in    std_logic_vector(1 downto 0);
        delcondmetinbotch2    :    in    std_logic_vector(0 downto 0);
        fifoovrinbotch2    :    in    std_logic_vector(0 downto 0);
        latencycompinbotch2    :    in    std_logic_vector(0 downto 0);
        insertincompleteinbotch2    :    in    std_logic_vector(0 downto 0);
        decdatabotch2    :    in    std_logic_vector(7 downto 0);
        decctlbotch2    :    in    std_logic_vector(0 downto 0);
        decdatavalidbotch2    :    in    std_logic_vector(0 downto 0);
        runningdispbotch2    :    in    std_logic_vector(1 downto 0);
        txdatatsbotch2    :    out    std_logic_vector(7 downto 0);
        txctltsbotch2    :    out    std_logic_vector(0 downto 0);
        fiforstrdqdbotch2    :    out    std_logic_vector(0 downto 0);
        endskwqdbotch2    :    out    std_logic_vector(0 downto 0);
        endskwrdptrsbotch2    :    out    std_logic_vector(0 downto 0);
        alignstatusbotch2    :    out    std_logic_vector(0 downto 0);
        alignstatussync0botch2    :    out    std_logic_vector(0 downto 0);
        fifordoutcomp0botch2    :    out    std_logic_vector(0 downto 0);
        cgcomprddallbotch2    :    out    std_logic_vector(0 downto 0);
        cgcompwrallbotch2    :    out    std_logic_vector(0 downto 0);
        delcondmet0botch2    :    out    std_logic_vector(0 downto 0);
        insertincomplete0botch2    :    out    std_logic_vector(0 downto 0);
        fifoovr0botch2    :    out    std_logic_vector(0 downto 0);
        latencycomp0botch2    :    out    std_logic_vector(0 downto 0);
        rxdatarsbotch2    :    out    std_logic_vector(7 downto 0);
        rxctlrsbotch2    :    out    std_logic_vector(0 downto 0)
    );
end component; --stratixv_hssi_8g_pcs_aggregate


component    stratixv_hssi_8g_rx_pcs
    generic    (
        prot_mode    :    string    :=    "gige";
        tx_rx_parallel_loopback    :    string    :=    "dis_plpbk";
        pma_dw    :    string    :=    "eight_bit";
        pcs_bypass    :    string    :=    "dis_pcs_bypass";
        polarity_inversion    :    string    :=    "dis_pol_inv";
        wa_pd    :    string    :=    "wa_pd_10";
        wa_pd_data    :    bit_vector    :=    B"0000000000000000000000000000000000000000";
        wa_boundary_lock_ctrl    :    string    :=    "bit_slip";
        wa_pld_controlled    :    string    :=    "dis_pld_ctrl";
        wa_sync_sm_ctrl    :    string    :=    "gige_sync_sm";
        wa_rknumber_data    :    bit_vector    :=    B"00000000";
        wa_renumber_data    :    bit_vector    :=    B"000000";
        wa_rgnumber_data    :    bit_vector    :=    B"00000000";
        wa_rosnumber_data    :    bit_vector    :=    B"00";
        wa_kchar    :    string    :=    "dis_kchar";
        wa_det_latency_sync_status_beh    :    string    :=    "assert_sync_status_non_imm";
        wa_clk_slip_spacing    :    string    :=    "min_clk_slip_spacing";
        wa_clk_slip_spacing_data    :    bit_vector    :=    B"0000010000";
        bit_reversal    :    string    :=    "dis_bit_reversal";
        symbol_swap    :    string    :=    "dis_symbol_swap";
        deskew_pattern    :    bit_vector    :=    B"1101101000";
        deskew_prog_pattern_only    :    string    :=    "en_deskew_prog_pat_only";
        rate_match    :    string    :=    "dis_rm";
        eightb_tenb_decoder    :    string    :=    "dis_8b10b";
        err_flags_sel    :    string    :=    "err_flags_wa";
        polinv_8b10b_dec    :    string    :=    "dis_polinv_8b10b_dec";
        eightbtenb_decoder_output_sel    :    string    :=    "data_8b10b_decoder";
        invalid_code_flag_only    :    string    :=    "dis_invalid_code_only";
        auto_error_replacement    :    string    :=    "dis_err_replace";
        pad_or_edb_error_replace    :    string    :=    "replace_edb";
        byte_deserializer    :    string    :=    "dis_bds";
        byte_order    :    string    :=    "dis_bo";
        re_bo_on_wa    :    string    :=    "dis_re_bo_on_wa";
        bo_pattern    :    bit_vector    :=    B"00000000000000000000";
        bo_pad    :    bit_vector    :=    B"0000000000";
        phase_compensation_fifo    :    string    :=    "low_latency";
        prbs_ver    :    string    :=    "dis_prbs";
        cid_pattern    :    string    :=    "cid_pattern_0";
        cid_pattern_len    :    bit_vector    :=    B"00000000";
        bist_ver    :    string    :=    "dis_bist";
        cdr_ctrl    :    string    :=    "dis_cdr_ctrl";
        cdr_ctrl_rxvalid_mask    :    string    :=    "dis_rxvalid_mask";
        wait_cnt    :    bit_vector    :=    B"00000000";
        mask_cnt    :    bit_vector    :=    B"1111111111";
        auto_deassert_pc_rst_cnt_data    :    bit_vector    :=    B"00000";
        auto_pc_en_cnt_data    :    bit_vector    :=    B"0000000";
        eidle_entry_sd    :    string    :=    "dis_eidle_sd";
        eidle_entry_eios    :    string    :=    "dis_eidle_eios";
        eidle_entry_iei    :    string    :=    "dis_eidle_iei";
        rx_rcvd_clk    :    string    :=    "rcvd_clk_rcvd_clk";
        rx_clk1    :    string    :=    "rcvd_clk_clk1";
        rx_clk2    :    string    :=    "rcvd_clk_clk2";
        rx_rd_clk    :    string    :=    "pld_rx_clk";
        dw_one_or_two_symbol_bo    :    string    :=    "donot_care_one_two_bo";
        comp_fifo_rst_pld_ctrl    :    string    :=    "dis_comp_fifo_rst_pld_ctrl";
        bypass_pipeline_reg    :    string    :=    "dis_bypass_pipeline";
        agg_block_sel    :    string    :=    "same_smrt_pack";
        test_bus_sel    :    string    :=    "test_bus_sel";
        wa_rvnumber_data    :    bit_vector    :=    B"0000000000000";
        ctrl_plane_bonding_compensation    :    string    :=    "dis_compensation";
        clock_gate_rx    :    string    :=    "dis_clk_gating";
        prbs_ver_clr_flag    :    string    :=    "dis_prbs_clr_flag";
        hip_mode    :    string    :=    "dis_hip";
        ctrl_plane_bonding_distribution    :    string    :=    "not_master_chnl_distr";
        ctrl_plane_bonding_consumption    :    string    :=    "individual";
        pma_done_count    :    bit_vector    :=    B"000000000000000000";
        test_mode    :    string    :=    "prbs";
        bist_ver_clr_flag    :    string    :=    "dis_bist_clr_flag";
        wa_disp_err_flag    :    string    :=    "dis_disp_err_flag";
        wait_for_phfifo_cnt_data    :    bit_vector    :=    B"000000";
        runlength_check    :    string    :=    "en_runlength_sw";
        test_bus_sel_val    :    bit_vector    :=    B"0000";
        runlength_val    :    bit_vector    :=    B"000000";
        force_signal_detect    :    string    :=    "en_force_signal_detect";
        deskew    :    string    :=    "dis_deskew";
        rx_wr_clk    :    string    :=    "rx_clk2_div_1_2_4";
        rx_clk_free_running    :    string    :=    "en_rx_clk_free_run";
        rx_pcs_urst    :    string    :=    "en_rx_pcs_urst";
        self_switch_dw_scaling    :    string    :=    "dis_self_switch_dw_scaling";
        pipe_if_enable    :    string    :=    "dis_pipe_rx";
        pc_fifo_rst_pld_ctrl    :    string    :=    "dis_pc_fifo_rst_pld_ctrl";
        auto_speed_nego_gen2    :    string    :=    "dis_auto_speed_nego_g2";
        auto_speed_nego_gen3    :    string    :=    "dis_auto_speed_nego_g3";
        ibm_invalid_code    :    string    :=    "dis_ibm_invalid_code";
        channel_number    :    string    :=    "int";
        rx_refclk    :    string    :=    "dis_refclk_sel"
    );
    port    (
        hrdrst    :    in    std_logic_vector(0 downto 0);
        rxpcsrst    :    in    std_logic_vector(0 downto 0);
        rmfifouserrst    :    in    std_logic_vector(0 downto 0);
        phfifouserrst    :    in    std_logic_vector(0 downto 0);
        scanmode    :    in    std_logic_vector(0 downto 0);
        enablecommadetect    :    in    std_logic_vector(0 downto 0);
        a1a2size    :    in    std_logic_vector(0 downto 0);
        bitslip    :    in    std_logic_vector(0 downto 0);
        rmfiforeadenable    :    in    std_logic_vector(0 downto 0);
        rmfifowriteenable    :    in    std_logic_vector(0 downto 0);
        pldrxclk    :    in    std_logic_vector(0 downto 0);
        softresetrclk1    :    out    std_logic_vector(0 downto 0);
        polinvrx    :    in    std_logic_vector(0 downto 0);
        bitreversalenable    :    in    std_logic_vector(0 downto 0);
        bytereversalenable    :    in    std_logic_vector(0 downto 0);
        rcvdclkpma    :    in    std_logic_vector(0 downto 0);
        datain    :    in    std_logic_vector(19 downto 0);
        sigdetfrompma    :    in    std_logic_vector(0 downto 0);
        fiforstrdqd    :    in    std_logic_vector(0 downto 0);
        endskwqd    :    in    std_logic_vector(0 downto 0);
        endskwrdptrs    :    in    std_logic_vector(0 downto 0);
        alignstatus    :    in    std_logic_vector(0 downto 0);
        fiforstrdqdtoporbot    :    in    std_logic_vector(0 downto 0);
        endskwqdtoporbot    :    in    std_logic_vector(0 downto 0);
        endskwrdptrstoporbot    :    in    std_logic_vector(0 downto 0);
        alignstatustoporbot    :    in    std_logic_vector(0 downto 0);
        datafrinaggblock    :    in    std_logic_vector(7 downto 0);
        ctrlfromaggblock    :    in    std_logic_vector(0 downto 0);
        rxdatarstoporbot    :    in    std_logic_vector(7 downto 0);
        rxcontrolrstoporbot    :    in    std_logic_vector(0 downto 0);
        rcvdclk0pma    :    in    std_logic_vector(0 downto 0);
        parallelloopback    :    in    std_logic_vector(19 downto 0);
        txpmaclk    :    in    std_logic_vector(0 downto 0);
        byteorder    :    in    std_logic_vector(0 downto 0);
        pxfifowrdisable    :    in    std_logic_vector(0 downto 0);
        pcfifordenable    :    in    std_logic_vector(0 downto 0);
        pmatestbus    :    in    std_logic_vector(7 downto 0);
        encodertestbus    :    in    std_logic_vector(9 downto 0);
        txctrltestbus    :    in    std_logic_vector(9 downto 0);
        phystatusinternal    :    in    std_logic_vector(0 downto 0);
        rxvalidinternal    :    in    std_logic_vector(0 downto 0);
        rxstatusinternal    :    in    std_logic_vector(2 downto 0);
        phystatuspcsgen3    :    in    std_logic_vector(0 downto 0);
        rxvalidpcsgen3    :    in    std_logic_vector(0 downto 0);
        rxstatuspcsgen3    :    in    std_logic_vector(2 downto 0);
        rxdatavalidpcsgen3    :    in    std_logic_vector(3 downto 0);
        rxblkstartpcsgen3    :    in    std_logic_vector(3 downto 0);
        rxsynchdrpcsgen3    :    in    std_logic_vector(1 downto 0);
        rxdatapcsgen3    :    in    std_logic_vector(63 downto 0);
        pipepowerdown    :    in    std_logic_vector(1 downto 0);
        rateswitchcontrol    :    in    std_logic_vector(0 downto 0);
        gen2ngen1    :    in    std_logic_vector(0 downto 0);
        gen2ngen1bundle    :    in    std_logic_vector(0 downto 0);
        eidleinfersel    :    in    std_logic_vector(2 downto 0);
        pipeloopbk    :    in    std_logic_vector(0 downto 0);
        pldltr    :    in    std_logic_vector(0 downto 0);
        prbscidenable    :    in    std_logic_vector(0 downto 0);
        txdiv2syncoutpipeup    :    in    std_logic_vector(0 downto 0);
        fifoselectoutpipeup    :    in    std_logic_vector(0 downto 0);
        txwrenableoutpipeup    :    in    std_logic_vector(0 downto 0);
        txrdenableoutpipeup    :    in    std_logic_vector(0 downto 0);
        txdiv2syncoutpipedown    :    in    std_logic_vector(0 downto 0);
        fifoselectoutpipedown    :    in    std_logic_vector(0 downto 0);
        txwrenableoutpipedown    :    in    std_logic_vector(0 downto 0);
        txrdenableoutpipedown    :    in    std_logic_vector(0 downto 0);
        alignstatussync0    :    in    std_logic_vector(0 downto 0);
        rmfifordincomp0    :    in    std_logic_vector(0 downto 0);
        cgcomprddall    :    in    std_logic_vector(0 downto 0);
        cgcompwrall    :    in    std_logic_vector(0 downto 0);
        delcondmet0    :    in    std_logic_vector(0 downto 0);
        fifoovr0    :    in    std_logic_vector(0 downto 0);
        latencycomp0    :    in    std_logic_vector(0 downto 0);
        insertincomplete0    :    in    std_logic_vector(0 downto 0);
        alignstatussync0toporbot    :    in    std_logic_vector(0 downto 0);
        fifordincomp0toporbot    :    in    std_logic_vector(0 downto 0);
        cgcomprddalltoporbot    :    in    std_logic_vector(0 downto 0);
        cgcompwralltoporbot    :    in    std_logic_vector(0 downto 0);
        delcondmet0toporbot    :    in    std_logic_vector(0 downto 0);
        fifoovr0toporbot    :    in    std_logic_vector(0 downto 0);
        latencycomp0toporbot    :    in    std_logic_vector(0 downto 0);
        insertincomplete0toporbot    :    in    std_logic_vector(0 downto 0);
        alignstatussync    :    out    std_logic_vector(0 downto 0);
        fifordoutcomp    :    out    std_logic_vector(0 downto 0);
        cgcomprddout    :    out    std_logic_vector(1 downto 0);
        cgcompwrout    :    out    std_logic_vector(1 downto 0);
        delcondmetout    :    out    std_logic_vector(0 downto 0);
        fifoovrout    :    out    std_logic_vector(0 downto 0);
        latencycompout    :    out    std_logic_vector(0 downto 0);
        insertincompleteout    :    out    std_logic_vector(0 downto 0);
        dataout    :    out    std_logic_vector(63 downto 0);
        parallelrevloopback    :    out    std_logic_vector(19 downto 0);
        clocktopld    :    out    std_logic_vector(0 downto 0);
        bisterr    :    out    std_logic_vector(0 downto 0);
        clk2b    :    out    std_logic_vector(0 downto 0);
        rcvdclkpmab    :    out    std_logic_vector(0 downto 0);
        syncstatus    :    out    std_logic_vector(0 downto 0);
        decoderdatavalid    :    out    std_logic_vector(0 downto 0);
        decoderdata    :    out    std_logic_vector(7 downto 0);
        decoderctrl    :    out    std_logic_vector(0 downto 0);
        runningdisparity    :    out    std_logic_vector(1 downto 0);
        selftestdone    :    out    std_logic_vector(0 downto 0);
        selftesterr    :    out    std_logic_vector(0 downto 0);
        errdata    :    out    std_logic_vector(15 downto 0);
        errctrl    :    out    std_logic_vector(1 downto 0);
        prbsdone    :    out    std_logic_vector(0 downto 0);
        prbserrlt    :    out    std_logic_vector(0 downto 0);
        signaldetectout    :    out    std_logic_vector(0 downto 0);
        aligndetsync    :    out    std_logic_vector(1 downto 0);
        rdalign    :    out    std_logic_vector(1 downto 0);
        bistdone    :    out    std_logic_vector(0 downto 0);
        runlengthviolation    :    out    std_logic_vector(0 downto 0);
        rlvlt    :    out    std_logic_vector(0 downto 0);
        rmfifopartialfull    :    out    std_logic_vector(0 downto 0);
        rmfifofull    :    out    std_logic_vector(0 downto 0);
        rmfifopartialempty    :    out    std_logic_vector(0 downto 0);
        rmfifoempty    :    out    std_logic_vector(0 downto 0);
        pcfifofull    :    out    std_logic_vector(0 downto 0);
        pcfifoempty    :    out    std_logic_vector(0 downto 0);
        a1a2k1k2flag    :    out    std_logic_vector(3 downto 0);
        byteordflag    :    out    std_logic_vector(0 downto 0);
        rxpipeclk    :    out    std_logic_vector(0 downto 0);
        channeltestbusout    :    out    std_logic_vector(9 downto 0);
        rxpipesoftreset    :    out    std_logic_vector(0 downto 0);
        phystatus    :    out    std_logic_vector(0 downto 0);
        rxvalid    :    out    std_logic_vector(0 downto 0);
        rxstatus    :    out    std_logic_vector(2 downto 0);
        pipedata    :    out    std_logic_vector(63 downto 0);
        rxdatavalid    :    out    std_logic_vector(3 downto 0);
        rxblkstart    :    out    std_logic_vector(3 downto 0);
        rxsynchdr    :    out    std_logic_vector(1 downto 0);
        speedchange    :    out    std_logic_vector(0 downto 0);
        eidledetected    :    out    std_logic_vector(0 downto 0);
        wordalignboundary    :    out    std_logic_vector(4 downto 0);
        rxclkslip    :    out    std_logic_vector(0 downto 0);
        eidleexit    :    out    std_logic_vector(0 downto 0);
        earlyeios    :    out    std_logic_vector(0 downto 0);
        ltr    :    out    std_logic_vector(0 downto 0);
        pcswrapbackin    :    in    std_logic_vector(69 downto 0);
        rxdivsyncinchnlup    :    in    std_logic_vector(1 downto 0);
        rxdivsyncinchnldown    :    in    std_logic_vector(1 downto 0);
        wrenableinchnlup    :    in    std_logic_vector(0 downto 0);
        wrenableinchnldown    :    in    std_logic_vector(0 downto 0);
        rdenableinchnlup    :    in    std_logic_vector(0 downto 0);
        rdenableinchnldown    :    in    std_logic_vector(0 downto 0);
        rxweinchnlup    :    in    std_logic_vector(1 downto 0);
        rxweinchnldown    :    in    std_logic_vector(1 downto 0);
        resetpcptrsinchnlup    :    in    std_logic_vector(0 downto 0);
        resetpcptrsinchnldown    :    in    std_logic_vector(0 downto 0);
        configselinchnlup    :    in    std_logic_vector(0 downto 0);
        configselinchnldown    :    in    std_logic_vector(0 downto 0);
        speedchangeinchnlup    :    in    std_logic_vector(0 downto 0);
        speedchangeinchnldown    :    in    std_logic_vector(0 downto 0);
        pcieswitch    :    out    std_logic_vector(0 downto 0);
        rxdivsyncoutchnlup    :    out    std_logic_vector(1 downto 0);
        rxweoutchnlup    :    out    std_logic_vector(1 downto 0);
        wrenableoutchnlup    :    out    std_logic_vector(0 downto 0);
        rdenableoutchnlup    :    out    std_logic_vector(0 downto 0);
        resetpcptrsoutchnlup    :    out    std_logic_vector(0 downto 0);
        speedchangeoutchnlup    :    out    std_logic_vector(0 downto 0);
        configseloutchnlup    :    out    std_logic_vector(0 downto 0);
        rxdivsyncoutchnldown    :    out    std_logic_vector(1 downto 0);
        rxweoutchnldown    :    out    std_logic_vector(1 downto 0);
        wrenableoutchnldown    :    out    std_logic_vector(0 downto 0);
        rdenableoutchnldown    :    out    std_logic_vector(0 downto 0);
        resetpcptrsoutchnldown    :    out    std_logic_vector(0 downto 0);
        speedchangeoutchnldown    :    out    std_logic_vector(0 downto 0);
        configseloutchnldown    :    out    std_logic_vector(0 downto 0);
        resetpcptrsinchnluppipe    :    out    std_logic_vector(0 downto 0);
        resetpcptrsinchnldownpipe    :    out    std_logic_vector(0 downto 0);
        speedchangeinchnluppipe    :    out    std_logic_vector(0 downto 0);
        speedchangeinchnldownpipe    :    out    std_logic_vector(0 downto 0);
        disablepcfifobyteserdes    :    out    std_logic_vector(0 downto 0);
        resetpcptrs    :    out    std_logic_vector(0 downto 0);
        rcvdclkagg    :    in    std_logic_vector(0 downto 0);
        rcvdclkaggtoporbot    :    in    std_logic_vector(0 downto 0);
        dispcbytegen3    :    in    std_logic_vector(0 downto 0);
        refclkdig    :    in    std_logic_vector(0 downto 0);
        txfifordclkraw    :    in    std_logic_vector(0 downto 0);
        resetpcptrsgen3    :    in    std_logic_vector(0 downto 0);
        syncdatain    :    out    std_logic_vector(0 downto 0);
        observablebyteserdesclock    :    out    std_logic_vector(0 downto 0)
    );
end component; --stratixv_hssi_8g_rx_pcs


component    stratixv_hssi_8g_tx_pcs
    generic    (
        prot_mode    :    string    :=    "basic";
        hip_mode    :    string    :=    "dis_hip";
        pma_dw    :    string    :=    "eight_bit";
        pcs_bypass    :    string    :=    "dis_pcs_bypass";
        phase_compensation_fifo    :    string    :=    "low_latency";
        tx_compliance_controlled_disparity    :    string    :=    "dis_txcompliance";
        force_kchar    :    string    :=    "dis_force_kchar";
        force_echar    :    string    :=    "dis_force_echar";
        byte_serializer    :    string    :=    "dis_bs";
        data_selection_8b10b_encoder_input    :    string    :=    "normal_data_path";
        eightb_tenb_disp_ctrl    :    string    :=    "dis_disp_ctrl";
        eightb_tenb_encoder    :    string    :=    "dis_8b10b";
        prbs_gen    :    string    :=    "dis_prbs";
        cid_pattern    :    string    :=    "cid_pattern_0";
        cid_pattern_len    :    bit_vector    :=    B"00000000";
        bist_gen    :    string    :=    "dis_bist";
        bit_reversal    :    string    :=    "dis_bit_reversal";
        symbol_swap    :    string    :=    "dis_symbol_swap";
        polarity_inversion    :    string    :=    "dis_polinv";
        tx_bitslip    :    string    :=    "dis_tx_bitslip";
        agg_block_sel    :    string    :=    "same_smrt_pack";
        revloop_back_rm    :    string    :=    "dis_rev_loopback_rx_rm";
        phfifo_write_clk_sel    :    string    :=    "pld_tx_clk";
        ctrl_plane_bonding_consumption    :    string    :=    "individual";
        bypass_pipeline_reg    :    string    :=    "dis_bypass_pipeline";
        ctrl_plane_bonding_distribution    :    string    :=    "not_master_chnl_distr";
        test_mode    :    string    :=    "prbs";
        clock_gate_tx    :    string    :=    "dis_clk_gating";
        self_switch_dw_scaling    :    string    :=    "dis_self_switch_dw_scaling";
        ctrl_plane_bonding_compensation    :    string    :=    "dis_compensation";
        refclk_b_clk_sel    :    string    :=    "tx_pma_clock";
        auto_speed_nego_gen2    :    string    :=    "dis_auto_speed_nego_g2";
        auto_speed_nego_gen3    :    string    :=    "dis_auto_speed_nego_g3";
        channel_number    :    string    :=    "int"
    );
    port    (
        txpcsreset    :    in    std_logic_vector(0 downto 0);
        refclkdig    :    in    std_logic_vector(0 downto 0);
        scanmode    :    in    std_logic_vector(0 downto 0);
        datain    :    in    std_logic_vector(43 downto 0);
        coreclk    :    in    std_logic_vector(0 downto 0);
        invpol    :    in    std_logic_vector(0 downto 0);
        xgmdatain    :    in    std_logic_vector(7 downto 0);
        xgmctrl    :    in    std_logic_vector(0 downto 0);
        xgmdataintoporbottom    :    in    std_logic_vector(7 downto 0);
        xgmctrltoporbottom    :    in    std_logic_vector(0 downto 0);
        txpmalocalclk    :    in    std_logic_vector(0 downto 0);
        enrevparallellpbk    :    in    std_logic_vector(0 downto 0);
        revparallellpbkdata    :    in    std_logic_vector(19 downto 0);
        phfifowrenable    :    in    std_logic_vector(0 downto 0);
        phfiforddisable    :    in    std_logic_vector(0 downto 0);
        phfiforeset    :    in    std_logic_vector(0 downto 0);
        detectrxloopin    :    in    std_logic_vector(0 downto 0);
        powerdn    :    in    std_logic_vector(1 downto 0);
        pipeenrevparallellpbkin    :    in    std_logic_vector(0 downto 0);
        pipetxswing    :    in    std_logic_vector(0 downto 0);
        pipetxdeemph    :    in    std_logic_vector(0 downto 0);
        pipetxmargin    :    in    std_logic_vector(2 downto 0);
        rxpolarityin    :    in    std_logic_vector(0 downto 0);
        polinvrxin    :    in    std_logic_vector(0 downto 0);
        elecidleinfersel    :    in    std_logic_vector(2 downto 0);
        rateswitch    :    in    std_logic_vector(0 downto 0);
        rateswitchbundle    :    in    std_logic_vector(0 downto 0);
        prbscidenable    :    in    std_logic_vector(0 downto 0);
        bitslipboundaryselect    :    in    std_logic_vector(4 downto 0);
        phfifooverflow    :    out    std_logic_vector(0 downto 0);
        phfifounderflow    :    out    std_logic_vector(0 downto 0);
        clkout    :    out    std_logic_vector(0 downto 0);
        clkoutgen3    :    out    std_logic_vector(0 downto 0);
        xgmdataout    :    out    std_logic_vector(7 downto 0);
        xgmctrlenable    :    out    std_logic_vector(0 downto 0);
        dataout    :    out    std_logic_vector(19 downto 0);
        rdenablesync    :    out    std_logic_vector(0 downto 0);
        refclkb    :    out    std_logic_vector(0 downto 0);
        parallelfdbkout    :    out    std_logic_vector(19 downto 0);
        txpipeclk    :    out    std_logic_vector(0 downto 0);
        encodertestbus    :    out    std_logic_vector(9 downto 0);
        txctrltestbus    :    out    std_logic_vector(9 downto 0);
        txpipesoftreset    :    out    std_logic_vector(0 downto 0);
        txpipeelectidle    :    out    std_logic_vector(0 downto 0);
        detectrxloopout    :    out    std_logic_vector(0 downto 0);
        pipepowerdownout    :    out    std_logic_vector(1 downto 0);
        pipeenrevparallellpbkout    :    out    std_logic_vector(0 downto 0);
        phfifotxswing    :    out    std_logic_vector(0 downto 0);
        phfifotxdeemph    :    out    std_logic_vector(0 downto 0);
        phfifotxmargin    :    out    std_logic_vector(2 downto 0);
        txdataouttogen3    :    out    std_logic_vector(31 downto 0);
        txdatakouttogen3    :    out    std_logic_vector(3 downto 0);
        txdatavalidouttogen3    :    out    std_logic_vector(3 downto 0);
        txblkstartout    :    out    std_logic_vector(3 downto 0);
        txsynchdrout    :    out    std_logic_vector(1 downto 0);
        txcomplianceout    :    out    std_logic_vector(0 downto 0);
        txelecidleout    :    out    std_logic_vector(0 downto 0);
        rxpolarityout    :    out    std_logic_vector(0 downto 0);
        polinvrxout    :    out    std_logic_vector(0 downto 0);
        grayelecidleinferselout    :    out    std_logic_vector(2 downto 0);
        txdivsyncinchnlup    :    in    std_logic_vector(1 downto 0);
        txdivsyncinchnldown    :    in    std_logic_vector(1 downto 0);
        wrenableinchnlup    :    in    std_logic_vector(0 downto 0);
        wrenableinchnldown    :    in    std_logic_vector(0 downto 0);
        rdenableinchnlup    :    in    std_logic_vector(0 downto 0);
        rdenableinchnldown    :    in    std_logic_vector(0 downto 0);
        fifoselectinchnlup    :    in    std_logic_vector(1 downto 0);
        fifoselectinchnldown    :    in    std_logic_vector(1 downto 0);
        resetpcptrs    :    in    std_logic_vector(0 downto 0);
        resetpcptrsinchnlup    :    in    std_logic_vector(0 downto 0);
        resetpcptrsinchnldown    :    in    std_logic_vector(0 downto 0);
        dispcbyte    :    in    std_logic_vector(0 downto 0);
        txdivsyncoutchnlup    :    out    std_logic_vector(1 downto 0);
        txdivsyncoutchnldown    :    out    std_logic_vector(1 downto 0);
        rdenableoutchnlup    :    out    std_logic_vector(0 downto 0);
        rdenableoutchnldown    :    out    std_logic_vector(0 downto 0);
        wrenableoutchnlup    :    out    std_logic_vector(0 downto 0);
        wrenableoutchnldown    :    out    std_logic_vector(0 downto 0);
        fifoselectoutchnlup    :    out    std_logic_vector(1 downto 0);
        fifoselectoutchnldown    :    out    std_logic_vector(1 downto 0);
        txfifordclkraw    :    out    std_logic_vector(0 downto 0);
        syncdatain    :    out    std_logic_vector(0 downto 0);
        observablebyteserdesclock    :    out    std_logic_vector(0 downto 0)
    );
end component; --stratixv_hssi_8g_tx_pcs


component    stratixv_hssi_common_pcs_pma_interface
    generic    (
        lpm_type    :    string    :=    "stratixv_hssi_common_pcs_pma_interface";
        auto_speed_ena    :    string    :=    "dis_auto_speed_ena";
        force_freqdet    :    string    :=    "force_freqdet_dis";
        func_mode    :    string    :=    "disable";
        pcie_gen3_cap    :    string    :=    "non_pcie_gen3_cap";
        pipe_if_g3pcs    :    string    :=    "pipe_if_8gpcs";
        pma_if_dft_en    :    string    :=    "dft_dis";
        pma_if_dft_val    :    string    :=    "dft_0";
        ppm_cnt_rst    :    string    :=    "ppm_cnt_rst_dis";
        ppm_deassert_early    :    string    :=    "deassert_early_dis";
        ppm_gen1_2_cnt    :    string    :=    "cnt_32k";
        ppm_post_eidle_delay    :    string    :=    "cnt_200_cycles";
        ppmsel    :    string    :=    "ppmsel_default";
        prot_mode    :    string    :=    "disabled_prot_mode";
        refclk_dig_sel    :    string    :=    "refclk_dig_dis";
        selectpcs    :    string    :=    "eight_g_pcs";
        sup_mode    :    string    :=    "full_mode"
    );
    port    (
        fref    :    in    std_logic;
        clklow    :    in    std_logic;
        pmapcieswdone    :    in    std_logic_vector(1 downto 0);
        pmarxfound    :    in    std_logic;
        pmarxdetectvalid    :    in    std_logic;
        pmahclk    :    in    std_logic;
        pldoffcalen    :    in    std_logic;
        aggrcvdclkagg    :    in    std_logic;
        aggtxdatats    :    in    std_logic_vector(7 downto 0);
        aggtxctlts    :    in    std_logic;
        aggfiforstrdqd    :    in    std_logic;
        aggendskwqd    :    in    std_logic;
        aggendskwrdptrs    :    in    std_logic;
        aggalignstatus    :    in    std_logic;
        aggalignstatussync0    :    in    std_logic;
        aggcgcomprddall    :    in    std_logic;
        aggcgcompwrall    :    in    std_logic;
        aggfifordincomp0    :    in    std_logic;
        aggdelcondmet0    :    in    std_logic;
        agginsertincomplete0    :    in    std_logic;
        aggfifoovr0    :    in    std_logic;
        agglatencycomp0    :    in    std_logic;
        aggrxdatars    :    in    std_logic_vector(7 downto 0);
        aggrxcontrolrs    :    in    std_logic;
        aggrcvdclkaggtoporbot    :    in    std_logic;
        aggtxdatatstoporbot    :    in    std_logic_vector(7 downto 0);
        aggtxctltstoporbot    :    in    std_logic;
        aggfiforstrdqdtoporbot    :    in    std_logic;
        aggendskwqdtoporbot    :    in    std_logic;
        aggendskwrdptrstoporbot    :    in    std_logic;
        aggalignstatustoporbot    :    in    std_logic;
        aggalignstatussync0toporbot    :    in    std_logic;
        aggcgcomprddalltoporbot    :    in    std_logic;
        aggcgcompwralltoporbot    :    in    std_logic;
        aggfifordincomp0toporbot    :    in    std_logic;
        aggdelcondmet0toporbot    :    in    std_logic;
        agginsertincomplete0toporbot    :    in    std_logic;
        aggfifoovr0toporbot    :    in    std_logic;
        agglatencycomp0toporbot    :    in    std_logic;
        aggrxdatarstoporbot    :    in    std_logic_vector(7 downto 0);
        aggrxcontrolrstoporbot    :    in    std_logic;
        pcsgen3pmapcieswitch    :    in    std_logic_vector(1 downto 0);
        pcsgen3pmatxmargin    :    in    std_logic_vector(2 downto 0);
        pcsgen3pmatxdeemph    :    in    std_logic;
        pcsgen3pmatxswing    :    in    std_logic;
        pcsgen3pmacurrentcoeff    :    in    std_logic_vector(17 downto 0);
        pcsgen3pmacurrentrxpreset    :    in    std_logic_vector(2 downto 0);
        pcsgen3pmatxelecidle    :    in    std_logic;
        pcsgen3pmatxdetectrx    :    in    std_logic;
        pcsgen3ppmeidleexit    :    in    std_logic;
        pcsgen3pmaltr    :    in    std_logic;
        pcsgen3pmaearlyeios    :    in    std_logic;
        pcs8gpcieswitch    :    in    std_logic;
        pcs8gtxelecidle    :    in    std_logic;
        pcs8gtxdetectrx    :    in    std_logic;
        pcs8gearlyeios    :    in    std_logic;
        pcs8gtxdeemphpma    :    in    std_logic;
        pcs8gtxmarginpma    :    in    std_logic_vector(2 downto 0);
        pcs8gtxswingpma    :    in    std_logic;
        pcs8gltrpma    :    in    std_logic;
        pcs8geidleexit    :    in    std_logic;
        pcsaggtxpcsrst    :    in    std_logic;
        pcsaggrxpcsrst    :    in    std_logic;
        pcsaggtxdatatc    :    in    std_logic_vector(7 downto 0);
        pcsaggtxctltc    :    in    std_logic;
        pcsaggrdenablesync    :    in    std_logic;
        pcsaggsyncstatus    :    in    std_logic;
        pcsaggaligndetsync    :    in    std_logic_vector(1 downto 0);
        pcsaggrdalign    :    in    std_logic_vector(1 downto 0);
        pcsaggalignstatussync    :    in    std_logic;
        pcsaggfifordoutcomp    :    in    std_logic;
        pcsaggcgcomprddout    :    in    std_logic_vector(1 downto 0);
        pcsaggcgcompwrout    :    in    std_logic_vector(1 downto 0);
        pcsaggdelcondmetout    :    in    std_logic;
        pcsaggfifoovrout    :    in    std_logic;
        pcsagglatencycompout    :    in    std_logic;
        pcsagginsertincompleteout    :    in    std_logic;
        pcsaggdecdatavalid    :    in    std_logic;
        pcsaggdecdata    :    in    std_logic_vector(7 downto 0);
        pcsaggdecctl    :    in    std_logic;
        pcsaggrunningdisp    :    in    std_logic_vector(1 downto 0);
        pldrxclkslip    :    in    std_logic;
        pldhardreset    :    in    std_logic;
        pcsscanmoden    :    in    std_logic;
        pcsscanshiftn    :    in    std_logic;
        pcsrefclkdig    :    in    std_logic;
        pcsaggscanmoden    :    in    std_logic;
        pcsaggscanshiftn    :    in    std_logic;
        pcsaggrefclkdig    :    in    std_logic;
        pcsgen3gen3datasel    :    in    std_logic;
        pldlccmurstb    :    in    std_logic;
        pmaoffcaldonein    :    in    std_logic;
        pmarxpmarstb    :    in    std_logic;
        pmahardreset    :    out    std_logic;
        freqlock    :    out    std_logic;
        pmapcieswitch    :    out    std_logic_vector(1 downto 0);
        pmaearlyeios    :    out    std_logic;
        pmatxdetectrx    :    out    std_logic;
        pmatxelecidle    :    out    std_logic;
        pmatxdeemph    :    out    std_logic;
        pmatxswing    :    out    std_logic;
        pmatxmargin    :    out    std_logic_vector(2 downto 0);
        pmacurrentcoeff    :    out    std_logic_vector(17 downto 0);
        pmacurrentrxpreset    :    out    std_logic_vector(2 downto 0);
        pmaoffcaldoneout    :    out    std_logic;
        pmalccmurstb    :    out    std_logic;
        pmaltr    :    out    std_logic;
        aggtxpcsrst    :    out    std_logic;
        aggrxpcsrst    :    out    std_logic;
        aggtxdatatc    :    out    std_logic_vector(7 downto 0);
        aggtxctltc    :    out    std_logic;
        aggrdenablesync    :    out    std_logic;
        aggsyncstatus    :    out    std_logic;
        aggaligndetsync    :    out    std_logic_vector(1 downto 0);
        aggrdalign    :    out    std_logic_vector(1 downto 0);
        aggalignstatussync    :    out    std_logic;
        aggfifordoutcomp    :    out    std_logic;
        aggcgcomprddout    :    out    std_logic_vector(1 downto 0);
        aggcgcompwrout    :    out    std_logic_vector(1 downto 0);
        aggdelcondmetout    :    out    std_logic;
        aggfifoovrout    :    out    std_logic;
        agglatencycompout    :    out    std_logic;
        agginsertincompleteout    :    out    std_logic;
        aggdecdatavalid    :    out    std_logic;
        aggdecdata    :    out    std_logic_vector(7 downto 0);
        aggdecctl    :    out    std_logic;
        aggrunningdisp    :    out    std_logic_vector(1 downto 0);
        pcsgen3pmarxdetectvalid    :    out    std_logic;
        pcsgen3pmarxfound    :    out    std_logic;
        pcsgen3pmapcieswdone    :    out    std_logic_vector(1 downto 0);
        pcsgen3pllfixedclk    :    out    std_logic;
        pcsaggrcvdclkagg    :    out    std_logic;
        pcsaggtxdatats    :    out    std_logic_vector(7 downto 0);
        pcsaggtxctlts    :    out    std_logic;
        pcsaggfiforstrdqd    :    out    std_logic;
        pcsaggendskwqd    :    out    std_logic;
        pcsaggendskwrdptrs    :    out    std_logic;
        pcsaggalignstatus    :    out    std_logic;
        pcsaggalignstatussync0    :    out    std_logic;
        pcsaggcgcomprddall    :    out    std_logic;
        pcsaggcgcompwrall    :    out    std_logic;
        pcsaggfifordincomp0    :    out    std_logic;
        pcsaggdelcondmet0    :    out    std_logic;
        pcsagginsertincomplete0    :    out    std_logic;
        pcsaggfifoovr0    :    out    std_logic;
        pcsagglatencycomp0    :    out    std_logic;
        pcsaggrxdatars    :    out    std_logic_vector(7 downto 0);
        pcsaggrxcontrolrs    :    out    std_logic;
        pcsaggrcvdclkaggtoporbot    :    out    std_logic;
        pcsaggtxdatatstoporbot    :    out    std_logic_vector(7 downto 0);
        pcsaggtxctltstoporbot    :    out    std_logic;
        pcsaggfiforstrdqdtoporbot    :    out    std_logic;
        pcsaggendskwqdtoporbot    :    out    std_logic;
        pcsaggendskwrdptrstoporbot    :    out    std_logic;
        pcsaggalignstatustoporbot    :    out    std_logic;
        pcsaggalignstatussync0toporbot    :    out    std_logic;
        pcsaggcgcomprddalltoporbot    :    out    std_logic;
        pcsaggcgcompwralltoporbot    :    out    std_logic;
        pcsaggfifordincomp0toporbot    :    out    std_logic;
        pcsaggdelcondmet0toporbot    :    out    std_logic;
        pcsagginsertincomplete0toporbot    :    out    std_logic;
        pcsaggfifoovr0toporbot    :    out    std_logic;
        pcsagglatencycomp0toporbot    :    out    std_logic;
        pcsaggrxdatarstoporbot    :    out    std_logic_vector(7 downto 0);
        pcsaggrxcontrolrstoporbot    :    out    std_logic;
        pcs8grxdetectvalid    :    out    std_logic;
        pcs8gpmarxfound    :    out    std_logic;
        pcs8ggen2ngen1    :    out    std_logic;
        pcs8gpowerstatetransitiondone    :    out    std_logic;
        ppmcntlatch    :    out    std_logic_vector(7 downto 0);
        pldhclkout    :    out    std_logic;
        aggscanmoden    :    out    std_logic;
        aggscanshiftn    :    out    std_logic;
        aggrefclkdig    :    out    std_logic;
        pmaoffcalen    :    out    std_logic;
        pmafrefout    :    out    std_logic;
        pmaclklowout    :    out    std_logic
    );
end component; --stratixv_hssi_common_pcs_pma_interface


component    stratixv_hssi_common_pld_pcs_interface
    generic    (
        lpm_type    :    string    :=    "stratixv_hssi_common_pld_pcs_interface";
        data_source    :    string    :=    "pld";
        emsip_enable    :    string    :=    "emsip_disable";
        selectpcs    :    string    :=    "eight_g_pcs"
    );
    port    (
        pldhardresetin    :    in    std_logic;
        pldscanmoden    :    in    std_logic;
        pldscanshiftn    :    in    std_logic;
        pldgen3refclkdig    :    in    std_logic;
        pld10grefclkdig    :    in    std_logic;
        pld8grefclkdig    :    in    std_logic;
        pldaggrefclkdig    :    in    std_logic;
        pldpcspmaifrefclkdig    :    in    std_logic;
        pldrate    :    in    std_logic_vector(1 downto 0);
        pldeidleinfersel    :    in    std_logic_vector(2 downto 0);
        pld8gsoftresetallhssi    :    in    std_logic;
        pld8gplniotri    :    in    std_logic;
        pld8gprbsciden    :    in    std_logic;
        pld8gltr    :    in    std_logic;
        pld8gtxelecidle    :    in    std_logic;
        pld8gtxdetectrxloopback    :    in    std_logic;
        pld8gtxdeemph    :    in    std_logic;
        pld8gtxmargin    :    in    std_logic_vector(2 downto 0);
        pld8gtxswing    :    in    std_logic;
        pld8grxpolarity    :    in    std_logic;
        pld8gpowerdown    :    in    std_logic_vector(1 downto 0);
        pldgen3currentcoeff    :    in    std_logic_vector(17 downto 0);
        pldgen3currentrxpreset    :    in    std_logic_vector(2 downto 0);
        pcs10gtestdata    :    in    std_logic_vector(19 downto 0);
        pcs8gchnltestbusout    :    in    std_logic_vector(9 downto 0);
        pcs8grxvalid    :    in    std_logic;
        pcs8grxelecidle    :    in    std_logic;
        pcs8grxstatus    :    in    std_logic_vector(2 downto 0);
        pcs8gphystatus    :    in    std_logic;
        pldhclkin    :    in    std_logic;
        pcsgen3pldasyncstatus    :    in    std_logic_vector(5 downto 0);
        pcsgen3testout    :    in    std_logic_vector(19 downto 0);
        emsippcsreset    :    in    std_logic_vector(2 downto 0);
        emsippcsctrl    :    in    std_logic_vector(38 downto 0);
        pmafref    :    in    std_logic;
        pmaclklow    :    in    std_logic;
        pmaoffcaldone    :    in    std_logic;
        pldoffcalenin    :    in    std_logic;
        pcsgen3masktxpll    :    in    std_logic;
        rcomemsip    :    in    std_logic;
        rcomhipena    :    in    std_logic;
        rcomblocksel    :    in    std_logic_vector(1 downto 0);
        pldtestdata    :    out    std_logic_vector(19 downto 0);
        pld8grxvalid    :    out    std_logic;
        pld8grxelecidle    :    out    std_logic;
        pld8grxstatus    :    out    std_logic_vector(2 downto 0);
        pld8gphystatus    :    out    std_logic;
        pldgen3pldasyncstatus    :    out    std_logic_vector(5 downto 0);
        pcs10ghardresetn    :    out    std_logic;
        pcs10gscanmoden    :    out    std_logic;
        pcs10gscanshiftn    :    out    std_logic;
        pcs10grefclkdig    :    out    std_logic;
        pcs8ghardreset    :    out    std_logic;
        pcs8gsoftresetallhssi    :    out    std_logic;
        pcs8gplniotri    :    out    std_logic;
        pcs8gscanmoden    :    out    std_logic;
        pcs8gscanshiftn    :    out    std_logic;
        pcs8grefclkdig    :    out    std_logic;
        pcs8gprbsciden    :    out    std_logic;
        pcs8gltr    :    out    std_logic;
        pcs8gtxelecidle    :    out    std_logic;
        pcs8gtxdetectrxloopback    :    out    std_logic;
        pcs8gtxdeemph    :    out    std_logic;
        pcs8gtxmargin    :    out    std_logic_vector(2 downto 0);
        pcs8gtxswing    :    out    std_logic;
        pcs8grxpolarity    :    out    std_logic;
        pcs8grate    :    out    std_logic;
        pcs8gpowerdown    :    out    std_logic_vector(1 downto 0);
        pcs8geidleinfersel    :    out    std_logic_vector(2 downto 0);
        pcsgen3pcsdigclk    :    out    std_logic;
        pcsgen3rate    :    out    std_logic_vector(1 downto 0);
        pcsgen3eidleinfersel    :    out    std_logic_vector(2 downto 0);
        pcsgen3scanmoden    :    out    std_logic;
        pcsgen3scanshiftn    :    out    std_logic;
        pcsgen3pldltr    :    out    std_logic;
        pldhardresetout    :    out    std_logic;
        pcsgen3currentcoeff    :    out    std_logic_vector(17 downto 0);
        pcsgen3currentrxpreset    :    out    std_logic_vector(2 downto 0);
        pcsaggrefclkdig    :    out    std_logic;
        pcspcspmaifrefclkdig    :    out    std_logic;
        pcsaggscanmoden    :    out    std_logic;
        pcsaggscanshiftn    :    out    std_logic;
        pcspcspmaifscanmoden    :    out    std_logic;
        pcspcspmaifscanshiftn    :    out    std_logic;
        emsippcsclkout    :    out    std_logic_vector(2 downto 0);
        emsippcsstatus    :    out    std_logic_vector(13 downto 0);
        pldfref    :    out    std_logic;
        pldclklow    :    out    std_logic;
        emsipenabledusermode    :    out    std_logic;
        pldoffcalenout    :    out    std_logic;
        pldoffcaldone    :    out    std_logic;
        pldgen3masktxpll    :    out    std_logic
    );
end component; --stratixv_hssi_common_pld_pcs_interface


component    stratixv_hssi_pipe_gen1_2
    generic    (
        prot_mode    :    string    :=    "pipe_g1";
        hip_mode    :    string    :=    "dis_hip";
        tx_pipe_enable    :    string    :=    "dis_pipe_tx";
        rx_pipe_enable    :    string    :=    "dis_pipe_rx";
        pipe_byte_de_serializer_en    :    string    :=    "dont_care_bds";
        txswing    :    string    :=    "dis_txswing";
        rxdetect_bypass    :    string    :=    "dis_rxdetect_bypass";
        error_replace_pad    :    string    :=    "replace_edb";
        ind_error_reporting    :    string    :=    "dis_ind_error_reporting";
        phystatus_rst_toggle    :    string    :=    "dis_phystatus_rst_toggle";
        elecidle_delay    :    string    :=    "elec_idle_delay";
        elec_idle_delay_val    :    bit_vector    :=    B"000";
        phy_status_delay    :    string    :=    "phystatus_delay";
        phystatus_delay_val    :    bit_vector    :=    B"000";
        ctrl_plane_bonding_consumption    :    string    :=    "individual";
        byte_deserializer    :    string    :=    "dis_bds"
    );
    port    (
        pipetxclk    :    in    std_logic_vector(0 downto 0);
        piperxclk    :    in    std_logic_vector(0 downto 0);
        refclkb    :    in    std_logic_vector(0 downto 0);
        txpipereset    :    in    std_logic_vector(0 downto 0);
        rxpipereset    :    in    std_logic_vector(0 downto 0);
        refclkbreset    :    in    std_logic_vector(0 downto 0);
        rrdwidthrx    :    in    std_logic_vector(0 downto 0);
        txdetectrxloopback    :    in    std_logic_vector(0 downto 0);
        txelecidlein    :    in    std_logic_vector(0 downto 0);
        powerdown    :    in    std_logic_vector(1 downto 0);
        txdeemph    :    in    std_logic_vector(0 downto 0);
        txmargin    :    in    std_logic_vector(2 downto 0);
        txswingport    :    in    std_logic_vector(0 downto 0);
        txdch    :    in    std_logic_vector(43 downto 0);
        rxpolarity    :    in    std_logic_vector(0 downto 0);
        sigdetni    :    in    std_logic_vector(0 downto 0);
        rxvalid    :    out    std_logic_vector(0 downto 0);
        rxelecidle    :    out    std_logic_vector(0 downto 0);
        rxstatus    :    out    std_logic_vector(2 downto 0);
        rxdch    :    out    std_logic_vector(63 downto 0);
        phystatus    :    out    std_logic_vector(0 downto 0);
        revloopback    :    in    std_logic_vector(0 downto 0);
        polinvrx    :    in    std_logic_vector(0 downto 0);
        txd    :    out    std_logic_vector(43 downto 0);
        revloopbk    :    out    std_logic_vector(0 downto 0);
        revloopbkpcsgen3    :    in    std_logic_vector(0 downto 0);
        rxelectricalidlepcsgen3    :    in    std_logic_vector(0 downto 0);
        txelecidlecomp    :    in    std_logic_vector(0 downto 0);
        rindvrx    :    in    std_logic_vector(0 downto 0);
        rmasterrx    :    in    std_logic_vector(1 downto 0);
        speedchange    :    in    std_logic_vector(0 downto 0);
        speedchangechnlup    :    in    std_logic_vector(0 downto 0);
        speedchangechnldown    :    in    std_logic_vector(0 downto 0);
        rxd    :    in    std_logic_vector(63 downto 0);
        txelecidleout    :    out    std_logic_vector(0 downto 0);
        txdetectrx    :    out    std_logic_vector(0 downto 0);
        powerstate    :    out    std_logic_vector(3 downto 0);
        rxfound    :    in    std_logic_vector(0 downto 0);
        rxdetectvalid    :    in    std_logic_vector(0 downto 0);
        rxelectricalidle    :    in    std_logic_vector(0 downto 0);
        powerstatetransitiondone    :    in    std_logic_vector(0 downto 0);
        powerstatetransitiondoneena    :    in    std_logic_vector(0 downto 0);
        txdeemphint    :    out    std_logic_vector(0 downto 0);
        txmarginint    :    out    std_logic_vector(2 downto 0);
        txswingint    :    out    std_logic_vector(0 downto 0);
        rxelectricalidleout    :    out    std_logic_vector(0 downto 0);
        rxpolaritypcsgen3    :    in    std_logic_vector(0 downto 0);
        polinvrxint    :    out    std_logic_vector(0 downto 0);
        speedchangeout    :    out    std_logic_vector(0 downto 0)
    );
end component; --stratixv_hssi_pipe_gen1_2


component    stratixv_hssi_pipe_gen3
    generic    (
        mode    :    string    :=    "pipe_g1";
        ctrl_plane_bonding    :    string    :=    "individual";
        pipe_clk_sel    :    string    :=    "func_clk";
        rate_match_pad_insertion    :    string    :=    "dis_rm_fifo_pad_ins";
        ind_error_reporting    :    string    :=    "dis_ind_error_reporting";
        phystatus_rst_toggle_g3    :    string    :=    "dis_phystatus_rst_toggle_g3";
        phystatus_rst_toggle_g12    :    string    :=    "dis_phystatus_rst_toggle";
        cdr_control    :    string    :=    "en_cdr_ctrl";
        cid_enable    :    string    :=    "en_cid_mode";
        parity_chk_ts1    :    string    :=    "en_ts1_parity_chk";
        rxvalid_mask    :    string    :=    "rxvalid_mask_en";
        ph_fifo_reg_mode    :    string    :=    "phfifo_reg_mode_dis";
        test_mode_timers    :    string    :=    "dis_test_mode_timers";
        inf_ei_enable    :    string    :=    "dis_inf_ei";
        spd_chnge_g2_sel    :    string    :=    "false";
        cp_up_mstr    :    string    :=    "false";
        cp_dwn_mstr    :    string    :=    "false";
        cp_cons_sel    :    string    :=    "cp_cons_default";
        elecidle_delay_g12_data    :    bit_vector    :=    B"000";
        elecidle_delay_g12    :    string    :=    "elecidle_delay_g12";
        elecidle_delay_g3_data    :    bit_vector    :=    B"000";
        elecidle_delay_g3    :    string    :=    "elecidle_delay_g3";
        phy_status_delay_g12_data    :    bit_vector    :=    B"000";
        phy_status_delay_g12    :    string    :=    "phy_status_delay_g12";
        phy_status_delay_g3_data    :    bit_vector    :=    B"000";
        phy_status_delay_g3    :    string    :=    "phy_status_delay_g3";
        sigdet_wait_counter_data    :    bit_vector    :=    B"00000000";
        sigdet_wait_counter    :    string    :=    "sigdet_wait_counter";
        data_mask_count_val    :    bit_vector    :=    B"0000000000";
        data_mask_count    :    string    :=    "data_mask_count";
        pma_done_counter_data    :    bit_vector    :=    B"000000000000000000";
        pma_done_counter    :    string    :=    "pma_done_count";
        pc_en_counter_data    :    bit_vector    :=    B"00000";
        pc_en_counter    :    string    :=    "pc_en_count";
        pc_rst_counter_data    :    bit_vector    :=    B"0000";
        pc_rst_counter    :    string    :=    "pc_rst_count";
        phfifo_flush_wait_data    :    bit_vector    :=    B"000000";
        phfifo_flush_wait    :    string    :=    "phfifo_flush_wait";
        asn_clk_enable    :    string    :=    "false";
        free_run_clk_enable    :    string    :=    "true";
        asn_enable    :    string    :=    "dis_asn"
    );
    port    (
        rcvdclk    :    in    std_logic_vector(0 downto 0);
        txpmaclk    :    in    std_logic_vector(0 downto 0);
        pcsdigclk    :    in    std_logic_vector(0 downto 0);
        pllfixedclk    :    in    std_logic_vector(0 downto 0);
        rtxgen3capen    :    in    std_logic_vector(0 downto 0);
        rrxgen3capen    :    in    std_logic_vector(0 downto 0);
        rtxdigclksel    :    in    std_logic_vector(0 downto 0);
        rrxdigclksel    :    in    std_logic_vector(0 downto 0);
        rxrstn    :    in    std_logic_vector(0 downto 0);
        txrstn    :    in    std_logic_vector(0 downto 0);
        scanmoden    :    in    std_logic_vector(0 downto 0);
        pldasyncstatus    :    out    std_logic_vector(5 downto 0);
        testout    :    out    std_logic_vector(19 downto 0);
        gen3datasel    :    out    std_logic_vector(0 downto 0);
        gen3clksel    :    out    std_logic_vector(0 downto 0);
        pcsrst    :    out    std_logic_vector(0 downto 0);
        dispcbyte    :    out    std_logic_vector(0 downto 0);
        resetpcprts    :    out    std_logic_vector(0 downto 0);
        shutdownclk    :    out    std_logic_vector(0 downto 0);
        txdata    :    in    std_logic_vector(31 downto 0);
        txdatak    :    in    std_logic_vector(3 downto 0);
        txdataskip    :    in    std_logic_vector(0 downto 0);
        txsynchdr    :    in    std_logic_vector(1 downto 0);
        txblkstart    :    in    std_logic_vector(0 downto 0);
        txelecidle    :    in    std_logic_vector(0 downto 0);
        txdetectrxloopback    :    in    std_logic_vector(0 downto 0);
        txcompliance    :    in    std_logic_vector(0 downto 0);
        rxpolarity    :    in    std_logic_vector(0 downto 0);
        powerdown    :    in    std_logic_vector(1 downto 0);
        rate    :    in    std_logic_vector(1 downto 0);
        txmargin    :    in    std_logic_vector(2 downto 0);
        txdeemph    :    in    std_logic_vector(0 downto 0);
        txswing    :    in    std_logic_vector(0 downto 0);
        eidleinfersel    :    in    std_logic_vector(2 downto 0);
        currentcoeff    :    in    std_logic_vector(17 downto 0);
        currentrxpreset    :    in    std_logic_vector(2 downto 0);
        rxupdatefc    :    in    std_logic_vector(0 downto 0);
        rxdataskip    :    out    std_logic_vector(3 downto 0);
        rxsynchdr    :    out    std_logic_vector(1 downto 0);
        rxblkstart    :    out    std_logic_vector(3 downto 0);
        rxvalid    :    out    std_logic_vector(0 downto 0);
        phystatus    :    out    std_logic_vector(0 downto 0);
        rxelecidle    :    out    std_logic_vector(0 downto 0);
        rxstatus    :    out    std_logic_vector(2 downto 0);
        rxdataint    :    in    std_logic_vector(31 downto 0);
        rxdatakint    :    in    std_logic_vector(3 downto 0);
        rxdataskipint    :    in    std_logic_vector(0 downto 0);
        rxsynchdrint    :    in    std_logic_vector(1 downto 0);
        rxblkstartint    :    in    std_logic_vector(0 downto 0);
        txdataint    :    out    std_logic_vector(31 downto 0);
        txdatakint    :    out    std_logic_vector(3 downto 0);
        txdataskipint    :    out    std_logic_vector(0 downto 0);
        txsynchdrint    :    out    std_logic_vector(1 downto 0);
        txblkstartint    :    out    std_logic_vector(0 downto 0);
        testinfei    :    out    std_logic_vector(18 downto 0);
        eidetint    :    in    std_logic_vector(0 downto 0);
        eipartialdetint    :    in    std_logic_vector(0 downto 0);
        idetint    :    in    std_logic_vector(0 downto 0);
        blkalgndint    :    in    std_logic_vector(0 downto 0);
        clkcompinsertint    :    in    std_logic_vector(0 downto 0);
        clkcompdeleteint    :    in    std_logic_vector(0 downto 0);
        clkcompoverflint    :    in    std_logic_vector(0 downto 0);
        clkcompundflint    :    in    std_logic_vector(0 downto 0);
        errdecodeint    :    in    std_logic_vector(0 downto 0);
        rcvlfsrchkint    :    in    std_logic_vector(0 downto 0);
        errencodeint    :    in    std_logic_vector(0 downto 0);
        rxpolarityint    :    out    std_logic_vector(0 downto 0);
        revlpbkint    :    out    std_logic_vector(0 downto 0);
        inferredrxvalidint    :    out    std_logic_vector(0 downto 0);
        rxd8gpcsin    :    in    std_logic_vector(63 downto 0);
        rxelecidle8gpcsin    :    in    std_logic_vector(0 downto 0);
        pldltr    :    in    std_logic_vector(0 downto 0);
        rxd8gpcsout    :    out    std_logic_vector(63 downto 0);
        revlpbk8gpcsout    :    out    std_logic_vector(0 downto 0);
        pmarxdetectvalid    :    in    std_logic_vector(0 downto 0);
        pmarxfound    :    in    std_logic_vector(0 downto 0);
        pmasignaldet    :    in    std_logic_vector(0 downto 0);
        pmapcieswdone    :    in    std_logic_vector(1 downto 0);
        pmapcieswitch    :    out    std_logic_vector(1 downto 0);
        pmatxmargin    :    out    std_logic_vector(2 downto 0);
        pmatxdeemph    :    out    std_logic_vector(0 downto 0);
        pmatxswing    :    out    std_logic_vector(0 downto 0);
        pmacurrentcoeff    :    out    std_logic_vector(17 downto 0);
        pmacurrentrxpreset    :    out    std_logic_vector(2 downto 0);
        pmatxelecidle    :    out    std_logic_vector(0 downto 0);
        pmatxdetectrx    :    out    std_logic_vector(0 downto 0);
        ppmeidleexit    :    out    std_logic_vector(0 downto 0);
        pmaltr    :    out    std_logic_vector(0 downto 0);
        pmaearlyeios    :    out    std_logic_vector(0 downto 0);
        pmarxdetpd    :    out    std_logic_vector(0 downto 0);
        bundlingindown    :    in    std_logic_vector(9 downto 0);
        bundlingoutdown    :    out    std_logic_vector(9 downto 0);
        rxpolarity8gpcsout    :    out    std_logic_vector(0 downto 0);
        speedchangeg2    :    in    std_logic_vector(0 downto 0);
        bundlingoutup    :    out    std_logic_vector(9 downto 0);
        bundlinginup    :    in    std_logic_vector(9 downto 0);
        masktxpll    :    out    std_logic_vector(0 downto 0)
    );
end component; --stratixv_hssi_pipe_gen3


component    stratixv_hssi_pma_cdr_refclk_select_mux
    generic    (
        lpm_type    :    string    :=    "stratixv_hssi_pma_cdr_refclk_select_mux";
        channel_number    :    integer    :=    0;
        refclk_select    :    string    :=    "ref_iqclk0";
        reference_clock_frequency    :    string    :=    "0 ps"
    );
    port    (
        calclk    :    in    std_logic;
        ffplloutbot    :    in    std_logic;
        ffpllouttop    :    in    std_logic;
        pldclk    :    in    std_logic;
        refiqclk0    :    in    std_logic;
        refiqclk1    :    in    std_logic;
        refiqclk10    :    in    std_logic;
        refiqclk2    :    in    std_logic;
        refiqclk3    :    in    std_logic;
        refiqclk4    :    in    std_logic;
        refiqclk5    :    in    std_logic;
        refiqclk6    :    in    std_logic;
        refiqclk7    :    in    std_logic;
        refiqclk8    :    in    std_logic;
        refiqclk9    :    in    std_logic;
        rxiqclk0    :    in    std_logic;
        rxiqclk1    :    in    std_logic;
        rxiqclk10    :    in    std_logic;
        rxiqclk2    :    in    std_logic;
        rxiqclk3    :    in    std_logic;
        rxiqclk4    :    in    std_logic;
        rxiqclk5    :    in    std_logic;
        rxiqclk6    :    in    std_logic;
        rxiqclk7    :    in    std_logic;
        rxiqclk8    :    in    std_logic;
        rxiqclk9    :    in    std_logic;
        clkout    :    out    std_logic
    );
end component; --stratixv_hssi_pma_cdr_refclk_select_mux


component    stratixv_hssi_pma_rx_buf
    generic    (
        lpm_type    :    string    :=    "stratixv_hssi_pma_rx_buf";
        adce_pd    :    string    :=    "false";
        bypass_eqz_stages_123    :    string    :=    "all_stages_enabled";
        eq_bw_sel    :    string    :=    "bw_full_12p5";
        input_vcm_sel    :    string    :=    "high_vcm";
        pdb_dfe    :    string    :=    "false";
        pdb_sd    :    string    :=    "false";
        qpi_enable    :    string    :=    "false";
        rx_dc_gain    :    string    :=    "dc_gain_0db";
        rx_sel_bias_source    :    string    :=    "bias_vcmdrv";
        sd_off    :    string    :=    "clk_divrx_2";
        sd_on    :    string    :=    "data_pulse_6";
        sd_threshold    :    string    :=    "sdlv_30mv";
        serial_loopback    :    string    :=    "lpbkp_dis";
        term_sel    :    string    :=    "r_100ohm";
        vccela_supply_voltage    :    string    :=    "vccela_1p0v";
        vcm_sel    :    string    :=    "vtt_0p7v";
        channel_number    :    integer    :=    0
    );
    port    (
        ck0sigdet    :    in    std_logic;
        datain    :    in    std_logic;
        fined2aout    :    in    std_logic;
        lpbkp    :    in    std_logic;
        occalen    :    in    std_logic;
        refclklpbk    :    in    std_logic;
        rstn    :    in    std_logic;
        rxqpipulldn    :    in    std_logic;
        slpbk    :    in    std_logic;
        dataout    :    out    std_logic;
        nonuserfrompmaux    :    out    std_logic;
        rdlpbkp    :    out    std_logic;
        rxpadce    :    out    std_logic;
        sd    :    out    std_logic
    );
end component; --stratixv_hssi_pma_rx_buf


component    stratixv_hssi_pma_rx_deser
    generic    (
        lpm_type    :    string    :=    "stratixv_hssi_pma_rx_deser";
        auto_negotiation    :    string    :=    "false";
        bit_slip_bypass    :    string    :=    "false";
        mode    :    integer    :=    8;
        sdclk_enable    :    string    :=    "false";
        vco_bypass    :    string    :=    "vco_bypass_normal";
        channel_number    :    integer    :=    0;
        clk_forward_only_mode    :    string    :=    "false"
    );
    port    (
        bslip    :    in    std_logic;
        clk90b    :    in    std_logic;
        clk270b    :    in    std_logic;
        deven    :    in    std_logic;
        dodd    :    in    std_logic;
        pciesw    :    in    std_logic_vector(1 downto 0);
        pfdmodelock    :    in    std_logic;
        rstn    :    in    std_logic;
        clk33pcs    :    out    std_logic;
        clkdivrx    :    out    std_logic;
        clkdivrxrx    :    out    std_logic;
        dout    :    out    std_logic_vector(39 downto 0);
        pciel    :    out    std_logic;
        pciem    :    out    std_logic
    );
end component; --stratixv_hssi_pma_rx_deser


component    stratixv_hssi_pma_tx_buf
    generic    (
        lpm_type    :    string    :=    "stratixv_hssi_pma_tx_buf";
        elec_idl_gate_ctrl    :    string    :=    "true";
        pre_emp_switching_ctrl_1st_post_tap    :    string    :=    "fir_1pt_disabled";
        pre_emp_switching_ctrl_2nd_post_tap    :    string    :=    "fir_2pt_disabled";
        pre_emp_switching_ctrl_pre_tap    :    string    :=    "fir_pre_disabled";
        qpi_en    :    string    :=    "false";
        rx_det    :    string    :=    "mode_0";
        rx_det_output_sel    :    string    :=    "rx_det_pcie_out";
        rx_det_pdb    :    string    :=    "true";
        sig_inv_2nd_tap    :    string    :=    "false";
        sig_inv_pre_tap    :    string    :=    "false";
        slew_rate_ctrl    :    string    :=    "slew_30ps";
        term_sel    :    string    :=    "r_100ohm";
        vod_switching_ctrl_main_tap    :    string    :=    "fir_main_2p0ma";
        channel_number    :    integer    :=    0
    );
    port    (
        datain    :    in    std_logic;
        rxdetclk    :    in    std_logic;
        txdetrx    :    in    std_logic;
        txelecidl    :    in    std_logic;
        txqpipulldn    :    in    std_logic;
        txqpipullup    :    in    std_logic;
        compass    :    out    std_logic;
        dataout    :    out    std_logic;
        detecton    :    out    std_logic_vector(1 downto 0);
        fixedclkout    :    out    std_logic;
        nonuserfrompmaux    :    out    std_logic;
        probepass    :    out    std_logic;
        rxdetectvalid    :    out    std_logic;
        rxfound    :    out    std_logic
    );
end component; --stratixv_hssi_pma_tx_buf


component    stratixv_hssi_pma_tx_cgb
    generic    (
        lpm_type    :    string    :=    "stratixv_hssi_pma_tx_cgb";
        auto_negotiation    :    string    :=    "false";
        x1_div_m_sel    :    integer    :=    1;
        channel_number    :    integer    :=    0;
        data_rate    :    string    :=    "";
        mode    :    integer    :=    8;
        rx_iqclk_sel    :    string    :=    "cgb_x1_n_div";
        tx_mux_power_down    :    string    :=    "normal";
        x1_clock_source_sel    :    string    :=    "x1_clk_unused";
        xn_clock_source_sel    :    string    :=    "cgb_xn_unused";
        xn_network_driver    :    string    :=    "enable_clock_entwork_driver";
        cgb_iqclk_sel    :    string    :=    "cgb_x1_n_div";
        ht_delay_enable    :    string    :=    "false"
    );
    port    (
        clkbcdr1adj    :    in    std_logic;
        clkbcdr1loc    :    in    std_logic;
        clkbcdrloc    :    in    std_logic;
        clkbdnseg    :    in    std_logic;
        clkbffpll    :    in    std_logic;
        clkblcb    :    in    std_logic;
        clkblct    :    in    std_logic;
        clkbupseg    :    in    std_logic;
        clkcdr1adj    :    in    std_logic;
        clkcdr1loc    :    in    std_logic;
        clkcdrloc    :    in    std_logic;
        clkdnseg    :    in    std_logic;
        clkffpll    :    in    std_logic;
        clklcb    :    in    std_logic;
        clklct    :    in    std_logic;
        clkupseg    :    in    std_logic;
        cpulsex6adj    :    in    std_logic;
        cpulsex6loc    :    in    std_logic;
        cpulsexndn    :    in    std_logic;
        cpulsexnup    :    in    std_logic;
        hfclknx6adj    :    in    std_logic;
        hfclknx6loc    :    in    std_logic;
        hfclknxndn    :    in    std_logic;
        hfclknxnup    :    in    std_logic;
        hfclkpx6adj    :    in    std_logic;
        hfclkpx6loc    :    in    std_logic;
        hfclkpxndn    :    in    std_logic;
        hfclkpxnup    :    in    std_logic;
        lfclknx6adj    :    in    std_logic;
        lfclknx6loc    :    in    std_logic;
        lfclknxndn    :    in    std_logic;
        lfclknxnup    :    in    std_logic;
        lfclkpx6adj    :    in    std_logic;
        lfclkpx6loc    :    in    std_logic;
        lfclkpxndn    :    in    std_logic;
        lfclkpxnup    :    in    std_logic;
        pciesw    :    in    std_logic_vector(1 downto 0);
        pclk0x6adj    :    in    std_logic;
        pclk0x6loc    :    in    std_logic;
        pclk0xndn    :    in    std_logic;
        pclk0xnup    :    in    std_logic;
        pclk1x6adj    :    in    std_logic;
        pclk1x6loc    :    in    std_logic;
        pclk1xndn    :    in    std_logic;
        pclk1xnup    :    in    std_logic;
        pclkx6adj    :    in    std_logic_vector(2 downto 0);
        pclkx6loc    :    in    std_logic_vector(2 downto 0);
        pclkxndn    :    in    std_logic_vector(2 downto 0);
        pclkxnup    :    in    std_logic_vector(2 downto 0);
        rxclk    :    in    std_logic;
        txpmarstb    :    in    std_logic;
        txpmasyncp    :    in    std_logic;
        xnresetin    :    in    std_logic;
        cpulse    :    out    std_logic;
        cpulseout    :    out    std_logic;
        hfclkn    :    out    std_logic;
        hfclknout    :    out    std_logic;
        hfclkp    :    out    std_logic;
        hfclkpout    :    out    std_logic;
        lfclkn    :    out    std_logic;
        lfclknout    :    out    std_logic;
        lfclkp    :    out    std_logic;
        lfclkpout    :    out    std_logic;
        pcieswdone    :    out    std_logic_vector(1 downto 0);
        pclk0    :    out    std_logic;
        pclk0out    :    out    std_logic;
        pclk1    :    out    std_logic;
        pclk1out    :    out    std_logic;
        pclk    :    out    std_logic_vector(2 downto 0);
        pclkout    :    out    std_logic_vector(2 downto 0);
        rxiqclk    :    out    std_logic;
        xnresetout    :    out    std_logic
    );
end component; --stratixv_hssi_pma_tx_cgb


component    stratixv_hssi_pma_tx_ser
    generic    (
        lpm_type    :    string    :=    "stratixv_hssi_pma_tx_ser";
        auto_negotiation    :    string    :=    "false";
        clk_divtx_deskew    :    string    :=    "deskew_delay1";
        mode    :    integer    :=    8;
        post_tap_1_en    :    string    :=    "false";
        post_tap_2_en    :    string    :=    "false";
        pre_tap_en    :    string    :=    "false";
        ser_loopback    :    string    :=    "false";
        pclksel    :    string    :=    "local_pclk";
        channel_number    :    integer    :=    0;
        clk_forward_only_mode    :    string    :=    "false"
    );
    port    (
        cpulse    :    in    std_logic;
        datain    :    in    std_logic_vector(39 downto 0);
        hfclk    :    in    std_logic;
        hfclkn    :    in    std_logic;
        lfclk    :    in    std_logic;
        lfclkn    :    in    std_logic;
        pciesw    :    in    std_logic_vector(1 downto 0);
        pclk0    :    in    std_logic;
        pclk1    :    in    std_logic;
        pclk2    :    in    std_logic;
        pclk    :    in    std_logic_vector(2 downto 0);
        rstn    :    in    std_logic;
        clkdivtx    :    out    std_logic;
        dataout    :    out    std_logic;
        div5    :    out    std_logic;
        lbvop    :    out    std_logic
    );
end component; --stratixv_hssi_pma_tx_ser


component    stratixv_hssi_rx_pcs_pma_interface
    generic    (
        lpm_type    :    string    :=    "stratixv_hssi_rx_pcs_pma_interface";
        clkslip_sel    :    string    :=    "pld";
        prot_mode    :    string    :=    "other_protocols";
        selectpcs    :    string    :=    "eight_g_pcs"
    );
    port    (
        clockinfrompma    :    in    std_logic;
        datainfrompma    :    in    std_logic_vector(39 downto 0);
        pmasigdet    :    in    std_logic;
        pmasignalok    :    in    std_logic;
        pcs10grxclkiqout    :    in    std_logic;
        pcsgen3rxclkiqout    :    in    std_logic;
        pcs8grxclkiqout    :    in    std_logic;
        pcs8grxclkslip    :    in    std_logic;
        pmaclkdiv33txorrxin    :    in    std_logic;
        pmarxplllockin    :    in    std_logic;
        pldrxpmarstb    :    in    std_logic;
        pldrxclkslip    :    in    std_logic;
        rrxblocksel    :    in    std_logic_vector(1 downto 0);
        rrxclkslipsel    :    in    std_logic;
        pmarxclkslip    :    out    std_logic;
        pmarxclkout    :    out    std_logic;
        clkoutto10gpcs    :    out    std_logic;
        dataoutto10gpcs    :    out    std_logic_vector(39 downto 0);
        pcs10gsignalok    :    out    std_logic;
        clockouttogen3pcs    :    out    std_logic;
        dataouttogen3pcs    :    out    std_logic_vector(31 downto 0);
        pcsgen3pmasignaldet    :    out    std_logic;
        clockoutto8gpcs    :    out    std_logic;
        dataoutto8gpcs    :    out    std_logic_vector(19 downto 0);
        pcs8gsigdetni    :    out    std_logic;
        pmaclkdiv33txorrxout    :    out    std_logic;
        pcs10gclkdiv33txorrx    :    out    std_logic;
        pmarxpmarstb    :    out    std_logic;
        pmarxplllockout    :    out    std_logic
    );
end component; --stratixv_hssi_rx_pcs_pma_interface


component    stratixv_hssi_rx_pld_pcs_interface
    generic    (
        lpm_type    :    string    :=    "stratixv_hssi_rx_pld_pcs_interface";
        data_source    :    string    :=    "pld";
        is_10g_0ppm    :    string    :=    "false";
        is_8g_0ppm    :    string    :=    "false";
        selectpcs    :    string    :=    "eight_g_pcs"
    );
    port    (
        pld10grxpldclk    :    in    std_logic;
        pld10grxpldrstn    :    in    std_logic;
        pld10grxalignen    :    in    std_logic;
        pld10grxalignclr    :    in    std_logic;
        pld10grxrden    :    in    std_logic;
        pld10grxdispclr    :    in    std_logic;
        pld10grxclrerrblkcnt    :    in    std_logic;
        pld10grxclrbercount    :    in    std_logic;
        pld10grxprbserrclr    :    in    std_logic;
        pld10grxbitslip    :    in    std_logic;
        pld8grxurstpma    :    in    std_logic;
        pld8grxurstpcs    :    in    std_logic;
        pld8gcmpfifourst    :    in    std_logic;
        pld8gphfifourstrx    :    in    std_logic;
        pld8gencdt    :    in    std_logic;
        pld8ga1a2size    :    in    std_logic;
        pld8gbitslip    :    in    std_logic;
        pld8grdenablermf    :    in    std_logic;
        pld8gwrenablermf    :    in    std_logic;
        pld8gpldrxclk    :    in    std_logic;
        pld8gpolinvrx    :    in    std_logic;
        pld8gbitlocreven    :    in    std_logic;
        pld8gbytereven    :    in    std_logic;
        pld8gbytordpld    :    in    std_logic;
        pld8gwrdisablerx    :    in    std_logic;
        pld8grdenablerx    :    in    std_logic;
        pldgen3rxrstn    :    in    std_logic;
        pldrxclkslipin    :    in    std_logic;
        pld8gpldextrain    :    in    std_logic_vector(3 downto 0);
        clockinfrom10gpcs    :    in    std_logic;
        pcs10grxdatavalid    :    in    std_logic;
        datainfrom10gpcs    :    in    std_logic_vector(63 downto 0);
        pcs10grxcontrol    :    in    std_logic_vector(9 downto 0);
        pcs10grxempty    :    in    std_logic;
        pcs10grxpempty    :    in    std_logic;
        pcs10grxpfull    :    in    std_logic;
        pcs10grxoflwerr    :    in    std_logic;
        pcs10grxalignval    :    in    std_logic;
        pcs10grxblklock    :    in    std_logic;
        pcs10grxhiber    :    in    std_logic;
        pcs10grxframelock    :    in    std_logic;
        pcs10grxrdpossts    :    in    std_logic;
        pcs10grxrdnegsts    :    in    std_logic;
        pcs10grxskipins    :    in    std_logic;
        pcs10grxrxframe    :    in    std_logic;
        pcs10grxpyldins    :    in    std_logic;
        pcs10grxsyncerr    :    in    std_logic;
        pcs10grxscrmerr    :    in    std_logic;
        pcs10grxskiperr    :    in    std_logic;
        pcs10grxdiagerr    :    in    std_logic;
        pcs10grxsherr    :    in    std_logic;
        pcs10grxmfrmerr    :    in    std_logic;
        pcs10grxcrc32err    :    in    std_logic;
        pcs10grxdiagstatus    :    in    std_logic_vector(1 downto 0);
        datainfrom8gpcs    :    in    std_logic_vector(63 downto 0);
        clockinfrom8gpcs    :    in    std_logic;
        pcs8gbisterr    :    in    std_logic;
        pcs8grcvdclkpmab    :    in    std_logic;
        pcs8gsignaldetectout    :    in    std_logic;
        pcs8gbistdone    :    in    std_logic;
        pcs8grlvlt    :    in    std_logic;
        pcs8gfullrmf    :    in    std_logic;
        pcs8gemptyrmf    :    in    std_logic;
        pcs8gfullrx    :    in    std_logic;
        pcs8gemptyrx    :    in    std_logic;
        pcs8ga1a2k1k2flag    :    in    std_logic_vector(3 downto 0);
        pcs8gbyteordflag    :    in    std_logic;
        pcs8gwaboundary    :    in    std_logic_vector(4 downto 0);
        pcs8grxdatavalid    :    in    std_logic_vector(3 downto 0);
        pcs8grxsynchdr    :    in    std_logic_vector(1 downto 0);
        pcs8grxblkstart    :    in    std_logic_vector(3 downto 0);
        pmaclkdiv33txorrx    :    in    std_logic;
        emsippcsrxclkin    :    in    std_logic_vector(2 downto 0);
        emsippcsrxreset    :    in    std_logic_vector(6 downto 0);
        emsippcsrxctrl    :    in    std_logic_vector(24 downto 0);
        pmarxplllock    :    in    std_logic;
        pldrxpmarstbin    :    in    std_logic;
        rrxblocksel    :    in    std_logic_vector(1 downto 0);
        rrxemsip    :    in    std_logic;
        emsipenabledusermode    :    in    std_logic;
        pcs10grxfifoinsert    :    in    std_logic;
        pld8gsyncsmeninput    :    in    std_logic;
        pcs10grxfifodel    :    in    std_logic;
        dataouttopld    :    out    std_logic_vector(63 downto 0);
        pld10grxclkout    :    out    std_logic;
        pld10grxdatavalid    :    out    std_logic;
        pld10grxcontrol    :    out    std_logic_vector(9 downto 0);
        pld10grxempty    :    out    std_logic;
        pld10grxpempty    :    out    std_logic;
        pld10grxpfull    :    out    std_logic;
        pld10grxoflwerr    :    out    std_logic;
        pld10grxalignval    :    out    std_logic;
        pld10grxblklock    :    out    std_logic;
        pld10grxhiber    :    out    std_logic;
        pld10grxframelock    :    out    std_logic;
        pld10grxrdpossts    :    out    std_logic;
        pld10grxrdnegsts    :    out    std_logic;
        pld10grxskipins    :    out    std_logic;
        pld10grxrxframe    :    out    std_logic;
        pld10grxpyldins    :    out    std_logic;
        pld10grxsyncerr    :    out    std_logic;
        pld10grxscrmerr    :    out    std_logic;
        pld10grxskiperr    :    out    std_logic;
        pld10grxdiagerr    :    out    std_logic;
        pld10grxsherr    :    out    std_logic;
        pld10grxmfrmerr    :    out    std_logic;
        pld10grxcrc32err    :    out    std_logic;
        pld10grxdiagstatus    :    out    std_logic_vector(1 downto 0);
        pld8grxclkout    :    out    std_logic;
        pld8gbisterr    :    out    std_logic;
        pld8grcvdclkpmab    :    out    std_logic;
        pld8gsignaldetectout    :    out    std_logic;
        pld8gbistdone    :    out    std_logic;
        pld8grlvlt    :    out    std_logic;
        pld8gfullrmf    :    out    std_logic;
        pld8gemptyrmf    :    out    std_logic;
        pld8gfullrx    :    out    std_logic;
        pld8gemptyrx    :    out    std_logic;
        pld8ga1a2k1k2flag    :    out    std_logic_vector(3 downto 0);
        pld8gbyteordflag    :    out    std_logic;
        pld8gwaboundary    :    out    std_logic_vector(4 downto 0);
        pld8grxdatavalid    :    out    std_logic_vector(3 downto 0);
        pld8grxsynchdr    :    out    std_logic_vector(1 downto 0);
        pld8grxblkstart    :    out    std_logic_vector(3 downto 0);
        pcs10grxpldclk    :    out    std_logic;
        pcs10grxpldrstn    :    out    std_logic;
        pcs10grxalignen    :    out    std_logic;
        pcs10grxalignclr    :    out    std_logic;
        pcs10grxrden    :    out    std_logic;
        pcs10grxdispclr    :    out    std_logic;
        pcs10grxclrerrblkcnt    :    out    std_logic;
        pcs10grxclrbercount    :    out    std_logic;
        pcs10grxprbserrclr    :    out    std_logic;
        pcs10grxbitslip    :    out    std_logic;
        pcs8grxurstpma    :    out    std_logic;
        pcs8grxurstpcs    :    out    std_logic;
        pcs8gcmpfifourst    :    out    std_logic;
        pcs8gphfifourstrx    :    out    std_logic;
        pcs8gencdt    :    out    std_logic;
        pcs8ga1a2size    :    out    std_logic;
        pcs8gbitslip    :    out    std_logic;
        pcs8grdenablermf    :    out    std_logic;
        pcs8gwrenablermf    :    out    std_logic;
        pcs8gpldrxclk    :    out    std_logic;
        pcs8gpolinvrx    :    out    std_logic;
        pcs8gbitlocreven    :    out    std_logic;
        pcs8gbytereven    :    out    std_logic;
        pcs8gbytordpld    :    out    std_logic;
        pcs8gwrdisablerx    :    out    std_logic;
        pcs8grdenablerx    :    out    std_logic;
        pcs8gpldextrain    :    out    std_logic_vector(3 downto 0);
        pcsgen3rxrstn    :    out    std_logic;
        pldrxclkslipout    :    out    std_logic;
        pldclkdiv33txorrx    :    out    std_logic;
        emsiprxdata    :    out    std_logic_vector(63 downto 0);
        emsippcsrxclkout    :    out    std_logic_vector(3 downto 0);
        emsippcsrxstatus    :    out    std_logic_vector(63 downto 0);
        pldrxpmarstbout    :    out    std_logic;
        pldrxplllock    :    out    std_logic;
        pld10grxfifodel    :    out    std_logic;
        pldrxiqclkout    :    out    std_logic;
        pld10grxfifoinsert    :    out    std_logic;
        pcs8gsyncsmenoutput    :    out    std_logic
    );
end component; --stratixv_hssi_rx_pld_pcs_interface


component    stratixv_hssi_tx_pcs_pma_interface
    generic    (
        lpm_type    :    string    :=    "stratixv_hssi_tx_pcs_pma_interface";
        selectpcs    :    string    :=    "eight_g_pcs"
    );
    port    (
        clockinfrompma    :    in    std_logic;
        datainfrom10gpcs    :    in    std_logic_vector(39 downto 0);
        pcs10gtxclkiqout    :    in    std_logic;
        pcsgen3txclkiqout    :    in    std_logic;
        datainfromgen3pcs    :    in    std_logic_vector(31 downto 0);
        pcs8gtxclkiqout    :    in    std_logic;
        datainfrom8gpcs    :    in    std_logic_vector(19 downto 0);
        pmaclkdiv33lcin    :    in    std_logic;
        pmatxlcplllockin    :    in    std_logic;
        pmatxcmuplllockin    :    in    std_logic;
        rtxblocksel    :    in    std_logic_vector(1 downto 0);
        pcsgen3gen3datasel    :    in    std_logic;
        pldtxpmasyncp    :    in    std_logic;
        dataouttopma    :    out    std_logic_vector(39 downto 0);
        pmatxclkout    :    out    std_logic;
        clockoutto10gpcs    :    out    std_logic;
        clockoutto8gpcs    :    out    std_logic;
        pmaclkdiv33lcout    :    out    std_logic;
        pcs10gclkdiv33lc    :    out    std_logic;
        pmatxlcplllockout    :    out    std_logic;
        pmatxcmuplllockout    :    out    std_logic;
        pmatxpmasyncp    :    out    std_logic
    );
end component; --stratixv_hssi_tx_pcs_pma_interface


component    stratixv_hssi_tx_pld_pcs_interface
    generic    (
        lpm_type    :    string    :=    "stratixv_hssi_tx_pld_pcs_interface";
        data_source    :    string    :=    "pld";
        is_10g_0ppm    :    string    :=    "false";
        is_8g_0ppm    :    string    :=    "false"
    );
    port    (
        datainfrompld    :    in    std_logic_vector(63 downto 0);
        pld10gtxpldclk    :    in    std_logic;
        pld10gtxpldrstn    :    in    std_logic;
        pld10gtxdatavalid    :    in    std_logic;
        pld10gtxcontrol    :    in    std_logic_vector(8 downto 0);
        pld10gtxbitslip    :    in    std_logic_vector(6 downto 0);
        pld10gtxdiagstatus    :    in    std_logic_vector(1 downto 0);
        pld10gtxwordslip    :    in    std_logic;
        pld10gtxbursten    :    in    std_logic;
        pld8gpldtxclk    :    in    std_logic;
        pld8gpolinvtx    :    in    std_logic;
        pld8grevloopbk    :    in    std_logic;
        pld8gwrenabletx    :    in    std_logic;
        pld8grddisabletx    :    in    std_logic;
        pld8gphfifoursttx    :    in    std_logic;
        pld8gtxboundarysel    :    in    std_logic_vector(4 downto 0);
        pld8gtxdatavalid    :    in    std_logic_vector(3 downto 0);
        pld8gtxsynchdr    :    in    std_logic_vector(1 downto 0);
        pld8gtxblkstart    :    in    std_logic_vector(3 downto 0);
        pldgen3txrstn    :    in    std_logic;
        pld8gtxurstpcs    :    in    std_logic;
        clockinfrom10gpcs    :    in    std_logic;
        pcs10gtxempty    :    in    std_logic;
        pcs10gtxpempty    :    in    std_logic;
        pcs10gtxpfull    :    in    std_logic;
        pcs10gtxfull    :    in    std_logic;
        pcs10gtxframe    :    in    std_logic;
        pcs10gtxburstenexe    :    in    std_logic;
        pcs10gtxwordslipexe    :    in    std_logic;
        pcs8gfulltx    :    in    std_logic;
        pcs8gemptytx    :    in    std_logic;
        clockinfrom8gpcs    :    in    std_logic;
        pmaclkdiv33lc    :    in    std_logic;
        emsiptxdata    :    in    std_logic_vector(63 downto 0);
        emsippcstxclkin    :    in    std_logic_vector(2 downto 0);
        emsippcstxreset    :    in    std_logic_vector(5 downto 0);
        emsippcstxctrl    :    in    std_logic_vector(43 downto 0);
        pmatxlcplllock    :    in    std_logic;
        pmatxcmuplllock    :    in    std_logic;
        pldtxpmarstbin    :    in    std_logic;
        pldlccmurstbin    :    in    std_logic;
        rtxemsip    :    in    std_logic;
        emsipenabledusermode    :    in    std_logic;
        pcs10gextraout    :    in    std_logic_vector(3 downto 0);
        pldtxpmasyncpin    :    in    std_logic;
        pcs10gtxfifoinsert    :    in    std_logic;
        pcs10gtxfifodel    :    in    std_logic;
        pld10gextrain    :    in    std_logic_vector(3 downto 0);
        pld10gtxclkout    :    out    std_logic;
        pld10gtxempty    :    out    std_logic;
        pld10gtxpempty    :    out    std_logic;
        pld10gtxpfull    :    out    std_logic;
        pld10gtxfull    :    out    std_logic;
        pld10gtxframe    :    out    std_logic;
        pld10gtxburstenexe    :    out    std_logic;
        pld10gtxwordslipexe    :    out    std_logic;
        pld8gfulltx    :    out    std_logic;
        pld8gemptytx    :    out    std_logic;
        pld8gtxclkout    :    out    std_logic;
        pcs10gtxpldclk    :    out    std_logic;
        pcs10gtxpldrstn    :    out    std_logic;
        pcs10gtxdatavalid    :    out    std_logic;
        dataoutto10gpcs    :    out    std_logic_vector(63 downto 0);
        pcs10gtxcontrol    :    out    std_logic_vector(8 downto 0);
        pcs10gtxbitslip    :    out    std_logic_vector(6 downto 0);
        pcs10gtxdiagstatus    :    out    std_logic_vector(1 downto 0);
        pcs10gtxwordslip    :    out    std_logic;
        pcs10gtxbursten    :    out    std_logic;
        pcs8gtxurstpcs    :    out    std_logic;
        dataoutto8gpcs    :    out    std_logic_vector(43 downto 0);
        pcs8gpldtxclk    :    out    std_logic;
        pcs8gpolinvtx    :    out    std_logic;
        pcs8grevloopbk    :    out    std_logic;
        pcs8gwrenabletx    :    out    std_logic;
        pcs8grddisabletx    :    out    std_logic;
        pcs8gphfifoursttx    :    out    std_logic;
        pcs8gtxboundarysel    :    out    std_logic_vector(4 downto 0);
        pcs8gtxdatavalid    :    out    std_logic_vector(3 downto 0);
        pcs8gtxsynchdr    :    out    std_logic_vector(1 downto 0);
        pcs8gtxblkstart    :    out    std_logic_vector(3 downto 0);
        pcsgen3txrstn    :    out    std_logic;
        pldclkdiv33lc    :    out    std_logic;
        emsippcstxclkout    :    out    std_logic_vector(2 downto 0);
        emsippcstxstatus    :    out    std_logic_vector(16 downto 0);
        pldtxpmarstbout    :    out    std_logic;
        pldlccmurstbout    :    out    std_logic;
        pldtxlcplllock    :    out    std_logic;
        pldtxcmuplllock    :    out    std_logic;
        pldtxiqclkout    :    out    std_logic;
        pcs10gextrain    :    out    std_logic_vector(3 downto 0);
        pld10gtxfifodel    :    out    std_logic;
        pldtxpmasyncpout    :    out    std_logic;
        pld10gtxfifoinsert    :    out    std_logic;
        pld10gextraout    :    out    std_logic_vector(3 downto 0)
    );
end component; --stratixv_hssi_tx_pld_pcs_interface

component    stratixv_hssi_avmm_interface
    port    (
    avmmrstn           : in  std_logic_vector(0 downto 0);
    avmmclk            : in  std_logic_vector(0 downto 0);
    avmmwrite          : in  std_logic_vector(0 downto 0);
    avmmread           : in  std_logic_vector(0 downto 0);
    avmmbyteen         : in  std_logic_vector(1 downto 0);
    avmmaddress        : in  std_logic_vector(10 downto 0);
    avmmwritedata      : in  std_logic_vector(15 downto 0);
    blockselect        : in  std_logic_vector(90-1 downto 0);
    readdatachnl       : in  std_logic_vector(90*16-1 downto 0);

    avmmreaddata       : out std_logic_vector(15 downto 0);

    clkchnl            : out std_logic_vector(0 downto 0);
    rstnchnl           : out std_logic_vector(0 downto 0);
    writedatachnl      : out std_logic_vector(15 downto 0);
    regaddrchnl        : out std_logic_vector(10 downto 0);
    writechnl          : out std_logic_vector(0 downto 0);
    readchnl           : out std_logic_vector(0 downto 0);
    byteenchnl         : out std_logic_vector(1 downto 0);

    -- The following ports are not modelled. They exist to match the avmm interface atom interface
    refclkdig          : in  std_logic_vector(0 downto 0);
    avmmreserevdin     : in  std_logic_vector(0 downto 0);
    
    avmmreservedout    : out std_logic_vector(0 downto 0);
    dpriorstntop       : out std_logic_vector(0 downto 0);
    dprioclktop        : out std_logic_vector(0 downto 0);
    mdiodistopchnl     : out std_logic_vector(0 downto 0);
    dpriorstnmid       : out std_logic_vector(0 downto 0);
    dprioclkmid        : out std_logic_vector(0 downto 0);
    mdiodismidchnl     : out std_logic_vector(0 downto 0);
    dpriorstnbot       : out std_logic_vector(0 downto 0);
    dprioclkbot        : out std_logic_vector(0 downto 0);
    mdiodisbotchnl     : out std_logic_vector(0 downto 0);
    dpriotestsitopchnl : out std_logic_vector(3 downto 0);
    dpriotestsimidchnl : out std_logic_vector(3 downto 0);
    dpriotestsibotchnl : out std_logic_vector(3 downto 0);
 
    -- The following ports belong to pm_adce and pm_tst_mux blocks in the PMA
    pmatestbus         : out std_logic_vector(23 downto 0);
    pmatestbussel      : in  std_logic_vector(11 downto 0);
    pmaadcestandby     : in  std_logic_vector(2 downto 0);
    pmaadcecapture     : in  std_logic_vector(2 downto 0)
   );
end component; --stratixv_hssi_avmm_interface

end STRATIXV_HSSI_COMPONENTS;

