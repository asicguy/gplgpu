///////////////////////////////////////////////////////////////////////////////
//
//  Copyright (C) 2014 Francis Bruno, All Rights Reserved
// 
//  This program is free software; you can redistribute it and/or modify it 
//  under the terms of the GNU General Public License as published by the Free 
//  Software Foundation; either version 3 of the License, or (at your option) 
//  any later version.
//
//  This program is distributed in the hope that it will be useful, but 
//  WITHOUT ANY WARRANTY; without even the implied warranty of MERCHANTABILITY 
//  or FITNESS FOR A PARTICULAR PURPOSE. 
//  See the GNU General Public License for more details.
//
//  You should have received a copy of the GNU General Public License along with
//  this program; if not, see <http://www.gnu.org/licenses>.
//
//  This code is available under licenses for commercial use. Please contact
//  Francis Bruno for more information.
//
//  http://www.gplgpu.com
//  http://www.asicsolutions.com
//
//  Title       :  CRT Controller
//  File        :  crtc.v
//  Author      :  Frank Bruno
//  Created     :  29-Dec-2005
//  RCS File    :  $Source:$
//  Status      :  $Id:$
//
//
///////////////////////////////////////////////////////////////////////////////
//
//  Description :
//   Few important signals generated by this module are
//    c_t_vsync - Vertical sync to Monitor
//    c_vert_blank - Indicates the vertical blanking period
//    c_vde - Vertical display timing strobe
//    c_pre_vde - Indicates Vertical Display will start next scan line
//    line_cmp - Indicates the succeeding lines will be in Screen B.
//
//////////////////////////////////////////////////////////////////////////////
//
//  Modules Instantiated:
//   transceiver
//   hcrt         - Horizontal CRT controller
//   vcrt         - Vertical CRT controller
//   clk_sel      - clock selection logic
//   crt_clk_gen  - CRT clock generator
//   crt_reg_dec  - Decoder CRXX and ERXX registers
//   crt_op_stage - CRT out put stage
//   crt_misc     - CRT Misc. module
//   txt_time     - Text time module
//
///////////////////////////////////////////////////////////////////////////////
//
//  Modification History:
//
//  $Log:$
//
///////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 10 ps
 module crtc
   (
    input [15:0]	h_io_addr, // Used for IO decoding.
    input   	        h_dec_3bx, // IO group decode of address range 03BX
    input   	        h_dec_3cx, // IO group decode of address range 03CX
    input   	        h_dec_3dx, // IO group decode of address range 03DX
    input   	        h_io_16,   // Indicates the current IO cycle is 16 bit.
    input               h_io_8,    // Indicates the current IO cycle is 16 bit.
    input   	        h_reset_n, // Power on reset to initialize
    input   	        h_iord,    // Indicates a read cycle.
    input   	        h_iowr,    // Indicates a write cycle.
    input               h_hclk,    // Host clock.
    input   	        t_crt_clk, // Main crt clock
    input   	        m_sr01_b0, // 8/9 dot clock
    input   	        m_sr01_b2, // shift and load 16
    input   	        m_sr01_b3, // dot clock divided by 2
    input   	        m_sr01_b4, // shift and load 32
    input               m_sr01_b5, // Disable video display control.'1' 
    input   	        a_ar10_b0, // graphics mode, graphics - 1, text - 0
    input   	        a_ar10_b5, // pixel panning compatibility
    input   	        a_ar10_b6, // pixel clock divided by 2
    input   	        t_sense_n, // switch sense bit
    input               a_arx_b5,  // Video display enable control bit
    input               a_is01_b5, // diagnostic
    input               a_is01_b4, // diagnostic
    input               m_dec_sr00_sr06, /* Valid IO decode of 03c5 
					  * index 0f 00 through 06 */
    input               m_dec_sr07, // Valid IO decode of 03c5 index of 07 
    input               m_soft_rst_n,
    input               a_ar13_b3,  // Pixel panning control bits 3-0
    input               a_ar13_b2,
    input               a_ar13_b1,
    input               a_ar13_b0,
    input [15:0] 	h_io_dbus,  // host I/O data bus
    input               vga_en,     // Disable CRT and REF reqs
    
    output [7:0] 	c_reg_ht,   // Horizontal total
    output [7:0] 	c_reg_hde,  //Horizontal Display End
    output [7:0] 	c_reg_hbs,  //Horizontal Blanking Start
    output [7:0] 	c_reg_hbe,  //Horizontal Blanking End
    output [7:0] 	c_reg_hss,  //Horizontal Sync Start
    output [7:0] 	c_reg_hse,  //Horizontal Sync End
    output [7:0] 	c_reg_cr06,
    output [7:0] 	c_reg_cr07,
    output [7:0] 	c_reg_cr10,
    output [7:0] 	c_reg_cr11,
    output [7:0] 	c_reg_cr12,
    output [7:0] 	c_reg_cr15,
    output [7:0] 	c_reg_cr16,
    output [7:0] 	c_reg_cr18,
    output [7:0] 	c_crtc_index,// crtc index register
    output [7:0] 	c_ext_index, // extension index register
    output [7:0] 	c_reg_ins0,
    output [7:0] 	c_reg_ins1,
    output [7:0] 	c_reg_fcr,   
    output [7:0] 	c_reg_cr17,
    output [7:0] 	c_reg_cr08,
    output [7:0] 	c_reg_cr09,
    output [7:0] 	c_reg_cr0a,   
    output [7:0] 	c_reg_cr0b,
    output [7:0] 	c_reg_cr14,
    output [7:0] 	c_reg_misc,
    output              c_cr24_rd,
    output              c_cr26_rd,
    output              c_9dot,
    output              c_mis_3c2_b5,
    output              c_misc_b0,
    output              c_cr0b_b5,  // Text cursor skew control 0
    output              c_cr0b_b6,  // Text cursor skew control 1
    output              c_cr0a_b5,
    output              c_cr14_b6,  // Double word mode
    output              c_cr17_b0,
    output              c_cr17_b1,
    output              c_cr17_b5,
    output              c_cr17_b6,
    output              c_gr_ext_en,  // enable Graphic's extension registers
    output [3:0]        c_ext_index_b, // lower 4 bits of ER's index register
    output              c_dec_3ba_or_3da,
    output      	c_vert_blank,  // vertical blanking period
    output  	        c_ready_n,    // current IO to CRT module is done
    output 	        c_t_clk_sel, // crt clock frequency select to pix_pll
    output  	        c_ahde,  // early horizontal display enable
    output  	        c_t_cblank_n, // composite blank to RAMDAC
    output  	        c_crt_line_end, // end of current scan line
    output  	        c_dclk_en, // Dot clock enable
    output  	        c_crt_ff_read, /* read data from CRT fifo into 
					* Attributes */
    output  	        c_shift_ld, // Load signal to Attribute serializer
    output  	        c_shift_ld_pulse, // Load signal to Attr serializer
    output  	        c_t_hsync, // Horizontal sync. to CRT monitor
    output  	        c_shift_clk, // Attribute serializer shift clock
    output  	        c_pre_vde, /* Indicates vertical display will start 
				    * next scan line */
    output  	        c_split_screen_pulse, /* Indicates screen B will start
					       * from next line untiil end of 
					       * vertical display */
    output              c_vde, // Vertical display timing strobe
    output              c_vdisp_end, // end of vertical display period.
    output  	        c_t_vsync, // Vertical sync. to CRT monitor
    output              c_attr_de, /* This signal indicates the actual display
				    * enable to the attribute control */
    output              c_uln_on, // under line on
    output              c_cursory,
    output [4:0]        c_slc_op, // scan line counter output
    output              c_row_end, // end of row
    output              c_cr0c_f13_22_hit,
    output              c_misc_b1,
    output              crt_mod_rd_en_hb,
    output              crt_mod_rd_en_lb,
    output              pre_load,
    output [10:0]       vcount
    );			 

  wire  	c_t_crt_int;
  wire 		c_raw_vsync;
  wire 		int_h_io_wr;
  wire [15:0]   crt_io_dbus;
  wire          cclk_en;
  wire          dclk_en;
  wire          pclk_en;
  wire          misc_b6;
  wire          cr11_b7;
  wire          line_cmp;
  wire          byte_pan_en;
  wire          misc_b7;
  wire          vsync_sel_ctl;
  wire          cr11_b4;
  wire          cr11_b5;
  wire          hblank;
  wire          hde;
  wire          vsync_vde;
  wire          clk_sel_strb;
  wire          final_crt_rd;
  wire          final_sh_ld;
  wire          sr_00_06_wr;
  wire          sr07_wr;
  wire          c_ahde_1;
  wire          c_ahde_1_u;
  wire          ade;
  wire          screen_off;
  wire          cr09_b5;       // Vertical Blanking start bit 9
  wire          cr09_b6;       //  Line compare bit 9
  wire          cr08_b5;
  wire          cr08_b6;
  wire          cr14_b5;
  wire          cr03_b7;      // Compatible read
  wire          misc_b0;
  wire          sel_sh_ld;
  wire          int_crt_line_end;
  wire          lncmp_zero;
  wire          txt_crt_line_end;
  wire          txt_crt_line_end_pulse;
  wire          cr17_b2;
  wire          cr17_b7;
  wire          lclk_or_by_2;
  wire          pel_pan_en;
  wire          int_split_screen_pulse;
  wire          cr17_b3;
  wire          dis_en_sta;
  
  assign        c_crt_ff_read   = final_crt_rd;
  assign        c_dclk_en       = dclk_en;
  assign        c_shift_clk     = pclk_en;
  assign        c_shift_ld      = sel_sh_ld;
  assign        c_misc_b0       = misc_b0;
   
  hcrt   HC
    (
     .m_sr01_b3                (m_sr01_b3),
     .h_reset_n                (h_reset_n),
     .cclk_en                  (cclk_en),
     .dclk_en                  (dclk_en),
     .h_hclk                   (h_hclk),
     .color_mode               (misc_b0),
     .h_io_16                  (h_io_16),
     .h_io_wr                  (int_h_io_wr),
     .h_addr                   (h_io_addr),
     .c_crtc_index             (c_crtc_index[5:0]),
     .c_ext_index              (c_ext_index),
     .misc_b6                  (misc_b6),
     .a_ar10_b0                (a_ar10_b0),
     .cr11_b7                  (cr11_b7),
     .line_cmp                 (line_cmp),
     .a_ar10_b5                (a_ar10_b5),
     .cr17_b2                  (cr17_b2),
     .byte_pan_en              (byte_pan_en),
     .cr08_b5                  (cr08_b5),
     .cr08_b6                  (cr08_b6),
     .cr17_b7                  (cr17_b7),
     .sr_00_06_wr              (sr_00_06_wr),
     .sr07_wr                  (sr07_wr),
     .t_crt_clk                (t_crt_clk),
     .h_io_dbus                (h_io_dbus[15:8]),
     
     .reg_ht                   (c_reg_ht),
     .reg_hde                  (c_reg_hde),
     .reg_hbs                  (c_reg_hbs),
     .reg_hbe                  (c_reg_hbe),
     .reg_hss                  (c_reg_hss),
     .reg_hse                  (c_reg_hse),
     .cr03_b7                  (cr03_b7),
     .c_t_hsync                (c_t_hsync),
     .c_ahde                   (c_ahde),
     .c_ahde_1                 (c_ahde_1),
     .c_ahde_1_u               (c_ahde_1_u),
     .hblank                   (hblank),
     .hde                      (hde),
     .lclk_or_by_2             (lclk_or_by_2),
     .int_crt_line_end         (int_crt_line_end)
     );


  vcrt VC
    (
     .m_soft_rst_n             (m_soft_rst_n),
     .h_reset_n                (h_reset_n),
     .h_hclk                   (h_hclk),
     .color_mode               (misc_b0),
     .h_io_16                  (h_io_16),
     .h_io_wr                  (int_h_io_wr),
     .h_addr                   (h_io_addr),
     .c_crtc_index             (c_crtc_index[5:0]),
     .c_ext_index              (c_ext_index),
     .cclk_en                  (cclk_en),
     .lclk_or_by_2             (lclk_or_by_2),
     .cr03_b7                  (cr03_b7),
     .cr17_b7                  (cr17_b7),
     .cr09_b6                  (cr09_b6),
     .cr09_b5                  (cr09_b5),
     .misc_b7                  (misc_b7),
     .vsync_sel_ctl            (vsync_sel_ctl),
     .int_crt_line_end         (int_crt_line_end),
     .t_crt_clk                (t_crt_clk),
     .h_io_dbus                (h_io_dbus[15:8]),
     .vga_en                   (vga_en),
     
     .reg_cr06                 (c_reg_cr06),
     .reg_cr07                 (c_reg_cr07),
     .reg_cr10                 (c_reg_cr10),
     .reg_cr11                 (c_reg_cr11),
     .reg_cr12                 (c_reg_cr12),
     .reg_cr15                 (c_reg_cr15),
     .reg_cr16                 (c_reg_cr16),
     .reg_cr18                 (c_reg_cr18),
     .vsync_vde                (vsync_vde),
     .cr11_b4                  (cr11_b4),
     .cr11_b5                  (cr11_b5),
     .cr11_b7                  (cr11_b7),
     .c_vde                    (c_vde),
     .c_pre_vde                (c_pre_vde),
     .c_vert_blank             (c_vert_blank),
     .c_t_vsync                (c_t_vsync),
     .line_cmp                 (line_cmp),
     .byte_pan_en              (byte_pan_en),
     .pel_pan_en               (pel_pan_en),
     .c_vdisp_end              (c_vdisp_end),
     .c_split_screen_pulse     (c_split_screen_pulse),
     .int_split_screen_pulse   (int_split_screen_pulse),
     .c_crt_line_end           (c_crt_line_end),
     .txt_crt_line_end         (txt_crt_line_end),
     .txt_crt_line_end_pulse   (txt_crt_line_end_pulse),
     .c_raw_vsync              (c_raw_vsync),
     .lncmp_zero               (lncmp_zero),
     .vcrt_cntr_op             (vcount)
     );
  
  clk_sel CS
    (
     .h_reset_n                (h_reset_n),
     .t_crt_clk                (t_crt_clk),
     .m_sr01_b3                (m_sr01_b3),
     .a_ar10_b6                (a_ar10_b6),
     .final_sh_ld              (final_sh_ld),
     .pre_load                 (pre_load),
     .cclk_en                  (cclk_en),
     
     .sel_sh_ld                (sel_sh_ld),
     .sel_sh_ld_pulse          (c_shift_ld_pulse),
     .dclk_en                  (dclk_en),
     .pclk_en                  (pclk_en)
     );
  
  crt_clk_gen CG
    (
     .t_crt_clk                (t_crt_clk),
     .line_cmp                 (line_cmp),
     .pix_pan                  (a_ar10_b5),
     .h_reset_n                (h_reset_n),
     .h_io_16                  (h_io_16),
     .h_io_wr                  (int_h_io_wr),
     .h_addr                   (h_io_addr),
     .c_ext_index              (c_ext_index),
     .m_sr01_b4                (m_sr01_b4),
     .m_sr01_b2                (m_sr01_b2),
     .m_sr01_b0                (m_sr01_b0),
     .a_ar10_b0                (a_ar10_b0),
     .a_ar10_b6                (a_ar10_b6),
     .a_ar13_b3                (a_ar13_b3),
     .a_ar13_b2                (a_ar13_b2),
     .a_ar13_b1                (a_ar13_b1),
     .a_ar13_b0                (a_ar13_b0),	 	 	 
     .cr14_b5                  (cr14_b5),
     .cr17_b3                  (cr17_b3),
     .c_ahde_1                 (c_ahde_1),
     .h_hclk                   (h_hclk),
     .ade                      (ade),
     .screen_off               (screen_off),
     .pel_pan_en               (pel_pan_en),
     .dclk_en                  (dclk_en),
     .h_io_dbus                (h_io_dbus),
     
     .reg_misc                 (c_reg_misc),
     .c_9dot                   (c_9dot),
     .misc_b0                  (misc_b0),
     .misc_b6                  (misc_b6),
     .misc_b7                  (misc_b7),
     .c_mis_3c2_b5             (c_mis_3c2_b5),
     .clk_sel_ctl              (c_t_clk_sel),
     .cclk_en                  (cclk_en),
     .final_sh_ld              (final_sh_ld),
     .final_crt_rd             (final_crt_rd),
     .c_misc_b1                (c_misc_b1),
     .pre_load                 (pre_load)
     );
  
  crt_reg_dec CD
    (
     .h_reset_n                (h_reset_n),
     .h_iord                   (h_iord),
     .h_iowr                   (h_iowr),
     .h_hclk                   (h_hclk),
     .h_io_16                  (h_io_16),
     .h_io_8                   (h_io_8),
     .misc_b0                  (misc_b0),
     .h_dec_3bx                (h_dec_3bx),
     .h_dec_3cx                (h_dec_3cx),
     .h_dec_3dx                (h_dec_3dx),
     .m_dec_sr07               (m_dec_sr07),
     .m_dec_sr00_sr06          (m_dec_sr00_sr06),
     .h_io_addr                (h_io_addr),
     .h_io_dbus                (h_io_dbus),

     .crtc_index               (c_crtc_index),
     .ext_index                (c_ext_index),
     .trim_wr                  (int_h_io_wr),
     .c_gr_ext_en              (c_gr_ext_en),
     .c_ext_index_b            (c_ext_index_b),
     .crt_mod_rd_en_hb         (crt_mod_rd_en_hb),
     .crt_mod_rd_en_lb         (crt_mod_rd_en_lb),
     .c_ready_n                (c_ready_n),
     .sr_00_06_wr              (sr_00_06_wr),
     .sr07_wr                  (sr07_wr),
     .cr24_rd                  (c_cr24_rd),
     .cr26_rd                  (c_cr26_rd),
     .c_dec_3ba_or_3da         (c_dec_3ba_or_3da),
     .c_cr0c_f13_22_hit        (c_cr0c_f13_22_hit)
     );
  

  crt_op_stage CO
    (
     .h_reset_n                (h_reset_n),
     .c_vde                    (c_vde),
     .cr11_b4                  (cr11_b4),
     .cr11_b5                  (cr11_b5),
     .a_arx_b5                 (a_arx_b5),
     .m_sr01_b5                (m_sr01_b5),
     .vblank                   (c_vert_blank),
     .hblank                   (hblank),
     .cclk_en                  (cclk_en),
     .dclk_en                  (dclk_en),
     .hde                      (hde),      
     .c_ahde                   (c_ahde),
     .int_crt_line_end         (int_crt_line_end),
     .t_crt_clk                (t_crt_clk),
     .a_ar10_b0                (a_ar10_b0),
     .vga_en                   (vga_en),
     
     .c_t_crt_int              (c_t_crt_int),
     .c_attr_de                (c_attr_de),
     .c_t_cblank_n             (c_t_cblank_n),
     .ade                      (ade),
     .screen_off               (screen_off),
     .dis_en_sta               (dis_en_sta)
     );
  
  crt_misc CM
    (
     .dis_en_sta               (dis_en_sta), 
     .c_raw_vsync              (c_raw_vsync),
     .h_reset_n                (h_reset_n),
     .h_hclk                   (h_hclk),
     .color_mode               (misc_b0),
     .h_io_16                  (h_io_16),
     .h_io_wr                  (int_h_io_wr),
     .h_addr                   (h_io_addr),
     .c_crtc_index             (c_crtc_index[5:0]),
     .c_ext_index              (c_ext_index),
     .t_sense_n                (t_sense_n),
     .c_t_crt_int              (c_t_crt_int),
     .a_is01_b5                (a_is01_b5),
     .a_is01_b4                (a_is01_b4),
     .vsync_vde                (vsync_vde),
     .h_io_dbus                (h_io_dbus),
     
     .reg_ins0                 (c_reg_ins0),
     .reg_ins1                 (c_reg_ins1),
     .reg_fcr                  (c_reg_fcr),   
     .reg_cr17                 (c_reg_cr17),
     .c_cr17_b0                (c_cr17_b0),
     .c_cr17_b1                (c_cr17_b1),
     .cr17_b2                  (cr17_b2),
     .cr17_b3                  (cr17_b3),
     .c_cr17_b5                (c_cr17_b5),
     .c_cr17_b6                (c_cr17_b6),
     .cr17_b7                  (cr17_b7),
     .vsync_sel_ctl            (vsync_sel_ctl)
     );

  txt_time   CT
    (
     .h_reset_n                (h_reset_n),
     .h_hclk                   (h_hclk),
     .color_mode               (misc_b0),
     .h_io_16                  (h_io_16),
     .h_io_wr                  (int_h_io_wr),
     .h_addr                   (h_io_addr),
     .c_crtc_index             (c_crtc_index[5:0]),
     .t_crt_clk                (t_crt_clk),
     .cclk_en                  (cclk_en),       // character clock
     .dclk_en                  (dclk_en),
     .int_pre_vde              (c_pre_vde), /* Indicates Vertical Display will
					     * start next scan line */
     .int_split_screen_pulse   (int_split_screen_pulse),
     .txt_crt_line_end         (txt_crt_line_end),
     .txt_crt_line_end_pulse   (txt_crt_line_end_pulse),
     .c_vdisp_end              (c_vdisp_end),
     .lncmp_zero               (lncmp_zero),
     .h_io_dbus                (h_io_dbus[15:8]),       // data bus
     
     .reg_cr08                 (c_reg_cr08),
     .reg_cr09                 (c_reg_cr09),
     .reg_cr0a                 (c_reg_cr0a),   
     .reg_cr0b                 (c_reg_cr0b),
     .reg_cr14                 (c_reg_cr14),
     .cr08_b5                  (cr08_b5),
     .cr08_b6                  (cr08_b6),
     .cr09_b5                  (cr09_b5),    // Vertical Blanking start bit 9
     .cr09_b6                  (cr09_b6),    // Line compare bit 9
     .c_cr0b_b5                (c_cr0b_b5),  // Text cursor skew control bit 0
     .c_cr0b_b6                (c_cr0b_b6),  // Text cursor skew control bit 1
     .c_cr0a_b5                (c_cr0a_b5),  // Disable Text cursor
     .cr14_b5                  (cr14_b5),    // Count by four
     .c_cr14_b6                (c_cr14_b6),  // Double word mode
     .c_uln_on                 (c_uln_on),   // under line on
     .c_cursor_on_line         (c_cursory), 
     .c_slc_op                 (c_slc_op),   // scan line counter output
     .c_row_end                (c_row_end)   // end of row
     );
endmodule

